// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:44:57"

// 
// Device: Altera 1SG280LU2F50E2VG Package FBGA2397
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_s10_12x12x32 (
	dout,
	clk,
	din_a,
	din_b);
output 	[27:0] dout;
input 	clk;
input 	[383:0] din_a;
input 	[383:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_12 ;
wire Xd_0__inst_inst_inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_17 ;
wire Xd_0__inst_inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_32 ;
wire Xd_0__inst_inst_inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_37 ;
wire Xd_0__inst_inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_52 ;
wire Xd_0__inst_inst_inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_57 ;
wire Xd_0__inst_inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_72 ;
wire Xd_0__inst_inst_inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_77 ;
wire Xd_0__inst_inst_inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_82 ;
wire Xd_0__inst_inst_inst_inst_add_0_86_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_87 ;
wire Xd_0__inst_inst_inst_inst_add_0_91_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_92 ;
wire Xd_0__inst_inst_inst_inst_add_0_96_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_97 ;
wire Xd_0__inst_inst_inst_inst_add_0_101_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_102 ;
wire Xd_0__inst_inst_inst_inst_add_0_106_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_107 ;
wire Xd_0__inst_inst_inst_inst_add_0_111_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_112 ;
wire Xd_0__inst_inst_inst_inst_add_0_116_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_117 ;
wire Xd_0__inst_inst_inst_inst_add_0_121_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_122 ;
wire Xd_0__inst_inst_inst_inst_add_0_126_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_127 ;
wire Xd_0__inst_inst_inst_inst_add_0_131_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_132 ;
wire Xd_0__inst_inst_inst_inst_add_0_136_sumout ;
wire Xd_0__inst_mult_2_205 ;
wire Xd_0__inst_mult_2_206 ;
wire Xd_0__inst_inst_inst_add_1_1_sumout ;
wire Xd_0__inst_inst_inst_add_1_2 ;
wire Xd_0__inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_add_0_2 ;
wire Xd_0__inst_mult_2_210 ;
wire Xd_0__inst_mult_2_211 ;
wire Xd_0__inst_inst_inst_add_1_6_sumout ;
wire Xd_0__inst_inst_inst_add_1_7 ;
wire Xd_0__inst_inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_add_1_11_sumout ;
wire Xd_0__inst_inst_inst_add_1_12 ;
wire Xd_0__inst_inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_inst_add_0_12 ;
wire Xd_0__inst_inst_inst_add_1_16_sumout ;
wire Xd_0__inst_inst_inst_add_1_17 ;
wire Xd_0__inst_inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_inst_add_0_17 ;
wire Xd_0__inst_inst_inst_add_1_21_sumout ;
wire Xd_0__inst_inst_inst_add_1_22 ;
wire Xd_0__inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_add_1_26_sumout ;
wire Xd_0__inst_inst_inst_add_1_27 ;
wire Xd_0__inst_inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_add_1_31_sumout ;
wire Xd_0__inst_inst_inst_add_1_32 ;
wire Xd_0__inst_inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_inst_add_0_32 ;
wire Xd_0__inst_inst_inst_add_1_36_sumout ;
wire Xd_0__inst_inst_inst_add_1_37 ;
wire Xd_0__inst_inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_inst_add_0_37 ;
wire Xd_0__inst_inst_inst_add_1_41_sumout ;
wire Xd_0__inst_inst_inst_add_1_42 ;
wire Xd_0__inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_add_1_46_sumout ;
wire Xd_0__inst_inst_inst_add_1_47 ;
wire Xd_0__inst_inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_add_1_51_sumout ;
wire Xd_0__inst_inst_inst_add_1_52 ;
wire Xd_0__inst_inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_inst_add_0_52 ;
wire Xd_0__inst_inst_inst_add_1_56_sumout ;
wire Xd_0__inst_inst_inst_add_1_57 ;
wire Xd_0__inst_inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_inst_add_0_57 ;
wire Xd_0__inst_inst_inst_add_1_61_sumout ;
wire Xd_0__inst_inst_inst_add_1_62 ;
wire Xd_0__inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_add_1_66_sumout ;
wire Xd_0__inst_inst_inst_add_1_67 ;
wire Xd_0__inst_inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_add_1_71_sumout ;
wire Xd_0__inst_inst_inst_add_1_72 ;
wire Xd_0__inst_inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_inst_add_0_72 ;
wire Xd_0__inst_inst_inst_add_1_76_sumout ;
wire Xd_0__inst_inst_inst_add_1_77 ;
wire Xd_0__inst_inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_inst_add_0_77 ;
wire Xd_0__inst_inst_inst_add_1_81_sumout ;
wire Xd_0__inst_inst_inst_add_1_82 ;
wire Xd_0__inst_inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_inst_add_0_82 ;
wire Xd_0__inst_inst_inst_add_1_86_sumout ;
wire Xd_0__inst_inst_inst_add_1_87 ;
wire Xd_0__inst_inst_inst_add_0_86_sumout ;
wire Xd_0__inst_inst_inst_add_0_87 ;
wire Xd_0__inst_inst_inst_add_1_91_sumout ;
wire Xd_0__inst_inst_inst_add_1_92 ;
wire Xd_0__inst_inst_inst_add_0_91_sumout ;
wire Xd_0__inst_inst_inst_add_0_92 ;
wire Xd_0__inst_inst_inst_add_1_96_sumout ;
wire Xd_0__inst_inst_inst_add_1_97 ;
wire Xd_0__inst_inst_inst_add_0_96_sumout ;
wire Xd_0__inst_inst_inst_add_0_97 ;
wire Xd_0__inst_inst_inst_add_1_101_sumout ;
wire Xd_0__inst_inst_inst_add_1_102 ;
wire Xd_0__inst_inst_inst_add_0_101_sumout ;
wire Xd_0__inst_inst_inst_add_0_102 ;
wire Xd_0__inst_inst_inst_add_1_106_sumout ;
wire Xd_0__inst_inst_inst_add_1_107 ;
wire Xd_0__inst_inst_inst_add_0_106_sumout ;
wire Xd_0__inst_inst_inst_add_0_107 ;
wire Xd_0__inst_inst_inst_add_1_111_sumout ;
wire Xd_0__inst_inst_inst_add_1_112 ;
wire Xd_0__inst_inst_inst_add_0_111_sumout ;
wire Xd_0__inst_inst_inst_add_0_112 ;
wire Xd_0__inst_inst_inst_add_1_116_sumout ;
wire Xd_0__inst_inst_inst_add_1_117 ;
wire Xd_0__inst_inst_inst_add_0_116_sumout ;
wire Xd_0__inst_inst_inst_add_0_117 ;
wire Xd_0__inst_inst_inst_add_1_121_sumout ;
wire Xd_0__inst_inst_inst_add_1_122 ;
wire Xd_0__inst_inst_inst_add_0_121_sumout ;
wire Xd_0__inst_inst_inst_add_0_122 ;
wire Xd_0__inst_inst_inst_add_1_126_sumout ;
wire Xd_0__inst_inst_inst_add_1_127 ;
wire Xd_0__inst_inst_inst_add_0_126_sumout ;
wire Xd_0__inst_inst_inst_add_0_127 ;
wire Xd_0__inst_inst_inst_add_1_131_sumout ;
wire Xd_0__inst_inst_inst_add_0_131_sumout ;
wire Xd_0__inst_mult_26_205 ;
wire Xd_0__inst_mult_26_206 ;
wire Xd_0__inst_mult_24_205 ;
wire Xd_0__inst_mult_24_206 ;
wire Xd_0__inst_mult_2_214 ;
wire Xd_0__inst_mult_2_215 ;
wire Xd_0__inst_inst_add_3_1_sumout ;
wire Xd_0__inst_inst_add_3_2 ;
wire Xd_0__inst_inst_add_2_1_sumout ;
wire Xd_0__inst_inst_add_2_2 ;
wire Xd_0__inst_mult_26_210 ;
wire Xd_0__inst_mult_26_35_sumout ;
wire Xd_0__inst_mult_26_36 ;
wire Xd_0__inst_mult_26_214 ;
wire Xd_0__inst_mult_26_215 ;
wire Xd_0__inst_inst_add_1_1_sumout ;
wire Xd_0__inst_inst_add_1_2 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_mult_24_210 ;
wire Xd_0__inst_mult_24_35_sumout ;
wire Xd_0__inst_mult_24_36 ;
wire Xd_0__inst_mult_24_214 ;
wire Xd_0__inst_mult_24_215 ;
wire Xd_0__inst_mult_2_219 ;
wire Xd_0__inst_mult_2_220 ;
wire Xd_0__inst_inst_add_3_6_sumout ;
wire Xd_0__inst_inst_add_3_7 ;
wire Xd_0__inst_inst_add_2_6_sumout ;
wire Xd_0__inst_inst_add_2_7 ;
wire Xd_0__inst_inst_add_1_6_sumout ;
wire Xd_0__inst_inst_add_1_7 ;
wire Xd_0__inst_inst_add_0_6_sumout ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_3_11_sumout ;
wire Xd_0__inst_inst_add_3_12 ;
wire Xd_0__inst_inst_add_2_11_sumout ;
wire Xd_0__inst_inst_add_2_12 ;
wire Xd_0__inst_inst_add_1_11_sumout ;
wire Xd_0__inst_inst_add_1_12 ;
wire Xd_0__inst_inst_add_0_11_sumout ;
wire Xd_0__inst_inst_add_0_12 ;
wire Xd_0__inst_inst_add_3_16_sumout ;
wire Xd_0__inst_inst_add_3_17 ;
wire Xd_0__inst_inst_add_2_16_sumout ;
wire Xd_0__inst_inst_add_2_17 ;
wire Xd_0__inst_inst_add_1_16_sumout ;
wire Xd_0__inst_inst_add_1_17 ;
wire Xd_0__inst_inst_add_0_16_sumout ;
wire Xd_0__inst_inst_add_0_17 ;
wire Xd_0__inst_inst_add_3_21_sumout ;
wire Xd_0__inst_inst_add_3_22 ;
wire Xd_0__inst_inst_add_2_21_sumout ;
wire Xd_0__inst_inst_add_2_22 ;
wire Xd_0__inst_inst_add_1_21_sumout ;
wire Xd_0__inst_inst_add_1_22 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_3_26_sumout ;
wire Xd_0__inst_inst_add_3_27 ;
wire Xd_0__inst_inst_add_2_26_sumout ;
wire Xd_0__inst_inst_add_2_27 ;
wire Xd_0__inst_inst_add_1_26_sumout ;
wire Xd_0__inst_inst_add_1_27 ;
wire Xd_0__inst_inst_add_0_26_sumout ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_3_31_sumout ;
wire Xd_0__inst_inst_add_3_32 ;
wire Xd_0__inst_inst_add_2_31_sumout ;
wire Xd_0__inst_inst_add_2_32 ;
wire Xd_0__inst_inst_add_1_31_sumout ;
wire Xd_0__inst_inst_add_1_32 ;
wire Xd_0__inst_inst_add_0_31_sumout ;
wire Xd_0__inst_inst_add_0_32 ;
wire Xd_0__inst_inst_add_3_36_sumout ;
wire Xd_0__inst_inst_add_3_37 ;
wire Xd_0__inst_inst_add_2_36_sumout ;
wire Xd_0__inst_inst_add_2_37 ;
wire Xd_0__inst_inst_add_1_36_sumout ;
wire Xd_0__inst_inst_add_1_37 ;
wire Xd_0__inst_inst_add_0_36_sumout ;
wire Xd_0__inst_inst_add_0_37 ;
wire Xd_0__inst_inst_add_3_41_sumout ;
wire Xd_0__inst_inst_add_3_42 ;
wire Xd_0__inst_inst_add_2_41_sumout ;
wire Xd_0__inst_inst_add_2_42 ;
wire Xd_0__inst_inst_add_1_41_sumout ;
wire Xd_0__inst_inst_add_1_42 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_3_46_sumout ;
wire Xd_0__inst_inst_add_3_47 ;
wire Xd_0__inst_inst_add_2_46_sumout ;
wire Xd_0__inst_inst_add_2_47 ;
wire Xd_0__inst_inst_add_1_46_sumout ;
wire Xd_0__inst_inst_add_1_47 ;
wire Xd_0__inst_inst_add_0_46_sumout ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_3_51_sumout ;
wire Xd_0__inst_inst_add_3_52 ;
wire Xd_0__inst_inst_add_2_51_sumout ;
wire Xd_0__inst_inst_add_2_52 ;
wire Xd_0__inst_inst_add_1_51_sumout ;
wire Xd_0__inst_inst_add_1_52 ;
wire Xd_0__inst_inst_add_0_51_sumout ;
wire Xd_0__inst_inst_add_0_52 ;
wire Xd_0__inst_inst_add_3_56_sumout ;
wire Xd_0__inst_inst_add_3_57 ;
wire Xd_0__inst_inst_add_2_56_sumout ;
wire Xd_0__inst_inst_add_2_57 ;
wire Xd_0__inst_inst_add_1_56_sumout ;
wire Xd_0__inst_inst_add_1_57 ;
wire Xd_0__inst_inst_add_0_56_sumout ;
wire Xd_0__inst_inst_add_0_57 ;
wire Xd_0__inst_inst_add_3_61_sumout ;
wire Xd_0__inst_inst_add_3_62 ;
wire Xd_0__inst_inst_add_2_61_sumout ;
wire Xd_0__inst_inst_add_2_62 ;
wire Xd_0__inst_inst_add_1_61_sumout ;
wire Xd_0__inst_inst_add_1_62 ;
wire Xd_0__inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_add_0_62 ;
wire Xd_0__inst_inst_add_3_66_sumout ;
wire Xd_0__inst_inst_add_3_67 ;
wire Xd_0__inst_inst_add_2_66_sumout ;
wire Xd_0__inst_inst_add_2_67 ;
wire Xd_0__inst_inst_add_1_66_sumout ;
wire Xd_0__inst_inst_add_1_67 ;
wire Xd_0__inst_inst_add_0_66_sumout ;
wire Xd_0__inst_inst_add_0_67 ;
wire Xd_0__inst_inst_add_3_71_sumout ;
wire Xd_0__inst_inst_add_3_72 ;
wire Xd_0__inst_inst_add_2_71_sumout ;
wire Xd_0__inst_inst_add_2_72 ;
wire Xd_0__inst_inst_add_1_71_sumout ;
wire Xd_0__inst_inst_add_1_72 ;
wire Xd_0__inst_inst_add_0_71_sumout ;
wire Xd_0__inst_inst_add_0_72 ;
wire Xd_0__inst_inst_add_3_76_sumout ;
wire Xd_0__inst_inst_add_3_77 ;
wire Xd_0__inst_inst_add_2_76_sumout ;
wire Xd_0__inst_inst_add_2_77 ;
wire Xd_0__inst_inst_add_1_76_sumout ;
wire Xd_0__inst_inst_add_1_77 ;
wire Xd_0__inst_inst_add_0_76_sumout ;
wire Xd_0__inst_inst_add_0_77 ;
wire Xd_0__inst_inst_add_3_81_sumout ;
wire Xd_0__inst_inst_add_3_82 ;
wire Xd_0__inst_inst_add_2_81_sumout ;
wire Xd_0__inst_inst_add_2_82 ;
wire Xd_0__inst_inst_add_1_81_sumout ;
wire Xd_0__inst_inst_add_1_82 ;
wire Xd_0__inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_add_0_82 ;
wire Xd_0__inst_inst_add_3_86_sumout ;
wire Xd_0__inst_inst_add_3_87 ;
wire Xd_0__inst_inst_add_2_86_sumout ;
wire Xd_0__inst_inst_add_2_87 ;
wire Xd_0__inst_inst_add_1_86_sumout ;
wire Xd_0__inst_inst_add_1_87 ;
wire Xd_0__inst_inst_add_0_86_sumout ;
wire Xd_0__inst_inst_add_0_87 ;
wire Xd_0__inst_inst_add_3_91_sumout ;
wire Xd_0__inst_inst_add_3_92 ;
wire Xd_0__inst_inst_add_2_91_sumout ;
wire Xd_0__inst_inst_add_2_92 ;
wire Xd_0__inst_inst_add_1_91_sumout ;
wire Xd_0__inst_inst_add_1_92 ;
wire Xd_0__inst_inst_add_0_91_sumout ;
wire Xd_0__inst_inst_add_0_92 ;
wire Xd_0__inst_inst_add_3_96_sumout ;
wire Xd_0__inst_inst_add_3_97 ;
wire Xd_0__inst_inst_add_2_96_sumout ;
wire Xd_0__inst_inst_add_2_97 ;
wire Xd_0__inst_inst_add_1_96_sumout ;
wire Xd_0__inst_inst_add_1_97 ;
wire Xd_0__inst_inst_add_0_96_sumout ;
wire Xd_0__inst_inst_add_0_97 ;
wire Xd_0__inst_inst_add_3_101_sumout ;
wire Xd_0__inst_inst_add_3_102 ;
wire Xd_0__inst_inst_add_2_101_sumout ;
wire Xd_0__inst_inst_add_2_102 ;
wire Xd_0__inst_inst_add_1_101_sumout ;
wire Xd_0__inst_inst_add_1_102 ;
wire Xd_0__inst_inst_add_0_101_sumout ;
wire Xd_0__inst_inst_add_0_102 ;
wire Xd_0__inst_inst_add_3_106_sumout ;
wire Xd_0__inst_inst_add_3_107 ;
wire Xd_0__inst_inst_add_2_106_sumout ;
wire Xd_0__inst_inst_add_2_107 ;
wire Xd_0__inst_inst_add_1_106_sumout ;
wire Xd_0__inst_inst_add_1_107 ;
wire Xd_0__inst_inst_add_0_106_sumout ;
wire Xd_0__inst_inst_add_0_107 ;
wire Xd_0__inst_inst_add_3_111_sumout ;
wire Xd_0__inst_inst_add_3_112 ;
wire Xd_0__inst_inst_add_2_111_sumout ;
wire Xd_0__inst_inst_add_2_112 ;
wire Xd_0__inst_inst_add_1_111_sumout ;
wire Xd_0__inst_inst_add_1_112 ;
wire Xd_0__inst_inst_add_0_111_sumout ;
wire Xd_0__inst_inst_add_0_112 ;
wire Xd_0__inst_inst_add_3_116_sumout ;
wire Xd_0__inst_inst_add_3_117 ;
wire Xd_0__inst_inst_add_2_116_sumout ;
wire Xd_0__inst_inst_add_2_117 ;
wire Xd_0__inst_inst_add_1_116_sumout ;
wire Xd_0__inst_inst_add_1_117 ;
wire Xd_0__inst_inst_add_0_116_sumout ;
wire Xd_0__inst_inst_add_0_117 ;
wire Xd_0__inst_inst_add_3_121_sumout ;
wire Xd_0__inst_inst_add_3_122 ;
wire Xd_0__inst_inst_add_2_121_sumout ;
wire Xd_0__inst_inst_add_2_122 ;
wire Xd_0__inst_inst_add_1_121_sumout ;
wire Xd_0__inst_inst_add_1_122 ;
wire Xd_0__inst_inst_add_0_121_sumout ;
wire Xd_0__inst_inst_add_0_122 ;
wire Xd_0__inst_inst_add_3_126_sumout ;
wire Xd_0__inst_inst_add_2_126_sumout ;
wire Xd_0__inst_inst_add_1_126_sumout ;
wire Xd_0__inst_inst_add_0_126_sumout ;
wire Xd_0__inst_mult_25_205 ;
wire Xd_0__inst_mult_25_206 ;
wire Xd_0__inst_mult_24_219 ;
wire Xd_0__inst_mult_24_220 ;
wire Xd_0__inst_mult_26_219 ;
wire Xd_0__inst_mult_26_220 ;
wire Xd_0__inst_mult_27_35_sumout ;
wire Xd_0__inst_mult_27_36 ;
wire Xd_0__inst_mult_26_40_sumout ;
wire Xd_0__inst_mult_26_41 ;
wire Xd_0__inst_mult_26_224 ;
wire Xd_0__inst_mult_26_225 ;
wire Xd_0__inst_mult_27_205 ;
wire Xd_0__inst_mult_27_206 ;
wire Xd_0__inst_mult_26_229 ;
wire Xd_0__inst_mult_26_230 ;
wire Xd_0__inst_mult_24_224 ;
wire Xd_0__inst_mult_24_225 ;
wire Xd_0__inst_mult_24_40_sumout ;
wire Xd_0__inst_mult_24_41 ;
wire Xd_0__inst_mult_24_229 ;
wire Xd_0__inst_mult_24_230 ;
wire Xd_0__inst_mult_2_224 ;
wire Xd_0__inst_mult_2_225 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_25_210 ;
wire Xd_0__inst_mult_25_35_sumout ;
wire Xd_0__inst_mult_25_36 ;
wire Xd_0__inst_mult_25_214 ;
wire Xd_0__inst_mult_25_215 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_24_234 ;
wire Xd_0__inst_mult_24_45_sumout ;
wire Xd_0__inst_mult_24_46 ;
wire Xd_0__inst_mult_24_239 ;
wire Xd_0__inst_mult_24_240 ;
wire Xd_0__inst_mult_26_234 ;
wire Xd_0__inst_mult_26_235 ;
wire Xd_0__inst_mult_26_239 ;
wire Xd_0__inst_mult_26_240 ;
wire Xd_0__inst_mult_27_40_sumout ;
wire Xd_0__inst_mult_27_41 ;
wire Xd_0__inst_mult_26_244 ;
wire Xd_0__inst_mult_26_249 ;
wire Xd_0__inst_mult_26_250 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_27_210 ;
wire Xd_0__inst_mult_27_45_sumout ;
wire Xd_0__inst_mult_27_46 ;
wire Xd_0__inst_mult_27_214 ;
wire Xd_0__inst_mult_27_215 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_2 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_2 ;
wire Xd_0__inst_mult_26_254 ;
wire Xd_0__inst_mult_26_45_sumout ;
wire Xd_0__inst_mult_26_46 ;
wire Xd_0__inst_mult_26_259 ;
wire Xd_0__inst_mult_26_260 ;
wire Xd_0__inst_mult_24_244 ;
wire Xd_0__inst_mult_24_245 ;
wire Xd_0__inst_mult_24_249 ;
wire Xd_0__inst_mult_24_250 ;
wire Xd_0__inst_mult_25_40_sumout ;
wire Xd_0__inst_mult_25_41 ;
wire Xd_0__inst_mult_24_254 ;
wire Xd_0__inst_mult_24_259 ;
wire Xd_0__inst_mult_24_260 ;
wire Xd_0__inst_mult_2_229 ;
wire Xd_0__inst_mult_2_230 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_7 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_12 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_17 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_22 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_27 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_32 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_37 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_42 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_47 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_52 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_57 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_62 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_67 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_72 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_77 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_82 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_86_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_87 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_91_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_92 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_96_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_97 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_101_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_102 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_106_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_107 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_111_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_112 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_116_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_117 ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_121_sumout ;
wire Xd_0__inst_a2_7__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_a2_6__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_mult_25_219 ;
wire Xd_0__inst_mult_25_220 ;
wire Xd_0__inst_mult_30_35_sumout ;
wire Xd_0__inst_mult_30_36 ;
wire Xd_0__inst_mult_25_45_sumout ;
wire Xd_0__inst_mult_25_46 ;
wire Xd_0__inst_mult_25_224 ;
wire Xd_0__inst_mult_25_225 ;
wire Xd_0__inst_a2_5__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_a2_4__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_mult_24_264 ;
wire Xd_0__inst_mult_24_265 ;
wire Xd_0__inst_mult_24_50_sumout ;
wire Xd_0__inst_mult_24_51 ;
wire Xd_0__inst_mult_24_269 ;
wire Xd_0__inst_mult_24_270 ;
wire Xd_0__inst_mult_26_264 ;
wire Xd_0__inst_mult_26_265 ;
wire Xd_0__inst_mult_26_269 ;
wire Xd_0__inst_mult_26_270 ;
wire Xd_0__inst_mult_26_274 ;
wire Xd_0__inst_mult_26_275 ;
wire Xd_0__inst_mult_26_279 ;
wire Xd_0__inst_mult_26_280 ;
wire Xd_0__inst_a2_3__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_a2_2__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_mult_27_219 ;
wire Xd_0__inst_mult_27_220 ;
wire Xd_0__inst_mult_27_50_sumout ;
wire Xd_0__inst_mult_27_51 ;
wire Xd_0__inst_mult_27_224 ;
wire Xd_0__inst_mult_27_225 ;
wire Xd_0__inst_a2_1__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_a2_0__adder2_inst_add_0_127_cout ;
wire Xd_0__inst_mult_26_284 ;
wire Xd_0__inst_mult_26_285 ;
wire Xd_0__inst_mult_26_50_sumout ;
wire Xd_0__inst_mult_26_51 ;
wire Xd_0__inst_mult_26_289 ;
wire Xd_0__inst_mult_26_290 ;
wire Xd_0__inst_mult_24_274 ;
wire Xd_0__inst_mult_24_275 ;
wire Xd_0__inst_mult_24_279 ;
wire Xd_0__inst_mult_24_280 ;
wire Xd_0__inst_mult_24_284 ;
wire Xd_0__inst_mult_24_285 ;
wire Xd_0__inst_mult_24_289 ;
wire Xd_0__inst_mult_24_290 ;
wire Xd_0__inst_mult_2_234 ;
wire Xd_0__inst_mult_2_235 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_21_205 ;
wire Xd_0__inst_mult_21_206 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_20_205 ;
wire Xd_0__inst_mult_20_206 ;
wire Xd_0__inst_mult_25_229 ;
wire Xd_0__inst_mult_25_234 ;
wire Xd_0__inst_mult_25_235 ;
wire Xd_0__inst_mult_25_239 ;
wire Xd_0__inst_mult_25_244 ;
wire Xd_0__inst_mult_25_245 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_23_205 ;
wire Xd_0__inst_mult_23_206 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_22_205 ;
wire Xd_0__inst_mult_22_206 ;
wire Xd_0__inst_mult_24_294 ;
wire Xd_0__inst_mult_24_299 ;
wire Xd_0__inst_mult_24_300 ;
wire Xd_0__inst_mult_24_304 ;
wire Xd_0__inst_mult_24_309 ;
wire Xd_0__inst_mult_24_310 ;
wire Xd_0__inst_mult_26_294 ;
wire Xd_0__inst_mult_26_295 ;
wire Xd_0__inst_mult_26_299 ;
wire Xd_0__inst_mult_26_300 ;
wire Xd_0__inst_mult_26_304 ;
wire Xd_0__inst_mult_26_309 ;
wire Xd_0__inst_mult_26_310 ;
wire Xd_0__inst_mult_26_314 ;
wire Xd_0__inst_mult_26_315 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_19_205 ;
wire Xd_0__inst_mult_19_206 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_17_205 ;
wire Xd_0__inst_mult_17_206 ;
wire Xd_0__inst_mult_27_229 ;
wire Xd_0__inst_mult_27_234 ;
wire Xd_0__inst_mult_27_235 ;
wire Xd_0__inst_mult_27_239 ;
wire Xd_0__inst_mult_27_244 ;
wire Xd_0__inst_mult_27_245 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_16_205 ;
wire Xd_0__inst_mult_16_206 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_2 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_2 ;
wire Xd_0__inst_mult_29_205 ;
wire Xd_0__inst_mult_29_206 ;
wire Xd_0__inst_mult_26_319 ;
wire Xd_0__inst_mult_26_324 ;
wire Xd_0__inst_mult_26_325 ;
wire Xd_0__inst_mult_26_329 ;
wire Xd_0__inst_mult_26_334 ;
wire Xd_0__inst_mult_26_335 ;
wire Xd_0__inst_mult_24_314 ;
wire Xd_0__inst_mult_24_315 ;
wire Xd_0__inst_mult_24_319 ;
wire Xd_0__inst_mult_24_320 ;
wire Xd_0__inst_mult_24_324 ;
wire Xd_0__inst_mult_24_329 ;
wire Xd_0__inst_mult_24_330 ;
wire Xd_0__inst_mult_24_334 ;
wire Xd_0__inst_mult_24_335 ;
wire Xd_0__inst_mult_2_239 ;
wire Xd_0__inst_mult_2_240 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_7 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_12 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_17 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_22 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_27 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_32 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_37 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_42 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_47 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_52 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_57 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_62 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_67 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_72 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_77 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_82 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_86_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_87 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_91_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_92 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_96_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_97 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_101_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_102 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_106_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_107 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_111_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_112 ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_116_sumout ;
wire Xd_0__inst_a1_15__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_14__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_21_210 ;
wire Xd_0__inst_mult_21_35_sumout ;
wire Xd_0__inst_mult_21_36 ;
wire Xd_0__inst_mult_21_214 ;
wire Xd_0__inst_mult_21_215 ;
wire Xd_0__inst_a1_13__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_12__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_20_210 ;
wire Xd_0__inst_mult_20_35_sumout ;
wire Xd_0__inst_mult_20_36 ;
wire Xd_0__inst_mult_20_214 ;
wire Xd_0__inst_mult_20_215 ;
wire Xd_0__inst_mult_25_249 ;
wire Xd_0__inst_mult_25_250 ;
wire Xd_0__inst_mult_25_254 ;
wire Xd_0__inst_mult_25_255 ;
wire Xd_0__inst_mult_25_259 ;
wire Xd_0__inst_mult_25_260 ;
wire Xd_0__inst_mult_25_264 ;
wire Xd_0__inst_mult_25_265 ;
wire Xd_0__inst_a1_11__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_10__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_23_210 ;
wire Xd_0__inst_mult_23_35_sumout ;
wire Xd_0__inst_mult_23_36 ;
wire Xd_0__inst_mult_23_214 ;
wire Xd_0__inst_mult_23_215 ;
wire Xd_0__inst_a1_9__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_8__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_22_210 ;
wire Xd_0__inst_mult_22_35_sumout ;
wire Xd_0__inst_mult_22_36 ;
wire Xd_0__inst_mult_22_214 ;
wire Xd_0__inst_mult_22_215 ;
wire Xd_0__inst_mult_24_339 ;
wire Xd_0__inst_mult_24_340 ;
wire Xd_0__inst_mult_24_344 ;
wire Xd_0__inst_mult_24_345 ;
wire Xd_0__inst_mult_24_349 ;
wire Xd_0__inst_mult_24_350 ;
wire Xd_0__inst_mult_24_354 ;
wire Xd_0__inst_mult_24_355 ;
wire Xd_0__inst_mult_26_339 ;
wire Xd_0__inst_mult_26_340 ;
wire Xd_0__inst_mult_26_344 ;
wire Xd_0__inst_mult_26_345 ;
wire Xd_0__inst_mult_26_349 ;
wire Xd_0__inst_mult_26_350 ;
wire Xd_0__inst_mult_26_354 ;
wire Xd_0__inst_mult_26_355 ;
wire Xd_0__inst_mult_26_359 ;
wire Xd_0__inst_mult_26_360 ;
wire Xd_0__inst_a1_7__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_6__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_19_210 ;
wire Xd_0__inst_mult_19_35_sumout ;
wire Xd_0__inst_mult_19_36 ;
wire Xd_0__inst_mult_19_214 ;
wire Xd_0__inst_mult_19_215 ;
wire Xd_0__inst_a1_5__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_4__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_17_210 ;
wire Xd_0__inst_mult_17_35_sumout ;
wire Xd_0__inst_mult_17_36 ;
wire Xd_0__inst_mult_17_214 ;
wire Xd_0__inst_mult_17_215 ;
wire Xd_0__inst_mult_27_249 ;
wire Xd_0__inst_mult_27_250 ;
wire Xd_0__inst_mult_27_254 ;
wire Xd_0__inst_mult_27_255 ;
wire Xd_0__inst_mult_27_259 ;
wire Xd_0__inst_mult_27_260 ;
wire Xd_0__inst_mult_27_264 ;
wire Xd_0__inst_mult_27_265 ;
wire Xd_0__inst_a1_3__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_2__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_16_210 ;
wire Xd_0__inst_mult_16_35_sumout ;
wire Xd_0__inst_mult_16_36 ;
wire Xd_0__inst_mult_16_214 ;
wire Xd_0__inst_mult_16_215 ;
wire Xd_0__inst_a1_1__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_a1_0__adder1_inst_add_0_122_cout ;
wire Xd_0__inst_mult_29_210 ;
wire Xd_0__inst_mult_29_35_sumout ;
wire Xd_0__inst_mult_29_36 ;
wire Xd_0__inst_mult_29_214 ;
wire Xd_0__inst_mult_29_215 ;
wire Xd_0__inst_mult_26_364 ;
wire Xd_0__inst_mult_26_365 ;
wire Xd_0__inst_mult_26_369 ;
wire Xd_0__inst_mult_26_370 ;
wire Xd_0__inst_mult_26_374 ;
wire Xd_0__inst_mult_26_375 ;
wire Xd_0__inst_mult_26_379 ;
wire Xd_0__inst_mult_26_380 ;
wire Xd_0__inst_mult_24_359 ;
wire Xd_0__inst_mult_24_360 ;
wire Xd_0__inst_mult_24_364 ;
wire Xd_0__inst_mult_24_365 ;
wire Xd_0__inst_mult_24_369 ;
wire Xd_0__inst_mult_24_370 ;
wire Xd_0__inst_mult_24_374 ;
wire Xd_0__inst_mult_24_375 ;
wire Xd_0__inst_mult_24_379 ;
wire Xd_0__inst_mult_24_380 ;
wire Xd_0__inst_mult_2_244 ;
wire Xd_0__inst_mult_2_245 ;
wire Xd_0__inst_mult_9_205 ;
wire Xd_0__inst_mult_9_206 ;
wire Xd_0__inst_mult_8_205 ;
wire Xd_0__inst_mult_8_206 ;
wire Xd_0__inst_i29_1_sumout ;
wire Xd_0__inst_i29_2 ;
wire Xd_0__inst_mult_21_219 ;
wire Xd_0__inst_mult_21_220 ;
wire Xd_0__inst_mult_13_35_sumout ;
wire Xd_0__inst_mult_13_36 ;
wire Xd_0__inst_mult_21_40_sumout ;
wire Xd_0__inst_mult_21_41 ;
wire Xd_0__inst_mult_21_224 ;
wire Xd_0__inst_mult_21_225 ;
wire Xd_0__inst_mult_11_205 ;
wire Xd_0__inst_mult_11_206 ;
wire Xd_0__inst_mult_10_205 ;
wire Xd_0__inst_mult_10_206 ;
wire Xd_0__inst_i29_6_sumout ;
wire Xd_0__inst_i29_7 ;
wire Xd_0__inst_mult_20_219 ;
wire Xd_0__inst_mult_20_220 ;
wire Xd_0__inst_mult_20_40_sumout ;
wire Xd_0__inst_mult_20_41 ;
wire Xd_0__inst_mult_20_45_sumout ;
wire Xd_0__inst_mult_20_46 ;
wire Xd_0__inst_mult_20_224 ;
wire Xd_0__inst_mult_20_225 ;
wire Xd_0__inst_mult_25_269 ;
wire Xd_0__inst_mult_25_270 ;
wire Xd_0__inst_mult_25_274 ;
wire Xd_0__inst_mult_25_275 ;
wire Xd_0__inst_mult_25_279 ;
wire Xd_0__inst_mult_25_280 ;
wire Xd_0__inst_mult_25_284 ;
wire Xd_0__inst_mult_25_285 ;
wire Xd_0__inst_mult_3_205 ;
wire Xd_0__inst_mult_3_206 ;
wire Xd_0__inst_mult_0_205 ;
wire Xd_0__inst_mult_0_206 ;
wire Xd_0__inst_i29_11_sumout ;
wire Xd_0__inst_i29_12 ;
wire Xd_0__inst_mult_23_219 ;
wire Xd_0__inst_mult_23_220 ;
wire Xd_0__inst_mult_23_40_sumout ;
wire Xd_0__inst_mult_23_41 ;
wire Xd_0__inst_mult_23_224 ;
wire Xd_0__inst_mult_23_225 ;
wire Xd_0__inst_mult_6_205 ;
wire Xd_0__inst_mult_6_206 ;
wire Xd_0__inst_mult_1_205 ;
wire Xd_0__inst_mult_1_206 ;
wire Xd_0__inst_i29_16_sumout ;
wire Xd_0__inst_i29_17 ;
wire Xd_0__inst_mult_22_219 ;
wire Xd_0__inst_mult_22_220 ;
wire Xd_0__inst_mult_22_40_sumout ;
wire Xd_0__inst_mult_22_41 ;
wire Xd_0__inst_mult_22_224 ;
wire Xd_0__inst_mult_22_225 ;
wire Xd_0__inst_mult_24_384 ;
wire Xd_0__inst_mult_24_385 ;
wire Xd_0__inst_mult_24_389 ;
wire Xd_0__inst_mult_24_390 ;
wire Xd_0__inst_mult_24_394 ;
wire Xd_0__inst_mult_24_395 ;
wire Xd_0__inst_mult_24_399 ;
wire Xd_0__inst_mult_24_400 ;
wire Xd_0__inst_mult_26_384 ;
wire Xd_0__inst_mult_26_385 ;
wire Xd_0__inst_mult_26_389 ;
wire Xd_0__inst_mult_26_390 ;
wire Xd_0__inst_mult_26_394 ;
wire Xd_0__inst_mult_26_395 ;
wire Xd_0__inst_mult_26_399 ;
wire Xd_0__inst_mult_26_400 ;
wire Xd_0__inst_mult_26_404 ;
wire Xd_0__inst_mult_26_405 ;
wire Xd_0__inst_mult_7_205 ;
wire Xd_0__inst_mult_7_206 ;
wire Xd_0__inst_mult_4_205 ;
wire Xd_0__inst_mult_4_206 ;
wire Xd_0__inst_i29_21_sumout ;
wire Xd_0__inst_i29_22 ;
wire Xd_0__inst_mult_19_219 ;
wire Xd_0__inst_mult_19_220 ;
wire Xd_0__inst_mult_19_40_sumout ;
wire Xd_0__inst_mult_19_41 ;
wire Xd_0__inst_mult_19_224 ;
wire Xd_0__inst_mult_19_225 ;
wire Xd_0__inst_mult_30_205 ;
wire Xd_0__inst_mult_30_206 ;
wire Xd_0__inst_mult_5_205 ;
wire Xd_0__inst_mult_5_206 ;
wire Xd_0__inst_i29_26_sumout ;
wire Xd_0__inst_i29_27 ;
wire Xd_0__inst_mult_17_219 ;
wire Xd_0__inst_mult_17_220 ;
wire Xd_0__inst_mult_17_40_sumout ;
wire Xd_0__inst_mult_17_41 ;
wire Xd_0__inst_mult_17_224 ;
wire Xd_0__inst_mult_17_225 ;
wire Xd_0__inst_mult_27_269 ;
wire Xd_0__inst_mult_27_270 ;
wire Xd_0__inst_mult_27_274 ;
wire Xd_0__inst_mult_27_275 ;
wire Xd_0__inst_mult_27_279 ;
wire Xd_0__inst_mult_27_280 ;
wire Xd_0__inst_mult_27_284 ;
wire Xd_0__inst_mult_27_285 ;
wire Xd_0__inst_mult_13_205 ;
wire Xd_0__inst_mult_13_206 ;
wire Xd_0__inst_mult_2_249 ;
wire Xd_0__inst_mult_2_250 ;
wire Xd_0__inst_i29_31_sumout ;
wire Xd_0__inst_i29_32 ;
wire Xd_0__inst_mult_16_219 ;
wire Xd_0__inst_mult_16_220 ;
wire Xd_0__inst_mult_16_40_sumout ;
wire Xd_0__inst_mult_16_41 ;
wire Xd_0__inst_mult_16_224 ;
wire Xd_0__inst_mult_16_225 ;
wire Xd_0__inst_mult_28_205 ;
wire Xd_0__inst_mult_28_206 ;
wire Xd_0__inst_mult_31_205 ;
wire Xd_0__inst_mult_31_206 ;
wire Xd_0__inst_i29_36_sumout ;
wire Xd_0__inst_i29_37 ;
wire Xd_0__inst_mult_29_219 ;
wire Xd_0__inst_mult_29_220 ;
wire Xd_0__inst_mult_29_40_sumout ;
wire Xd_0__inst_mult_29_41 ;
wire Xd_0__inst_mult_29_224 ;
wire Xd_0__inst_mult_29_225 ;
wire Xd_0__inst_mult_26_409 ;
wire Xd_0__inst_mult_26_410 ;
wire Xd_0__inst_mult_26_414 ;
wire Xd_0__inst_mult_26_415 ;
wire Xd_0__inst_mult_26_419 ;
wire Xd_0__inst_mult_26_420 ;
wire Xd_0__inst_mult_26_424 ;
wire Xd_0__inst_mult_26_425 ;
wire Xd_0__inst_mult_24_404 ;
wire Xd_0__inst_mult_24_405 ;
wire Xd_0__inst_mult_24_409 ;
wire Xd_0__inst_mult_24_410 ;
wire Xd_0__inst_mult_24_414 ;
wire Xd_0__inst_mult_24_415 ;
wire Xd_0__inst_mult_24_419 ;
wire Xd_0__inst_mult_24_420 ;
wire Xd_0__inst_mult_24_424 ;
wire Xd_0__inst_mult_24_425 ;
wire Xd_0__inst_mult_2_254 ;
wire Xd_0__inst_mult_2_255 ;
wire Xd_0__inst_mult_29_229 ;
wire Xd_0__inst_mult_29_230 ;
wire Xd_0__inst_mult_28_210 ;
wire Xd_0__inst_mult_28_211 ;
wire Xd_0__inst_mult_31_210 ;
wire Xd_0__inst_mult_31_211 ;
wire Xd_0__inst_mult_30_210 ;
wire Xd_0__inst_mult_30_211 ;
wire Xd_0__inst_mult_25_289 ;
wire Xd_0__inst_mult_25_290 ;
wire Xd_0__inst_mult_24_429 ;
wire Xd_0__inst_mult_24_430 ;
wire Xd_0__inst_mult_27_289 ;
wire Xd_0__inst_mult_27_290 ;
wire Xd_0__inst_mult_26_429 ;
wire Xd_0__inst_mult_26_430 ;
wire Xd_0__inst_mult_21_229 ;
wire Xd_0__inst_mult_21_230 ;
wire Xd_0__inst_mult_20_229 ;
wire Xd_0__inst_mult_20_230 ;
wire Xd_0__inst_mult_23_229 ;
wire Xd_0__inst_mult_23_230 ;
wire Xd_0__inst_mult_22_229 ;
wire Xd_0__inst_mult_22_230 ;
wire Xd_0__inst_mult_17_229 ;
wire Xd_0__inst_mult_17_230 ;
wire Xd_0__inst_mult_16_229 ;
wire Xd_0__inst_mult_16_230 ;
wire Xd_0__inst_mult_19_229 ;
wire Xd_0__inst_mult_19_230 ;
wire Xd_0__inst_mult_18_205 ;
wire Xd_0__inst_mult_18_206 ;
wire Xd_0__inst_mult_13_210 ;
wire Xd_0__inst_mult_13_211 ;
wire Xd_0__inst_mult_12_205 ;
wire Xd_0__inst_mult_12_206 ;
wire Xd_0__inst_mult_15_205 ;
wire Xd_0__inst_mult_15_206 ;
wire Xd_0__inst_mult_14_205 ;
wire Xd_0__inst_mult_14_206 ;
wire Xd_0__inst_mult_9_210 ;
wire Xd_0__inst_mult_9_211 ;
wire Xd_0__inst_mult_8_210 ;
wire Xd_0__inst_mult_8_211 ;
wire Xd_0__inst_mult_11_210 ;
wire Xd_0__inst_mult_11_211 ;
wire Xd_0__inst_mult_10_210 ;
wire Xd_0__inst_mult_10_211 ;
wire Xd_0__inst_mult_5_210 ;
wire Xd_0__inst_mult_5_211 ;
wire Xd_0__inst_mult_4_210 ;
wire Xd_0__inst_mult_4_211 ;
wire Xd_0__inst_mult_7_210 ;
wire Xd_0__inst_mult_7_211 ;
wire Xd_0__inst_mult_6_210 ;
wire Xd_0__inst_mult_6_211 ;
wire Xd_0__inst_mult_1_210 ;
wire Xd_0__inst_mult_1_211 ;
wire Xd_0__inst_mult_0_210 ;
wire Xd_0__inst_mult_0_211 ;
wire Xd_0__inst_mult_3_210 ;
wire Xd_0__inst_mult_3_211 ;
wire Xd_0__inst_mult_2_259 ;
wire Xd_0__inst_mult_2_260 ;
wire Xd_0__inst_mult_29_234 ;
wire Xd_0__inst_mult_29_235 ;
wire Xd_0__inst_mult_28_214 ;
wire Xd_0__inst_mult_28_215 ;
wire Xd_0__inst_mult_31_214 ;
wire Xd_0__inst_mult_31_215 ;
wire Xd_0__inst_mult_30_214 ;
wire Xd_0__inst_mult_30_215 ;
wire Xd_0__inst_mult_25_294 ;
wire Xd_0__inst_mult_25_295 ;
wire Xd_0__inst_mult_24_434 ;
wire Xd_0__inst_mult_24_435 ;
wire Xd_0__inst_mult_27_294 ;
wire Xd_0__inst_mult_27_295 ;
wire Xd_0__inst_mult_26_434 ;
wire Xd_0__inst_mult_26_435 ;
wire Xd_0__inst_mult_21_234 ;
wire Xd_0__inst_mult_21_235 ;
wire Xd_0__inst_mult_20_234 ;
wire Xd_0__inst_mult_20_235 ;
wire Xd_0__inst_mult_23_234 ;
wire Xd_0__inst_mult_23_235 ;
wire Xd_0__inst_mult_22_234 ;
wire Xd_0__inst_mult_22_235 ;
wire Xd_0__inst_mult_17_234 ;
wire Xd_0__inst_mult_17_235 ;
wire Xd_0__inst_mult_16_234 ;
wire Xd_0__inst_mult_16_235 ;
wire Xd_0__inst_mult_19_234 ;
wire Xd_0__inst_mult_19_235 ;
wire Xd_0__inst_mult_18_210 ;
wire Xd_0__inst_mult_18_211 ;
wire Xd_0__inst_mult_13_214 ;
wire Xd_0__inst_mult_13_215 ;
wire Xd_0__inst_mult_12_210 ;
wire Xd_0__inst_mult_12_211 ;
wire Xd_0__inst_mult_15_210 ;
wire Xd_0__inst_mult_15_211 ;
wire Xd_0__inst_mult_14_210 ;
wire Xd_0__inst_mult_14_211 ;
wire Xd_0__inst_mult_9_214 ;
wire Xd_0__inst_mult_9_215 ;
wire Xd_0__inst_mult_8_214 ;
wire Xd_0__inst_mult_8_215 ;
wire Xd_0__inst_mult_11_214 ;
wire Xd_0__inst_mult_11_215 ;
wire Xd_0__inst_mult_10_214 ;
wire Xd_0__inst_mult_10_215 ;
wire Xd_0__inst_mult_5_214 ;
wire Xd_0__inst_mult_5_215 ;
wire Xd_0__inst_mult_4_214 ;
wire Xd_0__inst_mult_4_215 ;
wire Xd_0__inst_mult_7_214 ;
wire Xd_0__inst_mult_7_215 ;
wire Xd_0__inst_mult_6_214 ;
wire Xd_0__inst_mult_6_215 ;
wire Xd_0__inst_mult_1_214 ;
wire Xd_0__inst_mult_1_215 ;
wire Xd_0__inst_mult_0_214 ;
wire Xd_0__inst_mult_0_215 ;
wire Xd_0__inst_mult_3_214 ;
wire Xd_0__inst_mult_3_215 ;
wire Xd_0__inst_mult_2_264 ;
wire Xd_0__inst_mult_2_265 ;
wire Xd_0__inst_mult_29_239 ;
wire Xd_0__inst_mult_29_240 ;
wire Xd_0__inst_mult_28_219 ;
wire Xd_0__inst_mult_28_220 ;
wire Xd_0__inst_mult_31_219 ;
wire Xd_0__inst_mult_31_220 ;
wire Xd_0__inst_mult_30_219 ;
wire Xd_0__inst_mult_30_220 ;
wire Xd_0__inst_mult_25_299 ;
wire Xd_0__inst_mult_25_300 ;
wire Xd_0__inst_mult_24_439 ;
wire Xd_0__inst_mult_24_440 ;
wire Xd_0__inst_mult_27_299 ;
wire Xd_0__inst_mult_27_300 ;
wire Xd_0__inst_mult_26_439 ;
wire Xd_0__inst_mult_26_440 ;
wire Xd_0__inst_mult_21_239 ;
wire Xd_0__inst_mult_21_240 ;
wire Xd_0__inst_mult_20_239 ;
wire Xd_0__inst_mult_20_240 ;
wire Xd_0__inst_mult_23_239 ;
wire Xd_0__inst_mult_23_240 ;
wire Xd_0__inst_mult_22_239 ;
wire Xd_0__inst_mult_22_240 ;
wire Xd_0__inst_mult_17_239 ;
wire Xd_0__inst_mult_17_240 ;
wire Xd_0__inst_mult_16_239 ;
wire Xd_0__inst_mult_16_240 ;
wire Xd_0__inst_mult_19_239 ;
wire Xd_0__inst_mult_19_240 ;
wire Xd_0__inst_mult_18_214 ;
wire Xd_0__inst_mult_18_215 ;
wire Xd_0__inst_mult_13_219 ;
wire Xd_0__inst_mult_13_220 ;
wire Xd_0__inst_mult_12_214 ;
wire Xd_0__inst_mult_12_215 ;
wire Xd_0__inst_mult_15_214 ;
wire Xd_0__inst_mult_15_215 ;
wire Xd_0__inst_mult_14_214 ;
wire Xd_0__inst_mult_14_215 ;
wire Xd_0__inst_mult_9_219 ;
wire Xd_0__inst_mult_9_220 ;
wire Xd_0__inst_mult_8_219 ;
wire Xd_0__inst_mult_8_220 ;
wire Xd_0__inst_mult_11_219 ;
wire Xd_0__inst_mult_11_220 ;
wire Xd_0__inst_mult_10_219 ;
wire Xd_0__inst_mult_10_220 ;
wire Xd_0__inst_mult_5_219 ;
wire Xd_0__inst_mult_5_220 ;
wire Xd_0__inst_mult_4_219 ;
wire Xd_0__inst_mult_4_220 ;
wire Xd_0__inst_mult_7_219 ;
wire Xd_0__inst_mult_7_220 ;
wire Xd_0__inst_mult_6_219 ;
wire Xd_0__inst_mult_6_220 ;
wire Xd_0__inst_mult_1_219 ;
wire Xd_0__inst_mult_1_220 ;
wire Xd_0__inst_mult_0_219 ;
wire Xd_0__inst_mult_0_220 ;
wire Xd_0__inst_mult_3_219 ;
wire Xd_0__inst_mult_3_220 ;
wire Xd_0__inst_mult_2_269 ;
wire Xd_0__inst_mult_2_270 ;
wire Xd_0__inst_mult_29_244 ;
wire Xd_0__inst_mult_29_245 ;
wire Xd_0__inst_mult_28_224 ;
wire Xd_0__inst_mult_28_225 ;
wire Xd_0__inst_mult_31_224 ;
wire Xd_0__inst_mult_31_225 ;
wire Xd_0__inst_mult_30_224 ;
wire Xd_0__inst_mult_30_225 ;
wire Xd_0__inst_mult_25_304 ;
wire Xd_0__inst_mult_25_305 ;
wire Xd_0__inst_mult_24_444 ;
wire Xd_0__inst_mult_24_445 ;
wire Xd_0__inst_mult_27_304 ;
wire Xd_0__inst_mult_27_305 ;
wire Xd_0__inst_mult_26_444 ;
wire Xd_0__inst_mult_26_445 ;
wire Xd_0__inst_mult_21_244 ;
wire Xd_0__inst_mult_21_245 ;
wire Xd_0__inst_mult_20_244 ;
wire Xd_0__inst_mult_20_245 ;
wire Xd_0__inst_mult_23_244 ;
wire Xd_0__inst_mult_23_245 ;
wire Xd_0__inst_mult_22_244 ;
wire Xd_0__inst_mult_22_245 ;
wire Xd_0__inst_mult_17_244 ;
wire Xd_0__inst_mult_17_245 ;
wire Xd_0__inst_mult_16_244 ;
wire Xd_0__inst_mult_16_245 ;
wire Xd_0__inst_mult_19_244 ;
wire Xd_0__inst_mult_19_245 ;
wire Xd_0__inst_mult_18_219 ;
wire Xd_0__inst_mult_18_220 ;
wire Xd_0__inst_mult_13_224 ;
wire Xd_0__inst_mult_13_225 ;
wire Xd_0__inst_mult_12_219 ;
wire Xd_0__inst_mult_12_220 ;
wire Xd_0__inst_mult_15_219 ;
wire Xd_0__inst_mult_15_220 ;
wire Xd_0__inst_mult_14_219 ;
wire Xd_0__inst_mult_14_220 ;
wire Xd_0__inst_mult_9_224 ;
wire Xd_0__inst_mult_9_225 ;
wire Xd_0__inst_mult_8_224 ;
wire Xd_0__inst_mult_8_225 ;
wire Xd_0__inst_mult_11_224 ;
wire Xd_0__inst_mult_11_225 ;
wire Xd_0__inst_mult_10_224 ;
wire Xd_0__inst_mult_10_225 ;
wire Xd_0__inst_mult_5_224 ;
wire Xd_0__inst_mult_5_225 ;
wire Xd_0__inst_mult_4_224 ;
wire Xd_0__inst_mult_4_225 ;
wire Xd_0__inst_mult_7_224 ;
wire Xd_0__inst_mult_7_225 ;
wire Xd_0__inst_mult_6_224 ;
wire Xd_0__inst_mult_6_225 ;
wire Xd_0__inst_mult_1_224 ;
wire Xd_0__inst_mult_1_225 ;
wire Xd_0__inst_mult_0_224 ;
wire Xd_0__inst_mult_0_225 ;
wire Xd_0__inst_mult_3_224 ;
wire Xd_0__inst_mult_3_225 ;
wire Xd_0__inst_mult_2_274 ;
wire Xd_0__inst_mult_2_275 ;
wire Xd_0__inst_mult_29_249 ;
wire Xd_0__inst_mult_29_250 ;
wire Xd_0__inst_mult_28_229 ;
wire Xd_0__inst_mult_28_230 ;
wire Xd_0__inst_mult_31_229 ;
wire Xd_0__inst_mult_31_230 ;
wire Xd_0__inst_mult_30_229 ;
wire Xd_0__inst_mult_30_230 ;
wire Xd_0__inst_mult_25_309 ;
wire Xd_0__inst_mult_25_310 ;
wire Xd_0__inst_mult_24_449 ;
wire Xd_0__inst_mult_24_450 ;
wire Xd_0__inst_mult_27_309 ;
wire Xd_0__inst_mult_27_310 ;
wire Xd_0__inst_mult_26_449 ;
wire Xd_0__inst_mult_26_450 ;
wire Xd_0__inst_mult_21_249 ;
wire Xd_0__inst_mult_21_250 ;
wire Xd_0__inst_mult_20_249 ;
wire Xd_0__inst_mult_20_250 ;
wire Xd_0__inst_mult_23_249 ;
wire Xd_0__inst_mult_23_250 ;
wire Xd_0__inst_mult_22_249 ;
wire Xd_0__inst_mult_22_250 ;
wire Xd_0__inst_mult_17_249 ;
wire Xd_0__inst_mult_17_250 ;
wire Xd_0__inst_mult_16_249 ;
wire Xd_0__inst_mult_16_250 ;
wire Xd_0__inst_mult_19_249 ;
wire Xd_0__inst_mult_19_250 ;
wire Xd_0__inst_mult_18_224 ;
wire Xd_0__inst_mult_18_225 ;
wire Xd_0__inst_mult_13_229 ;
wire Xd_0__inst_mult_13_230 ;
wire Xd_0__inst_mult_12_224 ;
wire Xd_0__inst_mult_12_225 ;
wire Xd_0__inst_mult_15_224 ;
wire Xd_0__inst_mult_15_225 ;
wire Xd_0__inst_mult_14_224 ;
wire Xd_0__inst_mult_14_225 ;
wire Xd_0__inst_mult_9_229 ;
wire Xd_0__inst_mult_9_230 ;
wire Xd_0__inst_mult_8_229 ;
wire Xd_0__inst_mult_8_230 ;
wire Xd_0__inst_mult_11_229 ;
wire Xd_0__inst_mult_11_230 ;
wire Xd_0__inst_mult_10_229 ;
wire Xd_0__inst_mult_10_230 ;
wire Xd_0__inst_mult_5_229 ;
wire Xd_0__inst_mult_5_230 ;
wire Xd_0__inst_mult_4_229 ;
wire Xd_0__inst_mult_4_230 ;
wire Xd_0__inst_mult_7_229 ;
wire Xd_0__inst_mult_7_230 ;
wire Xd_0__inst_mult_6_229 ;
wire Xd_0__inst_mult_6_230 ;
wire Xd_0__inst_mult_1_229 ;
wire Xd_0__inst_mult_1_230 ;
wire Xd_0__inst_mult_0_229 ;
wire Xd_0__inst_mult_0_230 ;
wire Xd_0__inst_mult_3_229 ;
wire Xd_0__inst_mult_3_230 ;
wire Xd_0__inst_mult_2_279 ;
wire Xd_0__inst_mult_2_280 ;
wire Xd_0__inst_mult_29_254 ;
wire Xd_0__inst_mult_29_255 ;
wire Xd_0__inst_mult_28_234 ;
wire Xd_0__inst_mult_28_235 ;
wire Xd_0__inst_mult_31_234 ;
wire Xd_0__inst_mult_31_235 ;
wire Xd_0__inst_mult_30_234 ;
wire Xd_0__inst_mult_30_235 ;
wire Xd_0__inst_mult_25_314 ;
wire Xd_0__inst_mult_25_315 ;
wire Xd_0__inst_mult_24_454 ;
wire Xd_0__inst_mult_24_455 ;
wire Xd_0__inst_mult_27_314 ;
wire Xd_0__inst_mult_27_315 ;
wire Xd_0__inst_mult_26_454 ;
wire Xd_0__inst_mult_26_455 ;
wire Xd_0__inst_mult_21_254 ;
wire Xd_0__inst_mult_21_255 ;
wire Xd_0__inst_mult_20_254 ;
wire Xd_0__inst_mult_20_255 ;
wire Xd_0__inst_mult_23_254 ;
wire Xd_0__inst_mult_23_255 ;
wire Xd_0__inst_mult_22_254 ;
wire Xd_0__inst_mult_22_255 ;
wire Xd_0__inst_mult_17_254 ;
wire Xd_0__inst_mult_17_255 ;
wire Xd_0__inst_mult_16_254 ;
wire Xd_0__inst_mult_16_255 ;
wire Xd_0__inst_mult_19_254 ;
wire Xd_0__inst_mult_19_255 ;
wire Xd_0__inst_mult_18_229 ;
wire Xd_0__inst_mult_18_230 ;
wire Xd_0__inst_mult_13_234 ;
wire Xd_0__inst_mult_13_235 ;
wire Xd_0__inst_mult_12_229 ;
wire Xd_0__inst_mult_12_230 ;
wire Xd_0__inst_mult_15_229 ;
wire Xd_0__inst_mult_15_230 ;
wire Xd_0__inst_mult_14_229 ;
wire Xd_0__inst_mult_14_230 ;
wire Xd_0__inst_mult_9_234 ;
wire Xd_0__inst_mult_9_235 ;
wire Xd_0__inst_mult_8_234 ;
wire Xd_0__inst_mult_8_235 ;
wire Xd_0__inst_mult_11_234 ;
wire Xd_0__inst_mult_11_235 ;
wire Xd_0__inst_mult_10_234 ;
wire Xd_0__inst_mult_10_235 ;
wire Xd_0__inst_mult_5_234 ;
wire Xd_0__inst_mult_5_235 ;
wire Xd_0__inst_mult_4_234 ;
wire Xd_0__inst_mult_4_235 ;
wire Xd_0__inst_mult_7_234 ;
wire Xd_0__inst_mult_7_235 ;
wire Xd_0__inst_mult_6_234 ;
wire Xd_0__inst_mult_6_235 ;
wire Xd_0__inst_mult_1_234 ;
wire Xd_0__inst_mult_1_235 ;
wire Xd_0__inst_mult_0_234 ;
wire Xd_0__inst_mult_0_235 ;
wire Xd_0__inst_mult_3_234 ;
wire Xd_0__inst_mult_3_235 ;
wire Xd_0__inst_mult_2_284 ;
wire Xd_0__inst_mult_2_285 ;
wire Xd_0__inst_mult_29_259 ;
wire Xd_0__inst_mult_29_260 ;
wire Xd_0__inst_mult_28_239 ;
wire Xd_0__inst_mult_28_240 ;
wire Xd_0__inst_mult_31_239 ;
wire Xd_0__inst_mult_31_240 ;
wire Xd_0__inst_mult_30_239 ;
wire Xd_0__inst_mult_30_240 ;
wire Xd_0__inst_mult_25_319 ;
wire Xd_0__inst_mult_25_320 ;
wire Xd_0__inst_mult_24_459 ;
wire Xd_0__inst_mult_24_460 ;
wire Xd_0__inst_mult_27_319 ;
wire Xd_0__inst_mult_27_320 ;
wire Xd_0__inst_mult_26_459 ;
wire Xd_0__inst_mult_26_460 ;
wire Xd_0__inst_mult_21_259 ;
wire Xd_0__inst_mult_21_260 ;
wire Xd_0__inst_mult_20_259 ;
wire Xd_0__inst_mult_20_260 ;
wire Xd_0__inst_mult_23_259 ;
wire Xd_0__inst_mult_23_260 ;
wire Xd_0__inst_mult_22_259 ;
wire Xd_0__inst_mult_22_260 ;
wire Xd_0__inst_mult_17_259 ;
wire Xd_0__inst_mult_17_260 ;
wire Xd_0__inst_mult_16_259 ;
wire Xd_0__inst_mult_16_260 ;
wire Xd_0__inst_mult_19_259 ;
wire Xd_0__inst_mult_19_260 ;
wire Xd_0__inst_mult_18_234 ;
wire Xd_0__inst_mult_18_235 ;
wire Xd_0__inst_mult_13_239 ;
wire Xd_0__inst_mult_13_240 ;
wire Xd_0__inst_mult_12_234 ;
wire Xd_0__inst_mult_12_235 ;
wire Xd_0__inst_mult_15_234 ;
wire Xd_0__inst_mult_15_235 ;
wire Xd_0__inst_mult_14_234 ;
wire Xd_0__inst_mult_14_235 ;
wire Xd_0__inst_mult_9_239 ;
wire Xd_0__inst_mult_9_240 ;
wire Xd_0__inst_mult_8_239 ;
wire Xd_0__inst_mult_8_240 ;
wire Xd_0__inst_mult_11_239 ;
wire Xd_0__inst_mult_11_240 ;
wire Xd_0__inst_mult_10_239 ;
wire Xd_0__inst_mult_10_240 ;
wire Xd_0__inst_mult_5_239 ;
wire Xd_0__inst_mult_5_240 ;
wire Xd_0__inst_mult_4_239 ;
wire Xd_0__inst_mult_4_240 ;
wire Xd_0__inst_mult_7_239 ;
wire Xd_0__inst_mult_7_240 ;
wire Xd_0__inst_mult_6_239 ;
wire Xd_0__inst_mult_6_240 ;
wire Xd_0__inst_mult_1_239 ;
wire Xd_0__inst_mult_1_240 ;
wire Xd_0__inst_mult_0_239 ;
wire Xd_0__inst_mult_0_240 ;
wire Xd_0__inst_mult_3_239 ;
wire Xd_0__inst_mult_3_240 ;
wire Xd_0__inst_mult_2_289 ;
wire Xd_0__inst_mult_2_290 ;
wire Xd_0__inst_mult_29_264 ;
wire Xd_0__inst_mult_29_265 ;
wire Xd_0__inst_mult_28_244 ;
wire Xd_0__inst_mult_28_245 ;
wire Xd_0__inst_mult_31_244 ;
wire Xd_0__inst_mult_31_245 ;
wire Xd_0__inst_mult_30_244 ;
wire Xd_0__inst_mult_30_245 ;
wire Xd_0__inst_mult_25_324 ;
wire Xd_0__inst_mult_25_325 ;
wire Xd_0__inst_mult_24_464 ;
wire Xd_0__inst_mult_24_465 ;
wire Xd_0__inst_mult_27_324 ;
wire Xd_0__inst_mult_27_325 ;
wire Xd_0__inst_mult_26_464 ;
wire Xd_0__inst_mult_26_465 ;
wire Xd_0__inst_mult_21_264 ;
wire Xd_0__inst_mult_21_265 ;
wire Xd_0__inst_mult_20_264 ;
wire Xd_0__inst_mult_20_265 ;
wire Xd_0__inst_mult_23_264 ;
wire Xd_0__inst_mult_23_265 ;
wire Xd_0__inst_mult_22_264 ;
wire Xd_0__inst_mult_22_265 ;
wire Xd_0__inst_mult_17_264 ;
wire Xd_0__inst_mult_17_265 ;
wire Xd_0__inst_mult_16_264 ;
wire Xd_0__inst_mult_16_265 ;
wire Xd_0__inst_mult_19_264 ;
wire Xd_0__inst_mult_19_265 ;
wire Xd_0__inst_mult_18_239 ;
wire Xd_0__inst_mult_18_240 ;
wire Xd_0__inst_mult_13_244 ;
wire Xd_0__inst_mult_13_245 ;
wire Xd_0__inst_mult_12_239 ;
wire Xd_0__inst_mult_12_240 ;
wire Xd_0__inst_mult_15_239 ;
wire Xd_0__inst_mult_15_240 ;
wire Xd_0__inst_mult_14_239 ;
wire Xd_0__inst_mult_14_240 ;
wire Xd_0__inst_mult_9_244 ;
wire Xd_0__inst_mult_9_245 ;
wire Xd_0__inst_mult_8_244 ;
wire Xd_0__inst_mult_8_245 ;
wire Xd_0__inst_mult_11_244 ;
wire Xd_0__inst_mult_11_245 ;
wire Xd_0__inst_mult_10_244 ;
wire Xd_0__inst_mult_10_245 ;
wire Xd_0__inst_mult_5_244 ;
wire Xd_0__inst_mult_5_245 ;
wire Xd_0__inst_mult_4_244 ;
wire Xd_0__inst_mult_4_245 ;
wire Xd_0__inst_mult_7_244 ;
wire Xd_0__inst_mult_7_245 ;
wire Xd_0__inst_mult_6_244 ;
wire Xd_0__inst_mult_6_245 ;
wire Xd_0__inst_mult_1_244 ;
wire Xd_0__inst_mult_1_245 ;
wire Xd_0__inst_mult_0_244 ;
wire Xd_0__inst_mult_0_245 ;
wire Xd_0__inst_mult_3_244 ;
wire Xd_0__inst_mult_3_245 ;
wire Xd_0__inst_mult_2_294 ;
wire Xd_0__inst_mult_2_295 ;
wire Xd_0__inst_mult_29_269 ;
wire Xd_0__inst_mult_29_270 ;
wire Xd_0__inst_mult_28_249 ;
wire Xd_0__inst_mult_28_250 ;
wire Xd_0__inst_mult_31_249 ;
wire Xd_0__inst_mult_31_250 ;
wire Xd_0__inst_mult_30_249 ;
wire Xd_0__inst_mult_30_250 ;
wire Xd_0__inst_mult_25_329 ;
wire Xd_0__inst_mult_25_330 ;
wire Xd_0__inst_mult_24_469 ;
wire Xd_0__inst_mult_24_470 ;
wire Xd_0__inst_mult_27_329 ;
wire Xd_0__inst_mult_27_330 ;
wire Xd_0__inst_mult_26_469 ;
wire Xd_0__inst_mult_26_470 ;
wire Xd_0__inst_mult_21_269 ;
wire Xd_0__inst_mult_21_270 ;
wire Xd_0__inst_mult_20_269 ;
wire Xd_0__inst_mult_20_270 ;
wire Xd_0__inst_mult_23_269 ;
wire Xd_0__inst_mult_23_270 ;
wire Xd_0__inst_mult_22_269 ;
wire Xd_0__inst_mult_22_270 ;
wire Xd_0__inst_mult_17_269 ;
wire Xd_0__inst_mult_17_270 ;
wire Xd_0__inst_mult_16_269 ;
wire Xd_0__inst_mult_16_270 ;
wire Xd_0__inst_mult_19_269 ;
wire Xd_0__inst_mult_19_270 ;
wire Xd_0__inst_mult_18_244 ;
wire Xd_0__inst_mult_18_245 ;
wire Xd_0__inst_mult_13_249 ;
wire Xd_0__inst_mult_13_250 ;
wire Xd_0__inst_mult_12_244 ;
wire Xd_0__inst_mult_12_245 ;
wire Xd_0__inst_mult_15_244 ;
wire Xd_0__inst_mult_15_245 ;
wire Xd_0__inst_mult_14_244 ;
wire Xd_0__inst_mult_14_245 ;
wire Xd_0__inst_mult_9_249 ;
wire Xd_0__inst_mult_9_250 ;
wire Xd_0__inst_mult_8_249 ;
wire Xd_0__inst_mult_8_250 ;
wire Xd_0__inst_mult_11_249 ;
wire Xd_0__inst_mult_11_250 ;
wire Xd_0__inst_mult_10_249 ;
wire Xd_0__inst_mult_10_250 ;
wire Xd_0__inst_mult_5_249 ;
wire Xd_0__inst_mult_5_250 ;
wire Xd_0__inst_mult_4_249 ;
wire Xd_0__inst_mult_4_250 ;
wire Xd_0__inst_mult_7_249 ;
wire Xd_0__inst_mult_7_250 ;
wire Xd_0__inst_mult_6_249 ;
wire Xd_0__inst_mult_6_250 ;
wire Xd_0__inst_mult_1_249 ;
wire Xd_0__inst_mult_1_250 ;
wire Xd_0__inst_mult_0_249 ;
wire Xd_0__inst_mult_0_250 ;
wire Xd_0__inst_mult_3_249 ;
wire Xd_0__inst_mult_3_250 ;
wire Xd_0__inst_mult_2_299 ;
wire Xd_0__inst_mult_2_300 ;
wire Xd_0__inst_mult_29_274 ;
wire Xd_0__inst_mult_29_275 ;
wire Xd_0__inst_mult_28_254 ;
wire Xd_0__inst_mult_28_255 ;
wire Xd_0__inst_mult_31_254 ;
wire Xd_0__inst_mult_31_255 ;
wire Xd_0__inst_mult_30_254 ;
wire Xd_0__inst_mult_30_255 ;
wire Xd_0__inst_mult_25_334 ;
wire Xd_0__inst_mult_25_335 ;
wire Xd_0__inst_mult_24_474 ;
wire Xd_0__inst_mult_24_475 ;
wire Xd_0__inst_mult_27_334 ;
wire Xd_0__inst_mult_27_335 ;
wire Xd_0__inst_mult_26_474 ;
wire Xd_0__inst_mult_26_475 ;
wire Xd_0__inst_mult_21_274 ;
wire Xd_0__inst_mult_21_275 ;
wire Xd_0__inst_mult_20_274 ;
wire Xd_0__inst_mult_20_275 ;
wire Xd_0__inst_mult_23_274 ;
wire Xd_0__inst_mult_23_275 ;
wire Xd_0__inst_mult_22_274 ;
wire Xd_0__inst_mult_22_275 ;
wire Xd_0__inst_mult_17_274 ;
wire Xd_0__inst_mult_17_275 ;
wire Xd_0__inst_mult_16_274 ;
wire Xd_0__inst_mult_16_275 ;
wire Xd_0__inst_mult_19_274 ;
wire Xd_0__inst_mult_19_275 ;
wire Xd_0__inst_mult_18_249 ;
wire Xd_0__inst_mult_18_250 ;
wire Xd_0__inst_mult_13_254 ;
wire Xd_0__inst_mult_13_255 ;
wire Xd_0__inst_mult_12_249 ;
wire Xd_0__inst_mult_12_250 ;
wire Xd_0__inst_mult_15_249 ;
wire Xd_0__inst_mult_15_250 ;
wire Xd_0__inst_mult_14_249 ;
wire Xd_0__inst_mult_14_250 ;
wire Xd_0__inst_mult_9_254 ;
wire Xd_0__inst_mult_9_255 ;
wire Xd_0__inst_mult_8_254 ;
wire Xd_0__inst_mult_8_255 ;
wire Xd_0__inst_mult_11_254 ;
wire Xd_0__inst_mult_11_255 ;
wire Xd_0__inst_mult_10_254 ;
wire Xd_0__inst_mult_10_255 ;
wire Xd_0__inst_mult_5_254 ;
wire Xd_0__inst_mult_5_255 ;
wire Xd_0__inst_mult_4_254 ;
wire Xd_0__inst_mult_4_255 ;
wire Xd_0__inst_mult_7_254 ;
wire Xd_0__inst_mult_7_255 ;
wire Xd_0__inst_mult_6_254 ;
wire Xd_0__inst_mult_6_255 ;
wire Xd_0__inst_mult_1_254 ;
wire Xd_0__inst_mult_1_255 ;
wire Xd_0__inst_mult_0_254 ;
wire Xd_0__inst_mult_0_255 ;
wire Xd_0__inst_mult_3_254 ;
wire Xd_0__inst_mult_3_255 ;
wire Xd_0__inst_mult_2_304 ;
wire Xd_0__inst_mult_2_305 ;
wire Xd_0__inst_mult_29_279 ;
wire Xd_0__inst_mult_29_280 ;
wire Xd_0__inst_mult_28_259 ;
wire Xd_0__inst_mult_28_260 ;
wire Xd_0__inst_mult_31_259 ;
wire Xd_0__inst_mult_31_260 ;
wire Xd_0__inst_mult_30_259 ;
wire Xd_0__inst_mult_30_260 ;
wire Xd_0__inst_mult_25_339 ;
wire Xd_0__inst_mult_25_340 ;
wire Xd_0__inst_mult_24_479 ;
wire Xd_0__inst_mult_24_480 ;
wire Xd_0__inst_mult_27_339 ;
wire Xd_0__inst_mult_27_340 ;
wire Xd_0__inst_mult_26_479 ;
wire Xd_0__inst_mult_26_480 ;
wire Xd_0__inst_mult_21_279 ;
wire Xd_0__inst_mult_21_280 ;
wire Xd_0__inst_mult_20_279 ;
wire Xd_0__inst_mult_20_280 ;
wire Xd_0__inst_mult_23_279 ;
wire Xd_0__inst_mult_23_280 ;
wire Xd_0__inst_mult_22_279 ;
wire Xd_0__inst_mult_22_280 ;
wire Xd_0__inst_mult_17_279 ;
wire Xd_0__inst_mult_17_280 ;
wire Xd_0__inst_mult_16_279 ;
wire Xd_0__inst_mult_16_280 ;
wire Xd_0__inst_mult_19_279 ;
wire Xd_0__inst_mult_19_280 ;
wire Xd_0__inst_mult_18_254 ;
wire Xd_0__inst_mult_18_255 ;
wire Xd_0__inst_mult_13_259 ;
wire Xd_0__inst_mult_13_260 ;
wire Xd_0__inst_mult_12_254 ;
wire Xd_0__inst_mult_12_255 ;
wire Xd_0__inst_mult_15_254 ;
wire Xd_0__inst_mult_15_255 ;
wire Xd_0__inst_mult_14_254 ;
wire Xd_0__inst_mult_14_255 ;
wire Xd_0__inst_mult_9_259 ;
wire Xd_0__inst_mult_9_260 ;
wire Xd_0__inst_mult_8_259 ;
wire Xd_0__inst_mult_8_260 ;
wire Xd_0__inst_mult_11_259 ;
wire Xd_0__inst_mult_11_260 ;
wire Xd_0__inst_mult_10_259 ;
wire Xd_0__inst_mult_10_260 ;
wire Xd_0__inst_mult_5_259 ;
wire Xd_0__inst_mult_5_260 ;
wire Xd_0__inst_mult_4_259 ;
wire Xd_0__inst_mult_4_260 ;
wire Xd_0__inst_mult_7_259 ;
wire Xd_0__inst_mult_7_260 ;
wire Xd_0__inst_mult_6_259 ;
wire Xd_0__inst_mult_6_260 ;
wire Xd_0__inst_mult_1_259 ;
wire Xd_0__inst_mult_1_260 ;
wire Xd_0__inst_mult_0_259 ;
wire Xd_0__inst_mult_0_260 ;
wire Xd_0__inst_mult_3_259 ;
wire Xd_0__inst_mult_3_260 ;
wire Xd_0__inst_mult_2_309 ;
wire Xd_0__inst_mult_2_310 ;
wire Xd_0__inst_mult_29_284 ;
wire Xd_0__inst_mult_29_285 ;
wire Xd_0__inst_mult_28_264 ;
wire Xd_0__inst_mult_28_265 ;
wire Xd_0__inst_mult_31_264 ;
wire Xd_0__inst_mult_31_265 ;
wire Xd_0__inst_mult_30_264 ;
wire Xd_0__inst_mult_30_265 ;
wire Xd_0__inst_mult_25_344 ;
wire Xd_0__inst_mult_25_345 ;
wire Xd_0__inst_mult_24_484 ;
wire Xd_0__inst_mult_24_485 ;
wire Xd_0__inst_mult_27_344 ;
wire Xd_0__inst_mult_27_345 ;
wire Xd_0__inst_mult_26_484 ;
wire Xd_0__inst_mult_26_485 ;
wire Xd_0__inst_mult_21_284 ;
wire Xd_0__inst_mult_21_285 ;
wire Xd_0__inst_mult_20_284 ;
wire Xd_0__inst_mult_20_285 ;
wire Xd_0__inst_mult_23_284 ;
wire Xd_0__inst_mult_23_285 ;
wire Xd_0__inst_mult_22_284 ;
wire Xd_0__inst_mult_22_285 ;
wire Xd_0__inst_mult_17_284 ;
wire Xd_0__inst_mult_17_285 ;
wire Xd_0__inst_mult_16_284 ;
wire Xd_0__inst_mult_16_285 ;
wire Xd_0__inst_mult_19_284 ;
wire Xd_0__inst_mult_19_285 ;
wire Xd_0__inst_mult_18_259 ;
wire Xd_0__inst_mult_18_260 ;
wire Xd_0__inst_mult_13_264 ;
wire Xd_0__inst_mult_13_265 ;
wire Xd_0__inst_mult_12_259 ;
wire Xd_0__inst_mult_12_260 ;
wire Xd_0__inst_mult_15_259 ;
wire Xd_0__inst_mult_15_260 ;
wire Xd_0__inst_mult_14_259 ;
wire Xd_0__inst_mult_14_260 ;
wire Xd_0__inst_mult_9_264 ;
wire Xd_0__inst_mult_9_265 ;
wire Xd_0__inst_mult_8_264 ;
wire Xd_0__inst_mult_8_265 ;
wire Xd_0__inst_mult_11_264 ;
wire Xd_0__inst_mult_11_265 ;
wire Xd_0__inst_mult_10_264 ;
wire Xd_0__inst_mult_10_265 ;
wire Xd_0__inst_mult_5_264 ;
wire Xd_0__inst_mult_5_265 ;
wire Xd_0__inst_mult_4_264 ;
wire Xd_0__inst_mult_4_265 ;
wire Xd_0__inst_mult_7_264 ;
wire Xd_0__inst_mult_7_265 ;
wire Xd_0__inst_mult_6_264 ;
wire Xd_0__inst_mult_6_265 ;
wire Xd_0__inst_mult_1_264 ;
wire Xd_0__inst_mult_1_265 ;
wire Xd_0__inst_mult_0_264 ;
wire Xd_0__inst_mult_0_265 ;
wire Xd_0__inst_mult_3_264 ;
wire Xd_0__inst_mult_3_265 ;
wire Xd_0__inst_mult_2_314 ;
wire Xd_0__inst_mult_2_315 ;
wire Xd_0__inst_mult_29_289 ;
wire Xd_0__inst_mult_29_290 ;
wire Xd_0__inst_mult_28_269 ;
wire Xd_0__inst_mult_28_270 ;
wire Xd_0__inst_mult_31_269 ;
wire Xd_0__inst_mult_31_270 ;
wire Xd_0__inst_mult_30_269 ;
wire Xd_0__inst_mult_30_270 ;
wire Xd_0__inst_mult_25_349 ;
wire Xd_0__inst_mult_25_350 ;
wire Xd_0__inst_mult_24_489 ;
wire Xd_0__inst_mult_24_490 ;
wire Xd_0__inst_mult_27_349 ;
wire Xd_0__inst_mult_27_350 ;
wire Xd_0__inst_mult_26_489 ;
wire Xd_0__inst_mult_26_490 ;
wire Xd_0__inst_mult_21_289 ;
wire Xd_0__inst_mult_21_290 ;
wire Xd_0__inst_mult_20_289 ;
wire Xd_0__inst_mult_20_290 ;
wire Xd_0__inst_mult_23_289 ;
wire Xd_0__inst_mult_23_290 ;
wire Xd_0__inst_mult_22_289 ;
wire Xd_0__inst_mult_22_290 ;
wire Xd_0__inst_mult_17_289 ;
wire Xd_0__inst_mult_17_290 ;
wire Xd_0__inst_mult_16_289 ;
wire Xd_0__inst_mult_16_290 ;
wire Xd_0__inst_mult_19_289 ;
wire Xd_0__inst_mult_19_290 ;
wire Xd_0__inst_mult_18_264 ;
wire Xd_0__inst_mult_18_265 ;
wire Xd_0__inst_mult_13_269 ;
wire Xd_0__inst_mult_13_270 ;
wire Xd_0__inst_mult_12_264 ;
wire Xd_0__inst_mult_12_265 ;
wire Xd_0__inst_mult_15_264 ;
wire Xd_0__inst_mult_15_265 ;
wire Xd_0__inst_mult_14_264 ;
wire Xd_0__inst_mult_14_265 ;
wire Xd_0__inst_mult_9_269 ;
wire Xd_0__inst_mult_9_270 ;
wire Xd_0__inst_mult_8_269 ;
wire Xd_0__inst_mult_8_270 ;
wire Xd_0__inst_mult_11_269 ;
wire Xd_0__inst_mult_11_270 ;
wire Xd_0__inst_mult_10_269 ;
wire Xd_0__inst_mult_10_270 ;
wire Xd_0__inst_mult_5_269 ;
wire Xd_0__inst_mult_5_270 ;
wire Xd_0__inst_mult_4_269 ;
wire Xd_0__inst_mult_4_270 ;
wire Xd_0__inst_mult_7_269 ;
wire Xd_0__inst_mult_7_270 ;
wire Xd_0__inst_mult_6_269 ;
wire Xd_0__inst_mult_6_270 ;
wire Xd_0__inst_mult_1_269 ;
wire Xd_0__inst_mult_1_270 ;
wire Xd_0__inst_mult_0_269 ;
wire Xd_0__inst_mult_0_270 ;
wire Xd_0__inst_mult_3_269 ;
wire Xd_0__inst_mult_3_270 ;
wire Xd_0__inst_mult_2_319 ;
wire Xd_0__inst_mult_2_320 ;
wire Xd_0__inst_mult_29_294 ;
wire Xd_0__inst_mult_29_295 ;
wire Xd_0__inst_mult_28_274 ;
wire Xd_0__inst_mult_28_275 ;
wire Xd_0__inst_mult_31_274 ;
wire Xd_0__inst_mult_31_275 ;
wire Xd_0__inst_mult_30_274 ;
wire Xd_0__inst_mult_30_275 ;
wire Xd_0__inst_mult_25_354 ;
wire Xd_0__inst_mult_25_355 ;
wire Xd_0__inst_mult_24_494 ;
wire Xd_0__inst_mult_24_495 ;
wire Xd_0__inst_mult_27_354 ;
wire Xd_0__inst_mult_27_355 ;
wire Xd_0__inst_mult_26_494 ;
wire Xd_0__inst_mult_26_495 ;
wire Xd_0__inst_mult_21_294 ;
wire Xd_0__inst_mult_21_295 ;
wire Xd_0__inst_mult_20_294 ;
wire Xd_0__inst_mult_20_295 ;
wire Xd_0__inst_mult_23_294 ;
wire Xd_0__inst_mult_23_295 ;
wire Xd_0__inst_mult_22_294 ;
wire Xd_0__inst_mult_22_295 ;
wire Xd_0__inst_mult_17_294 ;
wire Xd_0__inst_mult_17_295 ;
wire Xd_0__inst_mult_16_294 ;
wire Xd_0__inst_mult_16_295 ;
wire Xd_0__inst_mult_19_294 ;
wire Xd_0__inst_mult_19_295 ;
wire Xd_0__inst_mult_18_269 ;
wire Xd_0__inst_mult_18_270 ;
wire Xd_0__inst_mult_13_274 ;
wire Xd_0__inst_mult_13_275 ;
wire Xd_0__inst_mult_12_269 ;
wire Xd_0__inst_mult_12_270 ;
wire Xd_0__inst_mult_15_269 ;
wire Xd_0__inst_mult_15_270 ;
wire Xd_0__inst_mult_14_269 ;
wire Xd_0__inst_mult_14_270 ;
wire Xd_0__inst_mult_9_274 ;
wire Xd_0__inst_mult_9_275 ;
wire Xd_0__inst_mult_8_274 ;
wire Xd_0__inst_mult_8_275 ;
wire Xd_0__inst_mult_11_274 ;
wire Xd_0__inst_mult_11_275 ;
wire Xd_0__inst_mult_10_274 ;
wire Xd_0__inst_mult_10_275 ;
wire Xd_0__inst_mult_5_274 ;
wire Xd_0__inst_mult_5_275 ;
wire Xd_0__inst_mult_4_274 ;
wire Xd_0__inst_mult_4_275 ;
wire Xd_0__inst_mult_7_274 ;
wire Xd_0__inst_mult_7_275 ;
wire Xd_0__inst_mult_6_274 ;
wire Xd_0__inst_mult_6_275 ;
wire Xd_0__inst_mult_1_274 ;
wire Xd_0__inst_mult_1_275 ;
wire Xd_0__inst_mult_0_274 ;
wire Xd_0__inst_mult_0_275 ;
wire Xd_0__inst_mult_3_274 ;
wire Xd_0__inst_mult_3_275 ;
wire Xd_0__inst_mult_2_324 ;
wire Xd_0__inst_mult_2_325 ;
wire Xd_0__inst_mult_29_299 ;
wire Xd_0__inst_mult_29_300 ;
wire Xd_0__inst_mult_28_279 ;
wire Xd_0__inst_mult_28_280 ;
wire Xd_0__inst_mult_31_279 ;
wire Xd_0__inst_mult_31_280 ;
wire Xd_0__inst_mult_30_279 ;
wire Xd_0__inst_mult_30_280 ;
wire Xd_0__inst_mult_25_359 ;
wire Xd_0__inst_mult_25_360 ;
wire Xd_0__inst_mult_24_499 ;
wire Xd_0__inst_mult_24_500 ;
wire Xd_0__inst_mult_27_359 ;
wire Xd_0__inst_mult_27_360 ;
wire Xd_0__inst_mult_26_499 ;
wire Xd_0__inst_mult_26_500 ;
wire Xd_0__inst_mult_21_299 ;
wire Xd_0__inst_mult_21_300 ;
wire Xd_0__inst_mult_20_299 ;
wire Xd_0__inst_mult_20_300 ;
wire Xd_0__inst_mult_23_299 ;
wire Xd_0__inst_mult_23_300 ;
wire Xd_0__inst_mult_22_299 ;
wire Xd_0__inst_mult_22_300 ;
wire Xd_0__inst_mult_17_299 ;
wire Xd_0__inst_mult_17_300 ;
wire Xd_0__inst_mult_16_299 ;
wire Xd_0__inst_mult_16_300 ;
wire Xd_0__inst_mult_19_299 ;
wire Xd_0__inst_mult_19_300 ;
wire Xd_0__inst_mult_18_274 ;
wire Xd_0__inst_mult_18_275 ;
wire Xd_0__inst_mult_13_279 ;
wire Xd_0__inst_mult_13_280 ;
wire Xd_0__inst_mult_12_274 ;
wire Xd_0__inst_mult_12_275 ;
wire Xd_0__inst_mult_15_274 ;
wire Xd_0__inst_mult_15_275 ;
wire Xd_0__inst_mult_14_274 ;
wire Xd_0__inst_mult_14_275 ;
wire Xd_0__inst_mult_9_279 ;
wire Xd_0__inst_mult_9_280 ;
wire Xd_0__inst_mult_8_279 ;
wire Xd_0__inst_mult_8_280 ;
wire Xd_0__inst_mult_11_279 ;
wire Xd_0__inst_mult_11_280 ;
wire Xd_0__inst_mult_10_279 ;
wire Xd_0__inst_mult_10_280 ;
wire Xd_0__inst_mult_5_279 ;
wire Xd_0__inst_mult_5_280 ;
wire Xd_0__inst_mult_4_279 ;
wire Xd_0__inst_mult_4_280 ;
wire Xd_0__inst_mult_7_279 ;
wire Xd_0__inst_mult_7_280 ;
wire Xd_0__inst_mult_6_279 ;
wire Xd_0__inst_mult_6_280 ;
wire Xd_0__inst_mult_1_279 ;
wire Xd_0__inst_mult_1_280 ;
wire Xd_0__inst_mult_0_279 ;
wire Xd_0__inst_mult_0_280 ;
wire Xd_0__inst_mult_3_279 ;
wire Xd_0__inst_mult_3_280 ;
wire Xd_0__inst_mult_2_329 ;
wire Xd_0__inst_mult_2_330 ;
wire Xd_0__inst_mult_29_304 ;
wire Xd_0__inst_mult_29_305 ;
wire Xd_0__inst_mult_28_284 ;
wire Xd_0__inst_mult_28_285 ;
wire Xd_0__inst_mult_31_284 ;
wire Xd_0__inst_mult_31_285 ;
wire Xd_0__inst_mult_30_284 ;
wire Xd_0__inst_mult_30_285 ;
wire Xd_0__inst_mult_25_364 ;
wire Xd_0__inst_mult_25_365 ;
wire Xd_0__inst_mult_24_504 ;
wire Xd_0__inst_mult_24_505 ;
wire Xd_0__inst_mult_27_364 ;
wire Xd_0__inst_mult_27_365 ;
wire Xd_0__inst_mult_26_504 ;
wire Xd_0__inst_mult_26_505 ;
wire Xd_0__inst_mult_21_304 ;
wire Xd_0__inst_mult_21_305 ;
wire Xd_0__inst_mult_20_304 ;
wire Xd_0__inst_mult_20_305 ;
wire Xd_0__inst_mult_23_304 ;
wire Xd_0__inst_mult_23_305 ;
wire Xd_0__inst_mult_22_304 ;
wire Xd_0__inst_mult_22_305 ;
wire Xd_0__inst_mult_17_304 ;
wire Xd_0__inst_mult_17_305 ;
wire Xd_0__inst_mult_16_304 ;
wire Xd_0__inst_mult_16_305 ;
wire Xd_0__inst_mult_19_304 ;
wire Xd_0__inst_mult_19_305 ;
wire Xd_0__inst_mult_18_279 ;
wire Xd_0__inst_mult_18_280 ;
wire Xd_0__inst_mult_13_284 ;
wire Xd_0__inst_mult_13_285 ;
wire Xd_0__inst_mult_12_279 ;
wire Xd_0__inst_mult_12_280 ;
wire Xd_0__inst_mult_15_279 ;
wire Xd_0__inst_mult_15_280 ;
wire Xd_0__inst_mult_14_279 ;
wire Xd_0__inst_mult_14_280 ;
wire Xd_0__inst_mult_9_284 ;
wire Xd_0__inst_mult_9_285 ;
wire Xd_0__inst_mult_8_284 ;
wire Xd_0__inst_mult_8_285 ;
wire Xd_0__inst_mult_11_284 ;
wire Xd_0__inst_mult_11_285 ;
wire Xd_0__inst_mult_10_284 ;
wire Xd_0__inst_mult_10_285 ;
wire Xd_0__inst_mult_5_284 ;
wire Xd_0__inst_mult_5_285 ;
wire Xd_0__inst_mult_4_284 ;
wire Xd_0__inst_mult_4_285 ;
wire Xd_0__inst_mult_7_284 ;
wire Xd_0__inst_mult_7_285 ;
wire Xd_0__inst_mult_6_284 ;
wire Xd_0__inst_mult_6_285 ;
wire Xd_0__inst_mult_1_284 ;
wire Xd_0__inst_mult_1_285 ;
wire Xd_0__inst_mult_0_284 ;
wire Xd_0__inst_mult_0_285 ;
wire Xd_0__inst_mult_3_284 ;
wire Xd_0__inst_mult_3_285 ;
wire Xd_0__inst_mult_2_334 ;
wire Xd_0__inst_mult_2_335 ;
wire Xd_0__inst_mult_29_309 ;
wire Xd_0__inst_mult_28_289 ;
wire Xd_0__inst_mult_31_289 ;
wire Xd_0__inst_mult_30_289 ;
wire Xd_0__inst_mult_25_369 ;
wire Xd_0__inst_mult_24_509 ;
wire Xd_0__inst_mult_27_369 ;
wire Xd_0__inst_mult_26_509 ;
wire Xd_0__inst_mult_21_309 ;
wire Xd_0__inst_mult_20_309 ;
wire Xd_0__inst_mult_23_309 ;
wire Xd_0__inst_mult_22_309 ;
wire Xd_0__inst_mult_17_309 ;
wire Xd_0__inst_mult_16_309 ;
wire Xd_0__inst_mult_19_309 ;
wire Xd_0__inst_mult_18_284 ;
wire Xd_0__inst_mult_13_289 ;
wire Xd_0__inst_mult_12_284 ;
wire Xd_0__inst_mult_15_284 ;
wire Xd_0__inst_mult_14_284 ;
wire Xd_0__inst_mult_9_289 ;
wire Xd_0__inst_mult_8_289 ;
wire Xd_0__inst_mult_11_289 ;
wire Xd_0__inst_mult_10_289 ;
wire Xd_0__inst_mult_5_289 ;
wire Xd_0__inst_mult_4_289 ;
wire Xd_0__inst_mult_7_289 ;
wire Xd_0__inst_mult_6_289 ;
wire Xd_0__inst_mult_1_289 ;
wire Xd_0__inst_mult_0_289 ;
wire Xd_0__inst_mult_3_289 ;
wire Xd_0__inst_mult_2_339 ;
wire Xd_0__inst_i29_41_sumout ;
wire Xd_0__inst_i29_42 ;
wire Xd_0__inst_mult_31_35_sumout ;
wire Xd_0__inst_mult_31_36 ;
wire Xd_0__inst_mult_30_40_sumout ;
wire Xd_0__inst_mult_30_41 ;
wire Xd_0__inst_mult_9_294 ;
wire Xd_0__inst_mult_9_35_sumout ;
wire Xd_0__inst_mult_9_36 ;
wire Xd_0__inst_mult_9_299 ;
wire Xd_0__inst_mult_9_300 ;
wire Xd_0__inst_i29_46_sumout ;
wire Xd_0__inst_i29_47 ;
wire Xd_0__inst_i29_51_sumout ;
wire Xd_0__inst_i29_52 ;
wire Xd_0__inst_mult_29_45_sumout ;
wire Xd_0__inst_mult_29_46 ;
wire Xd_0__inst_mult_28_35_sumout ;
wire Xd_0__inst_mult_28_36 ;
wire Xd_0__inst_mult_8_294 ;
wire Xd_0__inst_mult_8_35_sumout ;
wire Xd_0__inst_mult_8_36 ;
wire Xd_0__inst_mult_8_299 ;
wire Xd_0__inst_mult_8_300 ;
wire Xd_0__inst_mult_21_314 ;
wire Xd_0__inst_mult_21_319 ;
wire Xd_0__inst_mult_21_320 ;
wire Xd_0__inst_mult_21_324 ;
wire Xd_0__inst_mult_21_329 ;
wire Xd_0__inst_mult_21_330 ;
wire Xd_0__inst_i29_56_sumout ;
wire Xd_0__inst_i29_57 ;
wire Xd_0__inst_mult_27_55_sumout ;
wire Xd_0__inst_mult_27_56 ;
wire Xd_0__inst_mult_26_55_sumout ;
wire Xd_0__inst_mult_26_56 ;
wire Xd_0__inst_mult_11_294 ;
wire Xd_0__inst_mult_11_35_sumout ;
wire Xd_0__inst_mult_11_36 ;
wire Xd_0__inst_mult_11_299 ;
wire Xd_0__inst_mult_11_300 ;
wire Xd_0__inst_i29_61_sumout ;
wire Xd_0__inst_i29_62 ;
wire Xd_0__inst_i29_66_sumout ;
wire Xd_0__inst_i29_67 ;
wire Xd_0__inst_mult_25_50_sumout ;
wire Xd_0__inst_mult_25_51 ;
wire Xd_0__inst_mult_24_55_sumout ;
wire Xd_0__inst_mult_24_56 ;
wire Xd_0__inst_mult_10_294 ;
wire Xd_0__inst_mult_10_35_sumout ;
wire Xd_0__inst_mult_10_36 ;
wire Xd_0__inst_mult_10_299 ;
wire Xd_0__inst_mult_10_300 ;
wire Xd_0__inst_mult_20_314 ;
wire Xd_0__inst_mult_20_319 ;
wire Xd_0__inst_mult_20_320 ;
wire Xd_0__inst_mult_14_35_sumout ;
wire Xd_0__inst_mult_14_36 ;
wire Xd_0__inst_mult_20_324 ;
wire Xd_0__inst_mult_20_329 ;
wire Xd_0__inst_mult_20_330 ;
wire Xd_0__inst_mult_25_374 ;
wire Xd_0__inst_mult_25_375 ;
wire Xd_0__inst_mult_25_379 ;
wire Xd_0__inst_mult_25_380 ;
wire Xd_0__inst_mult_25_384 ;
wire Xd_0__inst_mult_25_385 ;
wire Xd_0__inst_mult_25_389 ;
wire Xd_0__inst_mult_25_390 ;
wire Xd_0__inst_i29_71_sumout ;
wire Xd_0__inst_i29_72 ;
wire Xd_0__inst_mult_23_45_sumout ;
wire Xd_0__inst_mult_23_46 ;
wire Xd_0__inst_mult_22_45_sumout ;
wire Xd_0__inst_mult_22_46 ;
wire Xd_0__inst_mult_3_294 ;
wire Xd_0__inst_mult_3_35_sumout ;
wire Xd_0__inst_mult_3_36 ;
wire Xd_0__inst_mult_3_299 ;
wire Xd_0__inst_mult_3_300 ;
wire Xd_0__inst_i29_76_sumout ;
wire Xd_0__inst_i29_77 ;
wire Xd_0__inst_i29_81_sumout ;
wire Xd_0__inst_i29_82 ;
wire Xd_0__inst_mult_21_45_sumout ;
wire Xd_0__inst_mult_21_46 ;
wire Xd_0__inst_mult_20_50_sumout ;
wire Xd_0__inst_mult_20_51 ;
wire Xd_0__inst_mult_0_294 ;
wire Xd_0__inst_mult_0_35_sumout ;
wire Xd_0__inst_mult_0_36 ;
wire Xd_0__inst_mult_0_299 ;
wire Xd_0__inst_mult_0_300 ;
wire Xd_0__inst_mult_23_314 ;
wire Xd_0__inst_mult_23_319 ;
wire Xd_0__inst_mult_23_320 ;
wire Xd_0__inst_mult_23_324 ;
wire Xd_0__inst_mult_23_329 ;
wire Xd_0__inst_mult_23_330 ;
wire Xd_0__inst_i29_86_sumout ;
wire Xd_0__inst_i29_87 ;
wire Xd_0__inst_mult_19_45_sumout ;
wire Xd_0__inst_mult_19_46 ;
wire Xd_0__inst_mult_18_35_sumout ;
wire Xd_0__inst_mult_18_36 ;
wire Xd_0__inst_mult_6_294 ;
wire Xd_0__inst_mult_6_35_sumout ;
wire Xd_0__inst_mult_6_36 ;
wire Xd_0__inst_mult_6_299 ;
wire Xd_0__inst_mult_6_300 ;
wire Xd_0__inst_i29_91_sumout ;
wire Xd_0__inst_i29_92 ;
wire Xd_0__inst_i29_96_sumout ;
wire Xd_0__inst_i29_97 ;
wire Xd_0__inst_mult_17_45_sumout ;
wire Xd_0__inst_mult_17_46 ;
wire Xd_0__inst_mult_16_45_sumout ;
wire Xd_0__inst_mult_16_46 ;
wire Xd_0__inst_mult_1_294 ;
wire Xd_0__inst_mult_1_35_sumout ;
wire Xd_0__inst_mult_1_36 ;
wire Xd_0__inst_mult_1_299 ;
wire Xd_0__inst_mult_1_300 ;
wire Xd_0__inst_mult_22_314 ;
wire Xd_0__inst_mult_22_319 ;
wire Xd_0__inst_mult_22_320 ;
wire Xd_0__inst_mult_22_324 ;
wire Xd_0__inst_mult_22_329 ;
wire Xd_0__inst_mult_22_330 ;
wire Xd_0__inst_mult_24_514 ;
wire Xd_0__inst_mult_24_515 ;
wire Xd_0__inst_mult_24_519 ;
wire Xd_0__inst_mult_24_520 ;
wire Xd_0__inst_mult_24_524 ;
wire Xd_0__inst_mult_24_525 ;
wire Xd_0__inst_mult_24_529 ;
wire Xd_0__inst_mult_24_530 ;
wire Xd_0__inst_mult_26_514 ;
wire Xd_0__inst_mult_26_515 ;
wire Xd_0__inst_mult_26_519 ;
wire Xd_0__inst_mult_26_520 ;
wire Xd_0__inst_mult_26_524 ;
wire Xd_0__inst_mult_26_525 ;
wire Xd_0__inst_mult_26_529 ;
wire Xd_0__inst_mult_26_530 ;
wire Xd_0__inst_mult_26_534 ;
wire Xd_0__inst_mult_26_535 ;
wire Xd_0__inst_i29_101_sumout ;
wire Xd_0__inst_i29_102 ;
wire Xd_0__inst_mult_15_35_sumout ;
wire Xd_0__inst_mult_15_36 ;
wire Xd_0__inst_mult_14_40_sumout ;
wire Xd_0__inst_mult_14_41 ;
wire Xd_0__inst_mult_7_294 ;
wire Xd_0__inst_mult_7_35_sumout ;
wire Xd_0__inst_mult_7_36 ;
wire Xd_0__inst_mult_7_299 ;
wire Xd_0__inst_mult_7_300 ;
wire Xd_0__inst_i29_106_sumout ;
wire Xd_0__inst_i29_107 ;
wire Xd_0__inst_i29_111_sumout ;
wire Xd_0__inst_i29_112 ;
wire Xd_0__inst_mult_13_40_sumout ;
wire Xd_0__inst_mult_13_41 ;
wire Xd_0__inst_mult_12_35_sumout ;
wire Xd_0__inst_mult_12_36 ;
wire Xd_0__inst_mult_4_294 ;
wire Xd_0__inst_mult_4_35_sumout ;
wire Xd_0__inst_mult_4_36 ;
wire Xd_0__inst_mult_4_299 ;
wire Xd_0__inst_mult_4_300 ;
wire Xd_0__inst_mult_19_314 ;
wire Xd_0__inst_mult_19_319 ;
wire Xd_0__inst_mult_19_320 ;
wire Xd_0__inst_mult_19_324 ;
wire Xd_0__inst_mult_19_329 ;
wire Xd_0__inst_mult_19_330 ;
wire Xd_0__inst_i29_116_sumout ;
wire Xd_0__inst_i29_117 ;
wire Xd_0__inst_mult_11_40_sumout ;
wire Xd_0__inst_mult_11_41 ;
wire Xd_0__inst_mult_10_40_sumout ;
wire Xd_0__inst_mult_10_41 ;
wire Xd_0__inst_mult_30_294 ;
wire Xd_0__inst_mult_30_299 ;
wire Xd_0__inst_mult_30_300 ;
wire Xd_0__inst_i29_121_sumout ;
wire Xd_0__inst_i29_122 ;
wire Xd_0__inst_i29_126_sumout ;
wire Xd_0__inst_i29_127 ;
wire Xd_0__inst_mult_9_40_sumout ;
wire Xd_0__inst_mult_9_41 ;
wire Xd_0__inst_mult_8_40_sumout ;
wire Xd_0__inst_mult_8_41 ;
wire Xd_0__inst_mult_5_294 ;
wire Xd_0__inst_mult_5_35_sumout ;
wire Xd_0__inst_mult_5_36 ;
wire Xd_0__inst_mult_5_299 ;
wire Xd_0__inst_mult_5_300 ;
wire Xd_0__inst_mult_17_314 ;
wire Xd_0__inst_mult_17_319 ;
wire Xd_0__inst_mult_17_320 ;
wire Xd_0__inst_mult_17_324 ;
wire Xd_0__inst_mult_17_329 ;
wire Xd_0__inst_mult_17_330 ;
wire Xd_0__inst_mult_27_374 ;
wire Xd_0__inst_mult_27_375 ;
wire Xd_0__inst_mult_27_379 ;
wire Xd_0__inst_mult_27_380 ;
wire Xd_0__inst_mult_27_384 ;
wire Xd_0__inst_mult_27_385 ;
wire Xd_0__inst_mult_27_389 ;
wire Xd_0__inst_mult_27_390 ;
wire Xd_0__inst_i29_131_sumout ;
wire Xd_0__inst_i29_132 ;
wire Xd_0__inst_mult_7_40_sumout ;
wire Xd_0__inst_mult_7_41 ;
wire Xd_0__inst_mult_6_40_sumout ;
wire Xd_0__inst_mult_6_41 ;
wire Xd_0__inst_mult_13_294 ;
wire Xd_0__inst_mult_13_45_sumout ;
wire Xd_0__inst_mult_13_46 ;
wire Xd_0__inst_mult_13_299 ;
wire Xd_0__inst_mult_13_300 ;
wire Xd_0__inst_i29_136_sumout ;
wire Xd_0__inst_i29_137 ;
wire Xd_0__inst_i29_141_sumout ;
wire Xd_0__inst_i29_142 ;
wire Xd_0__inst_mult_5_40_sumout ;
wire Xd_0__inst_mult_5_41 ;
wire Xd_0__inst_mult_4_40_sumout ;
wire Xd_0__inst_mult_4_41 ;
wire Xd_0__inst_mult_2_344 ;
wire Xd_0__inst_mult_2_35_sumout ;
wire Xd_0__inst_mult_2_36 ;
wire Xd_0__inst_mult_2_349 ;
wire Xd_0__inst_mult_2_350 ;
wire Xd_0__inst_mult_16_314 ;
wire Xd_0__inst_mult_16_319 ;
wire Xd_0__inst_mult_16_320 ;
wire Xd_0__inst_mult_16_324 ;
wire Xd_0__inst_mult_16_329 ;
wire Xd_0__inst_mult_16_330 ;
wire Xd_0__inst_i29_146_sumout ;
wire Xd_0__inst_i29_147 ;
wire Xd_0__inst_mult_3_40_sumout ;
wire Xd_0__inst_mult_3_41 ;
wire Xd_0__inst_mult_2_40_sumout ;
wire Xd_0__inst_mult_2_41 ;
wire Xd_0__inst_mult_28_294 ;
wire Xd_0__inst_mult_28_40_sumout ;
wire Xd_0__inst_mult_28_41 ;
wire Xd_0__inst_mult_28_299 ;
wire Xd_0__inst_mult_28_300 ;
wire Xd_0__inst_i29_151_sumout ;
wire Xd_0__inst_i29_152 ;
wire Xd_0__inst_i29_156_sumout ;
wire Xd_0__inst_i29_157 ;
wire Xd_0__inst_mult_1_40_sumout ;
wire Xd_0__inst_mult_1_41 ;
wire Xd_0__inst_mult_0_40_sumout ;
wire Xd_0__inst_mult_0_41 ;
wire Xd_0__inst_mult_31_294 ;
wire Xd_0__inst_mult_31_40_sumout ;
wire Xd_0__inst_mult_31_41 ;
wire Xd_0__inst_mult_31_299 ;
wire Xd_0__inst_mult_31_300 ;
wire Xd_0__inst_mult_29_314 ;
wire Xd_0__inst_mult_29_319 ;
wire Xd_0__inst_mult_29_320 ;
wire Xd_0__inst_mult_29_324 ;
wire Xd_0__inst_mult_29_329 ;
wire Xd_0__inst_mult_29_330 ;
wire Xd_0__inst_mult_26_539 ;
wire Xd_0__inst_mult_26_540 ;
wire Xd_0__inst_mult_26_544 ;
wire Xd_0__inst_mult_26_545 ;
wire Xd_0__inst_mult_26_549 ;
wire Xd_0__inst_mult_26_550 ;
wire Xd_0__inst_mult_26_554 ;
wire Xd_0__inst_mult_26_555 ;
wire Xd_0__inst_mult_24_534 ;
wire Xd_0__inst_mult_24_535 ;
wire Xd_0__inst_mult_24_539 ;
wire Xd_0__inst_mult_24_540 ;
wire Xd_0__inst_mult_24_544 ;
wire Xd_0__inst_mult_24_545 ;
wire Xd_0__inst_mult_24_549 ;
wire Xd_0__inst_mult_24_550 ;
wire Xd_0__inst_mult_24_554 ;
wire Xd_0__inst_mult_24_555 ;
wire Xd_0__inst_mult_2_354 ;
wire Xd_0__inst_mult_2_355 ;
wire Xd_0__inst_mult_29_334 ;
wire Xd_0__inst_mult_29_335 ;
wire Xd_0__inst_mult_28_304 ;
wire Xd_0__inst_mult_28_305 ;
wire Xd_0__inst_mult_31_304 ;
wire Xd_0__inst_mult_31_305 ;
wire Xd_0__inst_mult_30_304 ;
wire Xd_0__inst_mult_30_305 ;
wire Xd_0__inst_mult_25_394 ;
wire Xd_0__inst_mult_25_395 ;
wire Xd_0__inst_mult_24_559 ;
wire Xd_0__inst_mult_24_560 ;
wire Xd_0__inst_mult_27_394 ;
wire Xd_0__inst_mult_27_395 ;
wire Xd_0__inst_mult_26_559 ;
wire Xd_0__inst_mult_26_560 ;
wire Xd_0__inst_mult_21_334 ;
wire Xd_0__inst_mult_21_335 ;
wire Xd_0__inst_mult_20_334 ;
wire Xd_0__inst_mult_20_335 ;
wire Xd_0__inst_mult_23_334 ;
wire Xd_0__inst_mult_23_335 ;
wire Xd_0__inst_mult_22_334 ;
wire Xd_0__inst_mult_22_335 ;
wire Xd_0__inst_mult_17_334 ;
wire Xd_0__inst_mult_17_335 ;
wire Xd_0__inst_mult_16_334 ;
wire Xd_0__inst_mult_16_335 ;
wire Xd_0__inst_mult_19_334 ;
wire Xd_0__inst_mult_19_335 ;
wire Xd_0__inst_mult_18_289 ;
wire Xd_0__inst_mult_18_290 ;
wire Xd_0__inst_mult_13_304 ;
wire Xd_0__inst_mult_13_305 ;
wire Xd_0__inst_mult_12_289 ;
wire Xd_0__inst_mult_12_290 ;
wire Xd_0__inst_mult_15_289 ;
wire Xd_0__inst_mult_15_290 ;
wire Xd_0__inst_mult_14_289 ;
wire Xd_0__inst_mult_14_290 ;
wire Xd_0__inst_mult_9_304 ;
wire Xd_0__inst_mult_9_305 ;
wire Xd_0__inst_mult_8_304 ;
wire Xd_0__inst_mult_8_305 ;
wire Xd_0__inst_mult_11_304 ;
wire Xd_0__inst_mult_11_305 ;
wire Xd_0__inst_mult_10_304 ;
wire Xd_0__inst_mult_10_305 ;
wire Xd_0__inst_mult_5_304 ;
wire Xd_0__inst_mult_5_305 ;
wire Xd_0__inst_mult_4_304 ;
wire Xd_0__inst_mult_4_305 ;
wire Xd_0__inst_mult_7_304 ;
wire Xd_0__inst_mult_7_305 ;
wire Xd_0__inst_mult_6_304 ;
wire Xd_0__inst_mult_6_305 ;
wire Xd_0__inst_mult_1_304 ;
wire Xd_0__inst_mult_1_305 ;
wire Xd_0__inst_mult_0_304 ;
wire Xd_0__inst_mult_0_305 ;
wire Xd_0__inst_mult_3_304 ;
wire Xd_0__inst_mult_3_305 ;
wire Xd_0__inst_mult_2_359 ;
wire Xd_0__inst_mult_2_360 ;
wire Xd_0__inst_mult_29_339 ;
wire Xd_0__inst_mult_29_340 ;
wire Xd_0__inst_mult_28_309 ;
wire Xd_0__inst_mult_28_310 ;
wire Xd_0__inst_mult_31_309 ;
wire Xd_0__inst_mult_31_310 ;
wire Xd_0__inst_mult_30_309 ;
wire Xd_0__inst_mult_30_310 ;
wire Xd_0__inst_mult_25_399 ;
wire Xd_0__inst_mult_25_400 ;
wire Xd_0__inst_mult_24_564 ;
wire Xd_0__inst_mult_24_565 ;
wire Xd_0__inst_mult_27_399 ;
wire Xd_0__inst_mult_27_400 ;
wire Xd_0__inst_mult_26_564 ;
wire Xd_0__inst_mult_26_565 ;
wire Xd_0__inst_mult_21_339 ;
wire Xd_0__inst_mult_21_340 ;
wire Xd_0__inst_mult_20_339 ;
wire Xd_0__inst_mult_20_340 ;
wire Xd_0__inst_mult_23_339 ;
wire Xd_0__inst_mult_23_340 ;
wire Xd_0__inst_mult_22_339 ;
wire Xd_0__inst_mult_22_340 ;
wire Xd_0__inst_mult_17_339 ;
wire Xd_0__inst_mult_17_340 ;
wire Xd_0__inst_mult_16_339 ;
wire Xd_0__inst_mult_16_340 ;
wire Xd_0__inst_mult_19_339 ;
wire Xd_0__inst_mult_19_340 ;
wire Xd_0__inst_mult_18_294 ;
wire Xd_0__inst_mult_18_295 ;
wire Xd_0__inst_mult_13_309 ;
wire Xd_0__inst_mult_13_310 ;
wire Xd_0__inst_mult_12_294 ;
wire Xd_0__inst_mult_12_295 ;
wire Xd_0__inst_mult_15_294 ;
wire Xd_0__inst_mult_15_295 ;
wire Xd_0__inst_mult_14_294 ;
wire Xd_0__inst_mult_14_295 ;
wire Xd_0__inst_mult_9_309 ;
wire Xd_0__inst_mult_9_310 ;
wire Xd_0__inst_mult_8_309 ;
wire Xd_0__inst_mult_8_310 ;
wire Xd_0__inst_mult_11_309 ;
wire Xd_0__inst_mult_11_310 ;
wire Xd_0__inst_mult_10_309 ;
wire Xd_0__inst_mult_10_310 ;
wire Xd_0__inst_mult_5_309 ;
wire Xd_0__inst_mult_5_310 ;
wire Xd_0__inst_mult_4_309 ;
wire Xd_0__inst_mult_4_310 ;
wire Xd_0__inst_mult_7_309 ;
wire Xd_0__inst_mult_7_310 ;
wire Xd_0__inst_mult_6_309 ;
wire Xd_0__inst_mult_6_310 ;
wire Xd_0__inst_mult_1_309 ;
wire Xd_0__inst_mult_1_310 ;
wire Xd_0__inst_mult_0_309 ;
wire Xd_0__inst_mult_0_310 ;
wire Xd_0__inst_mult_3_309 ;
wire Xd_0__inst_mult_3_310 ;
wire Xd_0__inst_mult_2_364 ;
wire Xd_0__inst_mult_2_365 ;
wire Xd_0__inst_mult_29_344 ;
wire Xd_0__inst_mult_29_345 ;
wire Xd_0__inst_mult_28_314 ;
wire Xd_0__inst_mult_28_315 ;
wire Xd_0__inst_mult_31_314 ;
wire Xd_0__inst_mult_31_315 ;
wire Xd_0__inst_mult_30_314 ;
wire Xd_0__inst_mult_30_315 ;
wire Xd_0__inst_mult_25_404 ;
wire Xd_0__inst_mult_25_405 ;
wire Xd_0__inst_mult_24_569 ;
wire Xd_0__inst_mult_24_570 ;
wire Xd_0__inst_mult_27_404 ;
wire Xd_0__inst_mult_27_405 ;
wire Xd_0__inst_mult_26_569 ;
wire Xd_0__inst_mult_26_570 ;
wire Xd_0__inst_mult_21_344 ;
wire Xd_0__inst_mult_21_345 ;
wire Xd_0__inst_mult_20_344 ;
wire Xd_0__inst_mult_20_345 ;
wire Xd_0__inst_mult_23_344 ;
wire Xd_0__inst_mult_23_345 ;
wire Xd_0__inst_mult_22_344 ;
wire Xd_0__inst_mult_22_345 ;
wire Xd_0__inst_mult_17_344 ;
wire Xd_0__inst_mult_17_345 ;
wire Xd_0__inst_mult_16_344 ;
wire Xd_0__inst_mult_16_345 ;
wire Xd_0__inst_mult_19_344 ;
wire Xd_0__inst_mult_19_345 ;
wire Xd_0__inst_mult_18_299 ;
wire Xd_0__inst_mult_18_300 ;
wire Xd_0__inst_mult_13_314 ;
wire Xd_0__inst_mult_13_315 ;
wire Xd_0__inst_mult_12_299 ;
wire Xd_0__inst_mult_12_300 ;
wire Xd_0__inst_mult_15_299 ;
wire Xd_0__inst_mult_15_300 ;
wire Xd_0__inst_mult_14_299 ;
wire Xd_0__inst_mult_14_300 ;
wire Xd_0__inst_mult_9_314 ;
wire Xd_0__inst_mult_9_315 ;
wire Xd_0__inst_mult_8_314 ;
wire Xd_0__inst_mult_8_315 ;
wire Xd_0__inst_mult_11_314 ;
wire Xd_0__inst_mult_11_315 ;
wire Xd_0__inst_mult_10_314 ;
wire Xd_0__inst_mult_10_315 ;
wire Xd_0__inst_mult_5_314 ;
wire Xd_0__inst_mult_5_315 ;
wire Xd_0__inst_mult_4_314 ;
wire Xd_0__inst_mult_4_315 ;
wire Xd_0__inst_mult_7_314 ;
wire Xd_0__inst_mult_7_315 ;
wire Xd_0__inst_mult_6_314 ;
wire Xd_0__inst_mult_6_315 ;
wire Xd_0__inst_mult_1_314 ;
wire Xd_0__inst_mult_1_315 ;
wire Xd_0__inst_mult_0_314 ;
wire Xd_0__inst_mult_0_315 ;
wire Xd_0__inst_mult_3_314 ;
wire Xd_0__inst_mult_3_315 ;
wire Xd_0__inst_mult_2_369 ;
wire Xd_0__inst_mult_2_370 ;
wire Xd_0__inst_mult_29_349 ;
wire Xd_0__inst_mult_29_350 ;
wire Xd_0__inst_mult_28_319 ;
wire Xd_0__inst_mult_28_320 ;
wire Xd_0__inst_mult_31_319 ;
wire Xd_0__inst_mult_31_320 ;
wire Xd_0__inst_mult_30_319 ;
wire Xd_0__inst_mult_30_320 ;
wire Xd_0__inst_mult_25_409 ;
wire Xd_0__inst_mult_25_410 ;
wire Xd_0__inst_mult_24_574 ;
wire Xd_0__inst_mult_24_575 ;
wire Xd_0__inst_mult_27_409 ;
wire Xd_0__inst_mult_27_410 ;
wire Xd_0__inst_mult_26_574 ;
wire Xd_0__inst_mult_26_575 ;
wire Xd_0__inst_mult_21_349 ;
wire Xd_0__inst_mult_21_350 ;
wire Xd_0__inst_mult_20_349 ;
wire Xd_0__inst_mult_20_350 ;
wire Xd_0__inst_mult_23_349 ;
wire Xd_0__inst_mult_23_350 ;
wire Xd_0__inst_mult_22_349 ;
wire Xd_0__inst_mult_22_350 ;
wire Xd_0__inst_mult_17_349 ;
wire Xd_0__inst_mult_17_350 ;
wire Xd_0__inst_mult_16_349 ;
wire Xd_0__inst_mult_16_350 ;
wire Xd_0__inst_mult_19_349 ;
wire Xd_0__inst_mult_19_350 ;
wire Xd_0__inst_mult_18_304 ;
wire Xd_0__inst_mult_18_305 ;
wire Xd_0__inst_mult_13_319 ;
wire Xd_0__inst_mult_13_320 ;
wire Xd_0__inst_mult_12_304 ;
wire Xd_0__inst_mult_12_305 ;
wire Xd_0__inst_mult_15_304 ;
wire Xd_0__inst_mult_15_305 ;
wire Xd_0__inst_mult_14_304 ;
wire Xd_0__inst_mult_14_305 ;
wire Xd_0__inst_mult_9_319 ;
wire Xd_0__inst_mult_9_320 ;
wire Xd_0__inst_mult_8_319 ;
wire Xd_0__inst_mult_8_320 ;
wire Xd_0__inst_mult_11_319 ;
wire Xd_0__inst_mult_11_320 ;
wire Xd_0__inst_mult_10_319 ;
wire Xd_0__inst_mult_10_320 ;
wire Xd_0__inst_mult_5_319 ;
wire Xd_0__inst_mult_5_320 ;
wire Xd_0__inst_mult_4_319 ;
wire Xd_0__inst_mult_4_320 ;
wire Xd_0__inst_mult_7_319 ;
wire Xd_0__inst_mult_7_320 ;
wire Xd_0__inst_mult_6_319 ;
wire Xd_0__inst_mult_6_320 ;
wire Xd_0__inst_mult_1_319 ;
wire Xd_0__inst_mult_1_320 ;
wire Xd_0__inst_mult_0_319 ;
wire Xd_0__inst_mult_0_320 ;
wire Xd_0__inst_mult_3_319 ;
wire Xd_0__inst_mult_3_320 ;
wire Xd_0__inst_mult_2_374 ;
wire Xd_0__inst_mult_2_375 ;
wire Xd_0__inst_mult_18_40_sumout ;
wire Xd_0__inst_mult_18_41 ;
wire Xd_0__inst_mult_17_50_sumout ;
wire Xd_0__inst_mult_17_51 ;
wire Xd_0__inst_mult_20_55_sumout ;
wire Xd_0__inst_mult_20_56 ;
wire Xd_0__inst_mult_2_45_sumout ;
wire Xd_0__inst_mult_2_46 ;
wire Xd_0__inst_mult_25_55_sumout ;
wire Xd_0__inst_mult_25_56 ;
wire Xd_0__inst_mult_28_45_sumout ;
wire Xd_0__inst_mult_28_46 ;
wire Xd_0__inst_mult_3_45_sumout ;
wire Xd_0__inst_mult_3_46 ;
wire Xd_0__inst_mult_6_45_sumout ;
wire Xd_0__inst_mult_6_46 ;
wire Xd_0__inst_mult_8_45_sumout ;
wire Xd_0__inst_mult_8_46 ;
wire Xd_0__inst_mult_8_50_sumout ;
wire Xd_0__inst_mult_8_51 ;
wire Xd_0__inst_mult_15_40_sumout ;
wire Xd_0__inst_mult_15_41 ;
wire Xd_0__inst_mult_5_45_sumout ;
wire Xd_0__inst_mult_5_46 ;
wire Xd_0__inst_mult_2_50_sumout ;
wire Xd_0__inst_mult_2_51 ;
wire Xd_0__inst_mult_14_45_sumout ;
wire Xd_0__inst_mult_14_46 ;
wire Xd_0__inst_mult_11_45_sumout ;
wire Xd_0__inst_mult_11_46 ;
wire Xd_0__inst_mult_4_45_sumout ;
wire Xd_0__inst_mult_4_46 ;
wire Xd_0__inst_mult_1_45_sumout ;
wire Xd_0__inst_mult_1_46 ;
wire Xd_0__inst_mult_2_55_sumout ;
wire Xd_0__inst_mult_2_56 ;
wire Xd_0__inst_mult_0_45_sumout ;
wire Xd_0__inst_mult_0_46 ;
wire Xd_0__inst_mult_31_45_sumout ;
wire Xd_0__inst_mult_31_46 ;
wire Xd_0__inst_mult_25_60_sumout ;
wire Xd_0__inst_mult_25_61 ;
wire Xd_0__inst_mult_28_50_sumout ;
wire Xd_0__inst_mult_28_51 ;
wire Xd_0__inst_mult_3_50_sumout ;
wire Xd_0__inst_mult_3_51 ;
wire Xd_0__inst_mult_27_60_sumout ;
wire Xd_0__inst_mult_27_61 ;
wire Xd_0__inst_mult_5_50_sumout ;
wire Xd_0__inst_mult_5_51 ;
wire Xd_0__inst_mult_8_55_sumout ;
wire Xd_0__inst_mult_8_56 ;
wire Xd_0__inst_mult_15_45_sumout ;
wire Xd_0__inst_mult_15_46 ;
wire Xd_0__inst_mult_6_50_sumout ;
wire Xd_0__inst_mult_6_51 ;
wire Xd_0__inst_mult_5_55_sumout ;
wire Xd_0__inst_mult_5_56 ;
wire Xd_0__inst_mult_18_45_sumout ;
wire Xd_0__inst_mult_18_46 ;
wire Xd_0__inst_mult_9_324 ;
wire Xd_0__inst_mult_9_325 ;
wire Xd_0__inst_mult_9_45_sumout ;
wire Xd_0__inst_mult_9_46 ;
wire Xd_0__inst_mult_9_329 ;
wire Xd_0__inst_mult_9_330 ;
wire Xd_0__inst_mult_5_60_sumout ;
wire Xd_0__inst_mult_5_61 ;
wire Xd_0__inst_mult_8_324 ;
wire Xd_0__inst_mult_8_325 ;
wire Xd_0__inst_mult_8_60_sumout ;
wire Xd_0__inst_mult_8_61 ;
wire Xd_0__inst_mult_8_329 ;
wire Xd_0__inst_mult_8_330 ;
wire Xd_0__inst_mult_21_354 ;
wire Xd_0__inst_mult_21_355 ;
wire Xd_0__inst_mult_21_359 ;
wire Xd_0__inst_mult_21_360 ;
wire Xd_0__inst_mult_21_364 ;
wire Xd_0__inst_mult_21_365 ;
wire Xd_0__inst_mult_21_369 ;
wire Xd_0__inst_mult_21_370 ;
wire Xd_0__inst_mult_11_324 ;
wire Xd_0__inst_mult_11_325 ;
wire Xd_0__inst_mult_11_329 ;
wire Xd_0__inst_mult_11_330 ;
wire Xd_0__inst_mult_10_324 ;
wire Xd_0__inst_mult_10_325 ;
wire Xd_0__inst_mult_10_45_sumout ;
wire Xd_0__inst_mult_10_46 ;
wire Xd_0__inst_mult_10_329 ;
wire Xd_0__inst_mult_10_330 ;
wire Xd_0__inst_mult_20_354 ;
wire Xd_0__inst_mult_20_355 ;
wire Xd_0__inst_mult_20_359 ;
wire Xd_0__inst_mult_20_360 ;
wire Xd_0__inst_mult_15_50_sumout ;
wire Xd_0__inst_mult_15_51 ;
wire Xd_0__inst_mult_20_364 ;
wire Xd_0__inst_mult_20_365 ;
wire Xd_0__inst_mult_20_369 ;
wire Xd_0__inst_mult_20_370 ;
wire Xd_0__inst_mult_25_414 ;
wire Xd_0__inst_mult_25_415 ;
wire Xd_0__inst_mult_25_419 ;
wire Xd_0__inst_mult_25_420 ;
wire Xd_0__inst_mult_25_424 ;
wire Xd_0__inst_mult_25_425 ;
wire Xd_0__inst_mult_25_429 ;
wire Xd_0__inst_mult_25_430 ;
wire Xd_0__inst_mult_3_324 ;
wire Xd_0__inst_mult_3_325 ;
wire Xd_0__inst_mult_15_55_sumout ;
wire Xd_0__inst_mult_15_56 ;
wire Xd_0__inst_mult_3_55_sumout ;
wire Xd_0__inst_mult_3_56 ;
wire Xd_0__inst_mult_3_329 ;
wire Xd_0__inst_mult_3_330 ;
wire Xd_0__inst_mult_0_324 ;
wire Xd_0__inst_mult_0_325 ;
wire Xd_0__inst_mult_0_329 ;
wire Xd_0__inst_mult_0_330 ;
wire Xd_0__inst_mult_23_354 ;
wire Xd_0__inst_mult_23_355 ;
wire Xd_0__inst_mult_23_359 ;
wire Xd_0__inst_mult_23_360 ;
wire Xd_0__inst_mult_23_364 ;
wire Xd_0__inst_mult_23_365 ;
wire Xd_0__inst_mult_23_369 ;
wire Xd_0__inst_mult_23_370 ;
wire Xd_0__inst_mult_17_55_sumout ;
wire Xd_0__inst_mult_17_56 ;
wire Xd_0__inst_mult_16_50_sumout ;
wire Xd_0__inst_mult_16_51 ;
wire Xd_0__inst_mult_6_324 ;
wire Xd_0__inst_mult_6_325 ;
wire Xd_0__inst_mult_6_55_sumout ;
wire Xd_0__inst_mult_6_56 ;
wire Xd_0__inst_mult_6_329 ;
wire Xd_0__inst_mult_6_330 ;
wire Xd_0__inst_mult_1_324 ;
wire Xd_0__inst_mult_1_325 ;
wire Xd_0__inst_mult_1_329 ;
wire Xd_0__inst_mult_1_330 ;
wire Xd_0__inst_mult_22_354 ;
wire Xd_0__inst_mult_22_355 ;
wire Xd_0__inst_mult_22_359 ;
wire Xd_0__inst_mult_22_360 ;
wire Xd_0__inst_mult_22_364 ;
wire Xd_0__inst_mult_22_365 ;
wire Xd_0__inst_mult_22_369 ;
wire Xd_0__inst_mult_22_370 ;
wire Xd_0__inst_mult_24_579 ;
wire Xd_0__inst_mult_24_580 ;
wire Xd_0__inst_mult_24_584 ;
wire Xd_0__inst_mult_24_585 ;
wire Xd_0__inst_mult_24_589 ;
wire Xd_0__inst_mult_24_590 ;
wire Xd_0__inst_mult_24_594 ;
wire Xd_0__inst_mult_24_595 ;
wire Xd_0__inst_mult_26_579 ;
wire Xd_0__inst_mult_26_580 ;
wire Xd_0__inst_mult_26_584 ;
wire Xd_0__inst_mult_26_585 ;
wire Xd_0__inst_mult_26_589 ;
wire Xd_0__inst_mult_26_590 ;
wire Xd_0__inst_mult_26_594 ;
wire Xd_0__inst_mult_26_595 ;
wire Xd_0__inst_mult_26_599 ;
wire Xd_0__inst_mult_26_600 ;
wire Xd_0__inst_mult_7_324 ;
wire Xd_0__inst_mult_7_325 ;
wire Xd_0__inst_mult_7_45_sumout ;
wire Xd_0__inst_mult_7_46 ;
wire Xd_0__inst_mult_7_329 ;
wire Xd_0__inst_mult_7_330 ;
wire Xd_0__inst_mult_4_324 ;
wire Xd_0__inst_mult_4_325 ;
wire Xd_0__inst_mult_4_329 ;
wire Xd_0__inst_mult_4_330 ;
wire Xd_0__inst_mult_19_354 ;
wire Xd_0__inst_mult_19_355 ;
wire Xd_0__inst_mult_19_359 ;
wire Xd_0__inst_mult_19_360 ;
wire Xd_0__inst_mult_19_364 ;
wire Xd_0__inst_mult_19_365 ;
wire Xd_0__inst_mult_19_369 ;
wire Xd_0__inst_mult_19_370 ;
wire Xd_0__inst_mult_30_324 ;
wire Xd_0__inst_mult_30_325 ;
wire Xd_0__inst_mult_30_45_sumout ;
wire Xd_0__inst_mult_30_46 ;
wire Xd_0__inst_mult_30_329 ;
wire Xd_0__inst_mult_30_330 ;
wire Xd_0__inst_mult_28_55_sumout ;
wire Xd_0__inst_mult_28_56 ;
wire Xd_0__inst_mult_5_324 ;
wire Xd_0__inst_mult_5_325 ;
wire Xd_0__inst_mult_5_65_sumout ;
wire Xd_0__inst_mult_5_66 ;
wire Xd_0__inst_mult_5_329 ;
wire Xd_0__inst_mult_5_330 ;
wire Xd_0__inst_mult_17_354 ;
wire Xd_0__inst_mult_17_355 ;
wire Xd_0__inst_mult_17_359 ;
wire Xd_0__inst_mult_17_360 ;
wire Xd_0__inst_mult_17_364 ;
wire Xd_0__inst_mult_17_365 ;
wire Xd_0__inst_mult_17_369 ;
wire Xd_0__inst_mult_17_370 ;
wire Xd_0__inst_mult_27_414 ;
wire Xd_0__inst_mult_27_415 ;
wire Xd_0__inst_mult_27_419 ;
wire Xd_0__inst_mult_27_420 ;
wire Xd_0__inst_mult_27_424 ;
wire Xd_0__inst_mult_27_425 ;
wire Xd_0__inst_mult_27_429 ;
wire Xd_0__inst_mult_27_430 ;
wire Xd_0__inst_mult_31_50_sumout ;
wire Xd_0__inst_mult_31_51 ;
wire Xd_0__inst_mult_13_324 ;
wire Xd_0__inst_mult_13_325 ;
wire Xd_0__inst_mult_18_50_sumout ;
wire Xd_0__inst_mult_18_51 ;
wire Xd_0__inst_mult_13_50_sumout ;
wire Xd_0__inst_mult_13_51 ;
wire Xd_0__inst_mult_13_329 ;
wire Xd_0__inst_mult_13_330 ;
wire Xd_0__inst_mult_2_379 ;
wire Xd_0__inst_mult_2_380 ;
wire Xd_0__inst_mult_2_384 ;
wire Xd_0__inst_mult_2_385 ;
wire Xd_0__inst_mult_16_354 ;
wire Xd_0__inst_mult_16_355 ;
wire Xd_0__inst_mult_16_359 ;
wire Xd_0__inst_mult_16_360 ;
wire Xd_0__inst_mult_16_364 ;
wire Xd_0__inst_mult_16_365 ;
wire Xd_0__inst_mult_16_369 ;
wire Xd_0__inst_mult_16_370 ;
wire Xd_0__inst_mult_28_324 ;
wire Xd_0__inst_mult_28_325 ;
wire Xd_0__inst_mult_28_60_sumout ;
wire Xd_0__inst_mult_28_61 ;
wire Xd_0__inst_mult_28_329 ;
wire Xd_0__inst_mult_28_330 ;
wire Xd_0__inst_mult_5_70_sumout ;
wire Xd_0__inst_mult_5_71 ;
wire Xd_0__inst_mult_31_324 ;
wire Xd_0__inst_mult_31_325 ;
wire Xd_0__inst_mult_31_329 ;
wire Xd_0__inst_mult_31_330 ;
wire Xd_0__inst_mult_29_354 ;
wire Xd_0__inst_mult_29_355 ;
wire Xd_0__inst_mult_29_359 ;
wire Xd_0__inst_mult_29_360 ;
wire Xd_0__inst_mult_29_364 ;
wire Xd_0__inst_mult_29_365 ;
wire Xd_0__inst_mult_29_369 ;
wire Xd_0__inst_mult_29_370 ;
wire Xd_0__inst_mult_26_604 ;
wire Xd_0__inst_mult_26_605 ;
wire Xd_0__inst_mult_26_609 ;
wire Xd_0__inst_mult_26_610 ;
wire Xd_0__inst_mult_26_614 ;
wire Xd_0__inst_mult_26_615 ;
wire Xd_0__inst_mult_26_619 ;
wire Xd_0__inst_mult_26_620 ;
wire Xd_0__inst_mult_24_599 ;
wire Xd_0__inst_mult_24_600 ;
wire Xd_0__inst_mult_24_604 ;
wire Xd_0__inst_mult_24_605 ;
wire Xd_0__inst_mult_24_609 ;
wire Xd_0__inst_mult_24_610 ;
wire Xd_0__inst_mult_24_614 ;
wire Xd_0__inst_mult_24_615 ;
wire Xd_0__inst_mult_24_619 ;
wire Xd_0__inst_mult_24_620 ;
wire Xd_0__inst_mult_2_389 ;
wire Xd_0__inst_mult_2_390 ;
wire Xd_0__inst_mult_29_374 ;
wire Xd_0__inst_mult_29_375 ;
wire Xd_0__inst_mult_29_379 ;
wire Xd_0__inst_mult_29_380 ;
wire Xd_0__inst_mult_28_334 ;
wire Xd_0__inst_mult_28_335 ;
wire Xd_0__inst_mult_28_339 ;
wire Xd_0__inst_mult_28_340 ;
wire Xd_0__inst_mult_31_334 ;
wire Xd_0__inst_mult_31_335 ;
wire Xd_0__inst_mult_31_339 ;
wire Xd_0__inst_mult_31_340 ;
wire Xd_0__inst_mult_12_40_sumout ;
wire Xd_0__inst_mult_12_41 ;
wire Xd_0__inst_mult_30_334 ;
wire Xd_0__inst_mult_30_335 ;
wire Xd_0__inst_mult_30_339 ;
wire Xd_0__inst_mult_30_340 ;
wire Xd_0__inst_mult_25_434 ;
wire Xd_0__inst_mult_25_435 ;
wire Xd_0__inst_mult_25_439 ;
wire Xd_0__inst_mult_25_440 ;
wire Xd_0__inst_mult_24_624 ;
wire Xd_0__inst_mult_24_625 ;
wire Xd_0__inst_mult_24_629 ;
wire Xd_0__inst_mult_24_630 ;
wire Xd_0__inst_mult_27_434 ;
wire Xd_0__inst_mult_27_435 ;
wire Xd_0__inst_mult_27_439 ;
wire Xd_0__inst_mult_27_440 ;
wire Xd_0__inst_mult_26_624 ;
wire Xd_0__inst_mult_26_625 ;
wire Xd_0__inst_mult_26_629 ;
wire Xd_0__inst_mult_26_630 ;
wire Xd_0__inst_mult_21_374 ;
wire Xd_0__inst_mult_21_375 ;
wire Xd_0__inst_mult_21_379 ;
wire Xd_0__inst_mult_21_380 ;
wire Xd_0__inst_mult_20_374 ;
wire Xd_0__inst_mult_20_375 ;
wire Xd_0__inst_mult_20_379 ;
wire Xd_0__inst_mult_20_380 ;
wire Xd_0__inst_mult_23_374 ;
wire Xd_0__inst_mult_23_375 ;
wire Xd_0__inst_mult_23_379 ;
wire Xd_0__inst_mult_23_380 ;
wire Xd_0__inst_mult_22_374 ;
wire Xd_0__inst_mult_22_375 ;
wire Xd_0__inst_mult_22_379 ;
wire Xd_0__inst_mult_22_380 ;
wire Xd_0__inst_mult_17_374 ;
wire Xd_0__inst_mult_17_375 ;
wire Xd_0__inst_mult_17_379 ;
wire Xd_0__inst_mult_17_380 ;
wire Xd_0__inst_mult_16_374 ;
wire Xd_0__inst_mult_16_375 ;
wire Xd_0__inst_mult_16_379 ;
wire Xd_0__inst_mult_16_380 ;
wire Xd_0__inst_mult_19_374 ;
wire Xd_0__inst_mult_19_375 ;
wire Xd_0__inst_mult_19_379 ;
wire Xd_0__inst_mult_19_380 ;
wire Xd_0__inst_mult_18_309 ;
wire Xd_0__inst_mult_18_310 ;
wire Xd_0__inst_mult_18_314 ;
wire Xd_0__inst_mult_18_315 ;
wire Xd_0__inst_mult_17_60_sumout ;
wire Xd_0__inst_mult_17_61 ;
wire Xd_0__inst_mult_13_334 ;
wire Xd_0__inst_mult_13_335 ;
wire Xd_0__inst_mult_13_339 ;
wire Xd_0__inst_mult_13_340 ;
wire Xd_0__inst_mult_12_309 ;
wire Xd_0__inst_mult_12_310 ;
wire Xd_0__inst_mult_12_314 ;
wire Xd_0__inst_mult_12_315 ;
wire Xd_0__inst_mult_15_60_sumout ;
wire Xd_0__inst_mult_15_61 ;
wire Xd_0__inst_mult_15_309 ;
wire Xd_0__inst_mult_15_310 ;
wire Xd_0__inst_mult_15_314 ;
wire Xd_0__inst_mult_15_315 ;
wire Xd_0__inst_mult_5_75_sumout ;
wire Xd_0__inst_mult_5_76 ;
wire Xd_0__inst_mult_14_309 ;
wire Xd_0__inst_mult_14_310 ;
wire Xd_0__inst_mult_14_314 ;
wire Xd_0__inst_mult_14_315 ;
wire Xd_0__inst_mult_3_60_sumout ;
wire Xd_0__inst_mult_3_61 ;
wire Xd_0__inst_mult_9_334 ;
wire Xd_0__inst_mult_9_335 ;
wire Xd_0__inst_mult_9_339 ;
wire Xd_0__inst_mult_9_340 ;
wire Xd_0__inst_mult_8_334 ;
wire Xd_0__inst_mult_8_335 ;
wire Xd_0__inst_mult_8_339 ;
wire Xd_0__inst_mult_8_340 ;
wire Xd_0__inst_mult_11_334 ;
wire Xd_0__inst_mult_11_335 ;
wire Xd_0__inst_mult_11_339 ;
wire Xd_0__inst_mult_11_340 ;
wire Xd_0__inst_mult_10_334 ;
wire Xd_0__inst_mult_10_335 ;
wire Xd_0__inst_mult_10_339 ;
wire Xd_0__inst_mult_10_340 ;
wire Xd_0__inst_mult_5_334 ;
wire Xd_0__inst_mult_5_335 ;
wire Xd_0__inst_mult_5_339 ;
wire Xd_0__inst_mult_5_340 ;
wire Xd_0__inst_mult_4_334 ;
wire Xd_0__inst_mult_4_335 ;
wire Xd_0__inst_mult_4_339 ;
wire Xd_0__inst_mult_4_340 ;
wire Xd_0__inst_mult_7_334 ;
wire Xd_0__inst_mult_7_335 ;
wire Xd_0__inst_mult_7_339 ;
wire Xd_0__inst_mult_7_340 ;
wire Xd_0__inst_mult_6_334 ;
wire Xd_0__inst_mult_6_335 ;
wire Xd_0__inst_mult_6_339 ;
wire Xd_0__inst_mult_6_340 ;
wire Xd_0__inst_mult_1_334 ;
wire Xd_0__inst_mult_1_335 ;
wire Xd_0__inst_mult_1_339 ;
wire Xd_0__inst_mult_1_340 ;
wire Xd_0__inst_mult_0_334 ;
wire Xd_0__inst_mult_0_335 ;
wire Xd_0__inst_mult_0_339 ;
wire Xd_0__inst_mult_0_340 ;
wire Xd_0__inst_mult_3_334 ;
wire Xd_0__inst_mult_3_335 ;
wire Xd_0__inst_mult_3_339 ;
wire Xd_0__inst_mult_3_340 ;
wire Xd_0__inst_mult_15_65_sumout ;
wire Xd_0__inst_mult_15_66 ;
wire Xd_0__inst_mult_2_394 ;
wire Xd_0__inst_mult_2_395 ;
wire Xd_0__inst_mult_2_399 ;
wire Xd_0__inst_mult_2_400 ;
wire Xd_0__inst_mult_18_55_sumout ;
wire Xd_0__inst_mult_18_56 ;
wire Xd_0__inst_mult_29_384 ;
wire Xd_0__inst_mult_29_385 ;
wire Xd_0__inst_mult_29_389 ;
wire Xd_0__inst_mult_29_390 ;
wire Xd_0__inst_mult_28_344 ;
wire Xd_0__inst_mult_28_345 ;
wire Xd_0__inst_mult_28_349 ;
wire Xd_0__inst_mult_28_350 ;
wire Xd_0__inst_mult_31_344 ;
wire Xd_0__inst_mult_31_345 ;
wire Xd_0__inst_mult_31_349 ;
wire Xd_0__inst_mult_31_350 ;
wire Xd_0__inst_mult_30_344 ;
wire Xd_0__inst_mult_30_345 ;
wire Xd_0__inst_mult_30_349 ;
wire Xd_0__inst_mult_30_350 ;
wire Xd_0__inst_mult_25_444 ;
wire Xd_0__inst_mult_25_445 ;
wire Xd_0__inst_mult_25_449 ;
wire Xd_0__inst_mult_25_450 ;
wire Xd_0__inst_mult_24_634 ;
wire Xd_0__inst_mult_24_635 ;
wire Xd_0__inst_mult_24_639 ;
wire Xd_0__inst_mult_24_640 ;
wire Xd_0__inst_mult_27_444 ;
wire Xd_0__inst_mult_27_445 ;
wire Xd_0__inst_mult_27_449 ;
wire Xd_0__inst_mult_27_450 ;
wire Xd_0__inst_mult_26_634 ;
wire Xd_0__inst_mult_26_635 ;
wire Xd_0__inst_mult_26_639 ;
wire Xd_0__inst_mult_26_640 ;
wire Xd_0__inst_mult_21_384 ;
wire Xd_0__inst_mult_21_385 ;
wire Xd_0__inst_mult_21_389 ;
wire Xd_0__inst_mult_21_390 ;
wire Xd_0__inst_mult_20_384 ;
wire Xd_0__inst_mult_20_385 ;
wire Xd_0__inst_mult_20_389 ;
wire Xd_0__inst_mult_20_390 ;
wire Xd_0__inst_mult_23_384 ;
wire Xd_0__inst_mult_23_385 ;
wire Xd_0__inst_mult_23_389 ;
wire Xd_0__inst_mult_23_390 ;
wire Xd_0__inst_mult_22_384 ;
wire Xd_0__inst_mult_22_385 ;
wire Xd_0__inst_mult_22_389 ;
wire Xd_0__inst_mult_22_390 ;
wire Xd_0__inst_mult_17_384 ;
wire Xd_0__inst_mult_17_385 ;
wire Xd_0__inst_mult_17_389 ;
wire Xd_0__inst_mult_17_390 ;
wire Xd_0__inst_mult_16_384 ;
wire Xd_0__inst_mult_16_385 ;
wire Xd_0__inst_mult_16_389 ;
wire Xd_0__inst_mult_16_390 ;
wire Xd_0__inst_mult_19_384 ;
wire Xd_0__inst_mult_19_385 ;
wire Xd_0__inst_mult_19_389 ;
wire Xd_0__inst_mult_19_390 ;
wire Xd_0__inst_mult_18_319 ;
wire Xd_0__inst_mult_18_320 ;
wire Xd_0__inst_mult_18_324 ;
wire Xd_0__inst_mult_18_325 ;
wire Xd_0__inst_mult_13_344 ;
wire Xd_0__inst_mult_13_345 ;
wire Xd_0__inst_mult_13_349 ;
wire Xd_0__inst_mult_13_350 ;
wire Xd_0__inst_mult_12_319 ;
wire Xd_0__inst_mult_12_320 ;
wire Xd_0__inst_mult_12_324 ;
wire Xd_0__inst_mult_12_325 ;
wire Xd_0__inst_mult_15_319 ;
wire Xd_0__inst_mult_15_320 ;
wire Xd_0__inst_mult_15_324 ;
wire Xd_0__inst_mult_15_325 ;
wire Xd_0__inst_mult_14_319 ;
wire Xd_0__inst_mult_14_320 ;
wire Xd_0__inst_mult_14_324 ;
wire Xd_0__inst_mult_14_325 ;
wire Xd_0__inst_mult_9_344 ;
wire Xd_0__inst_mult_9_345 ;
wire Xd_0__inst_mult_9_349 ;
wire Xd_0__inst_mult_9_350 ;
wire Xd_0__inst_mult_8_344 ;
wire Xd_0__inst_mult_8_345 ;
wire Xd_0__inst_mult_8_349 ;
wire Xd_0__inst_mult_8_350 ;
wire Xd_0__inst_mult_11_344 ;
wire Xd_0__inst_mult_11_345 ;
wire Xd_0__inst_mult_11_349 ;
wire Xd_0__inst_mult_11_350 ;
wire Xd_0__inst_mult_10_344 ;
wire Xd_0__inst_mult_10_345 ;
wire Xd_0__inst_mult_10_349 ;
wire Xd_0__inst_mult_10_350 ;
wire Xd_0__inst_mult_5_344 ;
wire Xd_0__inst_mult_5_345 ;
wire Xd_0__inst_mult_5_349 ;
wire Xd_0__inst_mult_5_350 ;
wire Xd_0__inst_mult_4_344 ;
wire Xd_0__inst_mult_4_345 ;
wire Xd_0__inst_mult_4_349 ;
wire Xd_0__inst_mult_4_350 ;
wire Xd_0__inst_mult_7_344 ;
wire Xd_0__inst_mult_7_345 ;
wire Xd_0__inst_mult_7_349 ;
wire Xd_0__inst_mult_7_350 ;
wire Xd_0__inst_mult_6_344 ;
wire Xd_0__inst_mult_6_345 ;
wire Xd_0__inst_mult_6_349 ;
wire Xd_0__inst_mult_6_350 ;
wire Xd_0__inst_mult_1_344 ;
wire Xd_0__inst_mult_1_345 ;
wire Xd_0__inst_mult_1_349 ;
wire Xd_0__inst_mult_1_350 ;
wire Xd_0__inst_mult_0_344 ;
wire Xd_0__inst_mult_0_345 ;
wire Xd_0__inst_mult_0_349 ;
wire Xd_0__inst_mult_0_350 ;
wire Xd_0__inst_mult_3_344 ;
wire Xd_0__inst_mult_3_345 ;
wire Xd_0__inst_mult_3_349 ;
wire Xd_0__inst_mult_3_350 ;
wire Xd_0__inst_mult_2_404 ;
wire Xd_0__inst_mult_2_405 ;
wire Xd_0__inst_mult_2_409 ;
wire Xd_0__inst_mult_2_410 ;
wire Xd_0__inst_mult_29_394 ;
wire Xd_0__inst_mult_29_395 ;
wire Xd_0__inst_mult_29_399 ;
wire Xd_0__inst_mult_29_400 ;
wire Xd_0__inst_mult_28_354 ;
wire Xd_0__inst_mult_28_355 ;
wire Xd_0__inst_mult_28_359 ;
wire Xd_0__inst_mult_28_360 ;
wire Xd_0__inst_mult_31_354 ;
wire Xd_0__inst_mult_31_355 ;
wire Xd_0__inst_mult_31_359 ;
wire Xd_0__inst_mult_31_360 ;
wire Xd_0__inst_mult_30_354 ;
wire Xd_0__inst_mult_30_355 ;
wire Xd_0__inst_mult_30_359 ;
wire Xd_0__inst_mult_30_360 ;
wire Xd_0__inst_mult_25_454 ;
wire Xd_0__inst_mult_25_455 ;
wire Xd_0__inst_mult_25_459 ;
wire Xd_0__inst_mult_25_460 ;
wire Xd_0__inst_mult_24_644 ;
wire Xd_0__inst_mult_24_645 ;
wire Xd_0__inst_mult_24_649 ;
wire Xd_0__inst_mult_24_650 ;
wire Xd_0__inst_mult_27_454 ;
wire Xd_0__inst_mult_27_455 ;
wire Xd_0__inst_mult_27_459 ;
wire Xd_0__inst_mult_27_460 ;
wire Xd_0__inst_mult_26_644 ;
wire Xd_0__inst_mult_26_645 ;
wire Xd_0__inst_mult_26_649 ;
wire Xd_0__inst_mult_26_650 ;
wire Xd_0__inst_mult_21_394 ;
wire Xd_0__inst_mult_21_395 ;
wire Xd_0__inst_mult_21_399 ;
wire Xd_0__inst_mult_21_400 ;
wire Xd_0__inst_mult_20_394 ;
wire Xd_0__inst_mult_20_395 ;
wire Xd_0__inst_mult_20_399 ;
wire Xd_0__inst_mult_20_400 ;
wire Xd_0__inst_mult_23_394 ;
wire Xd_0__inst_mult_23_395 ;
wire Xd_0__inst_mult_23_399 ;
wire Xd_0__inst_mult_23_400 ;
wire Xd_0__inst_mult_22_394 ;
wire Xd_0__inst_mult_22_395 ;
wire Xd_0__inst_mult_22_399 ;
wire Xd_0__inst_mult_22_400 ;
wire Xd_0__inst_mult_17_394 ;
wire Xd_0__inst_mult_17_395 ;
wire Xd_0__inst_mult_17_399 ;
wire Xd_0__inst_mult_17_400 ;
wire Xd_0__inst_mult_16_394 ;
wire Xd_0__inst_mult_16_395 ;
wire Xd_0__inst_mult_16_399 ;
wire Xd_0__inst_mult_16_400 ;
wire Xd_0__inst_mult_19_394 ;
wire Xd_0__inst_mult_19_395 ;
wire Xd_0__inst_mult_19_399 ;
wire Xd_0__inst_mult_19_400 ;
wire Xd_0__inst_mult_18_329 ;
wire Xd_0__inst_mult_18_330 ;
wire Xd_0__inst_mult_18_334 ;
wire Xd_0__inst_mult_18_335 ;
wire Xd_0__inst_mult_13_354 ;
wire Xd_0__inst_mult_13_355 ;
wire Xd_0__inst_mult_13_359 ;
wire Xd_0__inst_mult_13_360 ;
wire Xd_0__inst_mult_12_329 ;
wire Xd_0__inst_mult_12_330 ;
wire Xd_0__inst_mult_12_334 ;
wire Xd_0__inst_mult_12_335 ;
wire Xd_0__inst_mult_15_329 ;
wire Xd_0__inst_mult_15_330 ;
wire Xd_0__inst_mult_15_334 ;
wire Xd_0__inst_mult_15_335 ;
wire Xd_0__inst_mult_14_329 ;
wire Xd_0__inst_mult_14_330 ;
wire Xd_0__inst_mult_14_334 ;
wire Xd_0__inst_mult_14_335 ;
wire Xd_0__inst_mult_9_354 ;
wire Xd_0__inst_mult_9_355 ;
wire Xd_0__inst_mult_9_359 ;
wire Xd_0__inst_mult_9_360 ;
wire Xd_0__inst_mult_8_354 ;
wire Xd_0__inst_mult_8_355 ;
wire Xd_0__inst_mult_8_359 ;
wire Xd_0__inst_mult_8_360 ;
wire Xd_0__inst_mult_11_354 ;
wire Xd_0__inst_mult_11_355 ;
wire Xd_0__inst_mult_11_359 ;
wire Xd_0__inst_mult_11_360 ;
wire Xd_0__inst_mult_10_354 ;
wire Xd_0__inst_mult_10_355 ;
wire Xd_0__inst_mult_10_359 ;
wire Xd_0__inst_mult_10_360 ;
wire Xd_0__inst_mult_5_354 ;
wire Xd_0__inst_mult_5_355 ;
wire Xd_0__inst_mult_5_359 ;
wire Xd_0__inst_mult_5_360 ;
wire Xd_0__inst_mult_4_354 ;
wire Xd_0__inst_mult_4_355 ;
wire Xd_0__inst_mult_4_359 ;
wire Xd_0__inst_mult_4_360 ;
wire Xd_0__inst_mult_7_354 ;
wire Xd_0__inst_mult_7_355 ;
wire Xd_0__inst_mult_7_359 ;
wire Xd_0__inst_mult_7_360 ;
wire Xd_0__inst_mult_6_354 ;
wire Xd_0__inst_mult_6_355 ;
wire Xd_0__inst_mult_6_359 ;
wire Xd_0__inst_mult_6_360 ;
wire Xd_0__inst_mult_1_354 ;
wire Xd_0__inst_mult_1_355 ;
wire Xd_0__inst_mult_1_359 ;
wire Xd_0__inst_mult_1_360 ;
wire Xd_0__inst_mult_0_354 ;
wire Xd_0__inst_mult_0_355 ;
wire Xd_0__inst_mult_0_359 ;
wire Xd_0__inst_mult_0_360 ;
wire Xd_0__inst_mult_3_354 ;
wire Xd_0__inst_mult_3_355 ;
wire Xd_0__inst_mult_3_359 ;
wire Xd_0__inst_mult_3_360 ;
wire Xd_0__inst_mult_2_414 ;
wire Xd_0__inst_mult_2_415 ;
wire Xd_0__inst_mult_2_419 ;
wire Xd_0__inst_mult_2_420 ;
wire Xd_0__inst_mult_29_404 ;
wire Xd_0__inst_mult_29_405 ;
wire Xd_0__inst_mult_29_409 ;
wire Xd_0__inst_mult_29_410 ;
wire Xd_0__inst_mult_19_50_sumout ;
wire Xd_0__inst_mult_19_51 ;
wire Xd_0__inst_mult_28_364 ;
wire Xd_0__inst_mult_28_365 ;
wire Xd_0__inst_mult_28_369 ;
wire Xd_0__inst_mult_28_370 ;
wire Xd_0__inst_mult_22_50_sumout ;
wire Xd_0__inst_mult_22_51 ;
wire Xd_0__inst_mult_31_364 ;
wire Xd_0__inst_mult_31_365 ;
wire Xd_0__inst_mult_31_369 ;
wire Xd_0__inst_mult_31_370 ;
wire Xd_0__inst_mult_21_50_sumout ;
wire Xd_0__inst_mult_21_51 ;
wire Xd_0__inst_mult_30_364 ;
wire Xd_0__inst_mult_30_365 ;
wire Xd_0__inst_mult_30_369 ;
wire Xd_0__inst_mult_30_370 ;
wire Xd_0__inst_mult_20_60_sumout ;
wire Xd_0__inst_mult_20_61 ;
wire Xd_0__inst_mult_25_464 ;
wire Xd_0__inst_mult_25_465 ;
wire Xd_0__inst_mult_25_469 ;
wire Xd_0__inst_mult_25_470 ;
wire Xd_0__inst_mult_24_654 ;
wire Xd_0__inst_mult_24_655 ;
wire Xd_0__inst_mult_24_659 ;
wire Xd_0__inst_mult_24_660 ;
wire Xd_0__inst_mult_30_50_sumout ;
wire Xd_0__inst_mult_30_51 ;
wire Xd_0__inst_mult_27_464 ;
wire Xd_0__inst_mult_27_465 ;
wire Xd_0__inst_mult_27_469 ;
wire Xd_0__inst_mult_27_470 ;
wire Xd_0__inst_mult_29_50_sumout ;
wire Xd_0__inst_mult_29_51 ;
wire Xd_0__inst_mult_26_654 ;
wire Xd_0__inst_mult_26_655 ;
wire Xd_0__inst_mult_26_659 ;
wire Xd_0__inst_mult_26_660 ;
wire Xd_0__inst_mult_0_50_sumout ;
wire Xd_0__inst_mult_0_51 ;
wire Xd_0__inst_mult_21_404 ;
wire Xd_0__inst_mult_21_405 ;
wire Xd_0__inst_mult_21_409 ;
wire Xd_0__inst_mult_21_410 ;
wire Xd_0__inst_mult_7_50_sumout ;
wire Xd_0__inst_mult_7_51 ;
wire Xd_0__inst_mult_20_404 ;
wire Xd_0__inst_mult_20_405 ;
wire Xd_0__inst_mult_20_409 ;
wire Xd_0__inst_mult_20_410 ;
wire Xd_0__inst_mult_9_50_sumout ;
wire Xd_0__inst_mult_9_51 ;
wire Xd_0__inst_mult_23_404 ;
wire Xd_0__inst_mult_23_405 ;
wire Xd_0__inst_mult_23_409 ;
wire Xd_0__inst_mult_23_410 ;
wire Xd_0__inst_mult_8_65_sumout ;
wire Xd_0__inst_mult_8_66 ;
wire Xd_0__inst_mult_22_404 ;
wire Xd_0__inst_mult_22_405 ;
wire Xd_0__inst_mult_22_409 ;
wire Xd_0__inst_mult_22_410 ;
wire Xd_0__inst_mult_17_404 ;
wire Xd_0__inst_mult_17_405 ;
wire Xd_0__inst_mult_17_409 ;
wire Xd_0__inst_mult_17_410 ;
wire Xd_0__inst_mult_10_50_sumout ;
wire Xd_0__inst_mult_10_51 ;
wire Xd_0__inst_mult_16_404 ;
wire Xd_0__inst_mult_16_405 ;
wire Xd_0__inst_mult_16_409 ;
wire Xd_0__inst_mult_16_410 ;
wire Xd_0__inst_mult_3_65_sumout ;
wire Xd_0__inst_mult_3_66 ;
wire Xd_0__inst_mult_19_404 ;
wire Xd_0__inst_mult_19_405 ;
wire Xd_0__inst_mult_19_409 ;
wire Xd_0__inst_mult_19_410 ;
wire Xd_0__inst_mult_6_60_sumout ;
wire Xd_0__inst_mult_6_61 ;
wire Xd_0__inst_mult_18_339 ;
wire Xd_0__inst_mult_18_340 ;
wire Xd_0__inst_mult_18_344 ;
wire Xd_0__inst_mult_18_345 ;
wire Xd_0__inst_mult_13_364 ;
wire Xd_0__inst_mult_13_365 ;
wire Xd_0__inst_mult_13_369 ;
wire Xd_0__inst_mult_13_370 ;
wire Xd_0__inst_mult_12_339 ;
wire Xd_0__inst_mult_12_340 ;
wire Xd_0__inst_mult_12_344 ;
wire Xd_0__inst_mult_12_345 ;
wire Xd_0__inst_mult_15_339 ;
wire Xd_0__inst_mult_15_340 ;
wire Xd_0__inst_mult_15_344 ;
wire Xd_0__inst_mult_15_345 ;
wire Xd_0__inst_mult_14_339 ;
wire Xd_0__inst_mult_14_340 ;
wire Xd_0__inst_mult_14_344 ;
wire Xd_0__inst_mult_14_345 ;
wire Xd_0__inst_mult_9_364 ;
wire Xd_0__inst_mult_9_365 ;
wire Xd_0__inst_mult_9_369 ;
wire Xd_0__inst_mult_9_370 ;
wire Xd_0__inst_mult_8_364 ;
wire Xd_0__inst_mult_8_365 ;
wire Xd_0__inst_mult_8_369 ;
wire Xd_0__inst_mult_8_370 ;
wire Xd_0__inst_mult_11_364 ;
wire Xd_0__inst_mult_11_365 ;
wire Xd_0__inst_mult_11_369 ;
wire Xd_0__inst_mult_11_370 ;
wire Xd_0__inst_mult_10_364 ;
wire Xd_0__inst_mult_10_365 ;
wire Xd_0__inst_mult_10_369 ;
wire Xd_0__inst_mult_10_370 ;
wire Xd_0__inst_mult_30_55_sumout ;
wire Xd_0__inst_mult_30_56 ;
wire Xd_0__inst_mult_5_364 ;
wire Xd_0__inst_mult_5_365 ;
wire Xd_0__inst_mult_5_369 ;
wire Xd_0__inst_mult_5_370 ;
wire Xd_0__inst_mult_29_55_sumout ;
wire Xd_0__inst_mult_29_56 ;
wire Xd_0__inst_mult_4_364 ;
wire Xd_0__inst_mult_4_365 ;
wire Xd_0__inst_mult_4_369 ;
wire Xd_0__inst_mult_4_370 ;
wire Xd_0__inst_mult_0_55_sumout ;
wire Xd_0__inst_mult_0_56 ;
wire Xd_0__inst_mult_7_364 ;
wire Xd_0__inst_mult_7_365 ;
wire Xd_0__inst_mult_7_369 ;
wire Xd_0__inst_mult_7_370 ;
wire Xd_0__inst_mult_7_55_sumout ;
wire Xd_0__inst_mult_7_56 ;
wire Xd_0__inst_mult_6_364 ;
wire Xd_0__inst_mult_6_365 ;
wire Xd_0__inst_mult_6_369 ;
wire Xd_0__inst_mult_6_370 ;
wire Xd_0__inst_mult_10_55_sumout ;
wire Xd_0__inst_mult_10_56 ;
wire Xd_0__inst_mult_1_364 ;
wire Xd_0__inst_mult_1_365 ;
wire Xd_0__inst_mult_1_369 ;
wire Xd_0__inst_mult_1_370 ;
wire Xd_0__inst_mult_9_55_sumout ;
wire Xd_0__inst_mult_9_56 ;
wire Xd_0__inst_mult_0_364 ;
wire Xd_0__inst_mult_0_365 ;
wire Xd_0__inst_mult_0_369 ;
wire Xd_0__inst_mult_0_370 ;
wire Xd_0__inst_mult_12_45_sumout ;
wire Xd_0__inst_mult_12_46 ;
wire Xd_0__inst_mult_3_364 ;
wire Xd_0__inst_mult_3_365 ;
wire Xd_0__inst_mult_3_369 ;
wire Xd_0__inst_mult_3_370 ;
wire Xd_0__inst_mult_7_60_sumout ;
wire Xd_0__inst_mult_7_61 ;
wire Xd_0__inst_mult_2_424 ;
wire Xd_0__inst_mult_2_425 ;
wire Xd_0__inst_mult_10_60_sumout ;
wire Xd_0__inst_mult_10_61 ;
wire Xd_0__inst_mult_29_414 ;
wire Xd_0__inst_mult_29_415 ;
wire Xd_0__inst_mult_29_419 ;
wire Xd_0__inst_mult_29_420 ;
wire Xd_0__inst_mult_28_374 ;
wire Xd_0__inst_mult_28_375 ;
wire Xd_0__inst_mult_28_379 ;
wire Xd_0__inst_mult_28_380 ;
wire Xd_0__inst_mult_31_374 ;
wire Xd_0__inst_mult_31_375 ;
wire Xd_0__inst_mult_31_379 ;
wire Xd_0__inst_mult_31_380 ;
wire Xd_0__inst_mult_30_374 ;
wire Xd_0__inst_mult_30_375 ;
wire Xd_0__inst_mult_30_379 ;
wire Xd_0__inst_mult_30_380 ;
wire Xd_0__inst_mult_25_474 ;
wire Xd_0__inst_mult_25_475 ;
wire Xd_0__inst_mult_25_479 ;
wire Xd_0__inst_mult_25_480 ;
wire Xd_0__inst_mult_24_664 ;
wire Xd_0__inst_mult_24_665 ;
wire Xd_0__inst_mult_24_669 ;
wire Xd_0__inst_mult_24_670 ;
wire Xd_0__inst_mult_27_474 ;
wire Xd_0__inst_mult_27_475 ;
wire Xd_0__inst_mult_27_479 ;
wire Xd_0__inst_mult_27_480 ;
wire Xd_0__inst_mult_26_664 ;
wire Xd_0__inst_mult_26_665 ;
wire Xd_0__inst_mult_26_669 ;
wire Xd_0__inst_mult_26_670 ;
wire Xd_0__inst_mult_21_414 ;
wire Xd_0__inst_mult_21_415 ;
wire Xd_0__inst_mult_21_419 ;
wire Xd_0__inst_mult_21_420 ;
wire Xd_0__inst_mult_20_414 ;
wire Xd_0__inst_mult_20_415 ;
wire Xd_0__inst_mult_20_419 ;
wire Xd_0__inst_mult_20_420 ;
wire Xd_0__inst_mult_23_414 ;
wire Xd_0__inst_mult_23_415 ;
wire Xd_0__inst_mult_23_419 ;
wire Xd_0__inst_mult_23_420 ;
wire Xd_0__inst_mult_22_414 ;
wire Xd_0__inst_mult_22_415 ;
wire Xd_0__inst_mult_22_419 ;
wire Xd_0__inst_mult_22_420 ;
wire Xd_0__inst_mult_17_414 ;
wire Xd_0__inst_mult_17_415 ;
wire Xd_0__inst_mult_17_419 ;
wire Xd_0__inst_mult_17_420 ;
wire Xd_0__inst_mult_16_414 ;
wire Xd_0__inst_mult_16_415 ;
wire Xd_0__inst_mult_16_419 ;
wire Xd_0__inst_mult_16_420 ;
wire Xd_0__inst_mult_19_414 ;
wire Xd_0__inst_mult_19_415 ;
wire Xd_0__inst_mult_19_419 ;
wire Xd_0__inst_mult_19_420 ;
wire Xd_0__inst_mult_18_349 ;
wire Xd_0__inst_mult_18_350 ;
wire Xd_0__inst_mult_18_354 ;
wire Xd_0__inst_mult_18_355 ;
wire Xd_0__inst_mult_13_374 ;
wire Xd_0__inst_mult_13_375 ;
wire Xd_0__inst_mult_13_379 ;
wire Xd_0__inst_mult_13_380 ;
wire Xd_0__inst_mult_12_349 ;
wire Xd_0__inst_mult_12_350 ;
wire Xd_0__inst_mult_12_354 ;
wire Xd_0__inst_mult_12_355 ;
wire Xd_0__inst_mult_15_349 ;
wire Xd_0__inst_mult_15_350 ;
wire Xd_0__inst_mult_15_354 ;
wire Xd_0__inst_mult_15_355 ;
wire Xd_0__inst_mult_14_349 ;
wire Xd_0__inst_mult_14_350 ;
wire Xd_0__inst_mult_14_354 ;
wire Xd_0__inst_mult_14_355 ;
wire Xd_0__inst_mult_9_374 ;
wire Xd_0__inst_mult_9_375 ;
wire Xd_0__inst_mult_9_379 ;
wire Xd_0__inst_mult_9_380 ;
wire Xd_0__inst_mult_8_374 ;
wire Xd_0__inst_mult_8_375 ;
wire Xd_0__inst_mult_8_379 ;
wire Xd_0__inst_mult_8_380 ;
wire Xd_0__inst_mult_11_374 ;
wire Xd_0__inst_mult_11_375 ;
wire Xd_0__inst_mult_11_379 ;
wire Xd_0__inst_mult_11_380 ;
wire Xd_0__inst_mult_10_374 ;
wire Xd_0__inst_mult_10_375 ;
wire Xd_0__inst_mult_10_379 ;
wire Xd_0__inst_mult_10_380 ;
wire Xd_0__inst_mult_5_374 ;
wire Xd_0__inst_mult_5_375 ;
wire Xd_0__inst_mult_5_379 ;
wire Xd_0__inst_mult_5_380 ;
wire Xd_0__inst_mult_4_374 ;
wire Xd_0__inst_mult_4_375 ;
wire Xd_0__inst_mult_4_379 ;
wire Xd_0__inst_mult_4_380 ;
wire Xd_0__inst_mult_7_374 ;
wire Xd_0__inst_mult_7_375 ;
wire Xd_0__inst_mult_7_379 ;
wire Xd_0__inst_mult_7_380 ;
wire Xd_0__inst_mult_6_374 ;
wire Xd_0__inst_mult_6_375 ;
wire Xd_0__inst_mult_6_379 ;
wire Xd_0__inst_mult_6_380 ;
wire Xd_0__inst_mult_1_374 ;
wire Xd_0__inst_mult_1_375 ;
wire Xd_0__inst_mult_1_379 ;
wire Xd_0__inst_mult_1_380 ;
wire Xd_0__inst_mult_0_374 ;
wire Xd_0__inst_mult_0_375 ;
wire Xd_0__inst_mult_0_379 ;
wire Xd_0__inst_mult_0_380 ;
wire Xd_0__inst_mult_3_374 ;
wire Xd_0__inst_mult_3_375 ;
wire Xd_0__inst_mult_3_379 ;
wire Xd_0__inst_mult_3_380 ;
wire Xd_0__inst_mult_2_429 ;
wire Xd_0__inst_mult_2_430 ;
wire Xd_0__inst_mult_29_424 ;
wire Xd_0__inst_mult_29_425 ;
wire Xd_0__inst_mult_29_429 ;
wire Xd_0__inst_mult_29_430 ;
wire Xd_0__inst_mult_28_384 ;
wire Xd_0__inst_mult_28_385 ;
wire Xd_0__inst_mult_28_389 ;
wire Xd_0__inst_mult_28_390 ;
wire Xd_0__inst_mult_31_384 ;
wire Xd_0__inst_mult_31_385 ;
wire Xd_0__inst_mult_31_389 ;
wire Xd_0__inst_mult_31_390 ;
wire Xd_0__inst_mult_30_384 ;
wire Xd_0__inst_mult_30_385 ;
wire Xd_0__inst_mult_30_389 ;
wire Xd_0__inst_mult_30_390 ;
wire Xd_0__inst_mult_25_484 ;
wire Xd_0__inst_mult_25_485 ;
wire Xd_0__inst_mult_25_489 ;
wire Xd_0__inst_mult_25_490 ;
wire Xd_0__inst_mult_24_674 ;
wire Xd_0__inst_mult_24_675 ;
wire Xd_0__inst_mult_24_679 ;
wire Xd_0__inst_mult_24_680 ;
wire Xd_0__inst_mult_27_484 ;
wire Xd_0__inst_mult_27_485 ;
wire Xd_0__inst_mult_27_489 ;
wire Xd_0__inst_mult_27_490 ;
wire Xd_0__inst_mult_26_674 ;
wire Xd_0__inst_mult_26_675 ;
wire Xd_0__inst_mult_26_679 ;
wire Xd_0__inst_mult_26_680 ;
wire Xd_0__inst_mult_21_424 ;
wire Xd_0__inst_mult_21_425 ;
wire Xd_0__inst_mult_21_429 ;
wire Xd_0__inst_mult_21_430 ;
wire Xd_0__inst_mult_20_424 ;
wire Xd_0__inst_mult_20_425 ;
wire Xd_0__inst_mult_20_429 ;
wire Xd_0__inst_mult_20_430 ;
wire Xd_0__inst_mult_23_424 ;
wire Xd_0__inst_mult_23_425 ;
wire Xd_0__inst_mult_23_429 ;
wire Xd_0__inst_mult_23_430 ;
wire Xd_0__inst_mult_22_424 ;
wire Xd_0__inst_mult_22_425 ;
wire Xd_0__inst_mult_22_429 ;
wire Xd_0__inst_mult_22_430 ;
wire Xd_0__inst_mult_17_424 ;
wire Xd_0__inst_mult_17_425 ;
wire Xd_0__inst_mult_17_429 ;
wire Xd_0__inst_mult_17_430 ;
wire Xd_0__inst_mult_16_424 ;
wire Xd_0__inst_mult_16_425 ;
wire Xd_0__inst_mult_16_429 ;
wire Xd_0__inst_mult_16_430 ;
wire Xd_0__inst_mult_19_424 ;
wire Xd_0__inst_mult_19_425 ;
wire Xd_0__inst_mult_19_429 ;
wire Xd_0__inst_mult_19_430 ;
wire Xd_0__inst_mult_18_359 ;
wire Xd_0__inst_mult_18_360 ;
wire Xd_0__inst_mult_18_364 ;
wire Xd_0__inst_mult_18_365 ;
wire Xd_0__inst_mult_13_384 ;
wire Xd_0__inst_mult_13_385 ;
wire Xd_0__inst_mult_13_389 ;
wire Xd_0__inst_mult_13_390 ;
wire Xd_0__inst_mult_12_359 ;
wire Xd_0__inst_mult_12_360 ;
wire Xd_0__inst_mult_12_364 ;
wire Xd_0__inst_mult_12_365 ;
wire Xd_0__inst_mult_15_359 ;
wire Xd_0__inst_mult_15_360 ;
wire Xd_0__inst_mult_15_364 ;
wire Xd_0__inst_mult_15_365 ;
wire Xd_0__inst_mult_14_359 ;
wire Xd_0__inst_mult_14_360 ;
wire Xd_0__inst_mult_14_364 ;
wire Xd_0__inst_mult_14_365 ;
wire Xd_0__inst_mult_9_384 ;
wire Xd_0__inst_mult_9_385 ;
wire Xd_0__inst_mult_9_389 ;
wire Xd_0__inst_mult_9_390 ;
wire Xd_0__inst_mult_8_384 ;
wire Xd_0__inst_mult_8_385 ;
wire Xd_0__inst_mult_8_389 ;
wire Xd_0__inst_mult_8_390 ;
wire Xd_0__inst_mult_11_384 ;
wire Xd_0__inst_mult_11_385 ;
wire Xd_0__inst_mult_11_389 ;
wire Xd_0__inst_mult_11_390 ;
wire Xd_0__inst_mult_10_384 ;
wire Xd_0__inst_mult_10_385 ;
wire Xd_0__inst_mult_10_389 ;
wire Xd_0__inst_mult_10_390 ;
wire Xd_0__inst_mult_5_384 ;
wire Xd_0__inst_mult_5_385 ;
wire Xd_0__inst_mult_5_389 ;
wire Xd_0__inst_mult_5_390 ;
wire Xd_0__inst_mult_4_384 ;
wire Xd_0__inst_mult_4_385 ;
wire Xd_0__inst_mult_4_389 ;
wire Xd_0__inst_mult_4_390 ;
wire Xd_0__inst_mult_7_384 ;
wire Xd_0__inst_mult_7_385 ;
wire Xd_0__inst_mult_7_389 ;
wire Xd_0__inst_mult_7_390 ;
wire Xd_0__inst_mult_6_384 ;
wire Xd_0__inst_mult_6_385 ;
wire Xd_0__inst_mult_6_389 ;
wire Xd_0__inst_mult_6_390 ;
wire Xd_0__inst_mult_1_384 ;
wire Xd_0__inst_mult_1_385 ;
wire Xd_0__inst_mult_1_389 ;
wire Xd_0__inst_mult_1_390 ;
wire Xd_0__inst_mult_0_384 ;
wire Xd_0__inst_mult_0_385 ;
wire Xd_0__inst_mult_0_389 ;
wire Xd_0__inst_mult_0_390 ;
wire Xd_0__inst_mult_3_384 ;
wire Xd_0__inst_mult_3_385 ;
wire Xd_0__inst_mult_3_389 ;
wire Xd_0__inst_mult_3_390 ;
wire Xd_0__inst_mult_2_434 ;
wire Xd_0__inst_mult_2_435 ;
wire Xd_0__inst_mult_29_434 ;
wire Xd_0__inst_mult_29_435 ;
wire Xd_0__inst_mult_29_439 ;
wire Xd_0__inst_mult_29_440 ;
wire Xd_0__inst_mult_28_394 ;
wire Xd_0__inst_mult_28_395 ;
wire Xd_0__inst_mult_28_399 ;
wire Xd_0__inst_mult_28_400 ;
wire Xd_0__inst_mult_31_394 ;
wire Xd_0__inst_mult_31_395 ;
wire Xd_0__inst_mult_31_399 ;
wire Xd_0__inst_mult_31_400 ;
wire Xd_0__inst_mult_30_394 ;
wire Xd_0__inst_mult_30_395 ;
wire Xd_0__inst_mult_30_399 ;
wire Xd_0__inst_mult_30_400 ;
wire Xd_0__inst_mult_25_494 ;
wire Xd_0__inst_mult_25_495 ;
wire Xd_0__inst_mult_24_684 ;
wire Xd_0__inst_mult_24_685 ;
wire Xd_0__inst_mult_27_494 ;
wire Xd_0__inst_mult_27_495 ;
wire Xd_0__inst_mult_26_684 ;
wire Xd_0__inst_mult_26_685 ;
wire Xd_0__inst_mult_21_434 ;
wire Xd_0__inst_mult_21_435 ;
wire Xd_0__inst_mult_21_439 ;
wire Xd_0__inst_mult_21_440 ;
wire Xd_0__inst_mult_20_434 ;
wire Xd_0__inst_mult_20_435 ;
wire Xd_0__inst_mult_20_439 ;
wire Xd_0__inst_mult_20_440 ;
wire Xd_0__inst_mult_23_434 ;
wire Xd_0__inst_mult_23_435 ;
wire Xd_0__inst_mult_23_439 ;
wire Xd_0__inst_mult_23_440 ;
wire Xd_0__inst_mult_22_434 ;
wire Xd_0__inst_mult_22_435 ;
wire Xd_0__inst_mult_22_439 ;
wire Xd_0__inst_mult_22_440 ;
wire Xd_0__inst_mult_17_434 ;
wire Xd_0__inst_mult_17_435 ;
wire Xd_0__inst_mult_17_439 ;
wire Xd_0__inst_mult_17_440 ;
wire Xd_0__inst_mult_16_434 ;
wire Xd_0__inst_mult_16_435 ;
wire Xd_0__inst_mult_16_439 ;
wire Xd_0__inst_mult_16_440 ;
wire Xd_0__inst_mult_19_434 ;
wire Xd_0__inst_mult_19_435 ;
wire Xd_0__inst_mult_19_439 ;
wire Xd_0__inst_mult_19_440 ;
wire Xd_0__inst_mult_18_369 ;
wire Xd_0__inst_mult_18_370 ;
wire Xd_0__inst_mult_18_374 ;
wire Xd_0__inst_mult_18_375 ;
wire Xd_0__inst_mult_13_394 ;
wire Xd_0__inst_mult_13_395 ;
wire Xd_0__inst_mult_13_399 ;
wire Xd_0__inst_mult_13_400 ;
wire Xd_0__inst_mult_12_369 ;
wire Xd_0__inst_mult_12_370 ;
wire Xd_0__inst_mult_12_374 ;
wire Xd_0__inst_mult_12_375 ;
wire Xd_0__inst_mult_15_369 ;
wire Xd_0__inst_mult_15_370 ;
wire Xd_0__inst_mult_15_374 ;
wire Xd_0__inst_mult_15_375 ;
wire Xd_0__inst_mult_14_369 ;
wire Xd_0__inst_mult_14_370 ;
wire Xd_0__inst_mult_14_374 ;
wire Xd_0__inst_mult_14_375 ;
wire Xd_0__inst_mult_9_394 ;
wire Xd_0__inst_mult_9_395 ;
wire Xd_0__inst_mult_9_399 ;
wire Xd_0__inst_mult_9_400 ;
wire Xd_0__inst_mult_8_394 ;
wire Xd_0__inst_mult_8_395 ;
wire Xd_0__inst_mult_8_399 ;
wire Xd_0__inst_mult_8_400 ;
wire Xd_0__inst_mult_11_394 ;
wire Xd_0__inst_mult_11_395 ;
wire Xd_0__inst_mult_11_399 ;
wire Xd_0__inst_mult_11_400 ;
wire Xd_0__inst_mult_10_394 ;
wire Xd_0__inst_mult_10_395 ;
wire Xd_0__inst_mult_10_399 ;
wire Xd_0__inst_mult_10_400 ;
wire Xd_0__inst_mult_5_394 ;
wire Xd_0__inst_mult_5_395 ;
wire Xd_0__inst_mult_5_399 ;
wire Xd_0__inst_mult_5_400 ;
wire Xd_0__inst_mult_4_394 ;
wire Xd_0__inst_mult_4_395 ;
wire Xd_0__inst_mult_4_399 ;
wire Xd_0__inst_mult_4_400 ;
wire Xd_0__inst_mult_7_394 ;
wire Xd_0__inst_mult_7_395 ;
wire Xd_0__inst_mult_7_399 ;
wire Xd_0__inst_mult_7_400 ;
wire Xd_0__inst_mult_6_394 ;
wire Xd_0__inst_mult_6_395 ;
wire Xd_0__inst_mult_6_399 ;
wire Xd_0__inst_mult_6_400 ;
wire Xd_0__inst_mult_1_394 ;
wire Xd_0__inst_mult_1_395 ;
wire Xd_0__inst_mult_1_399 ;
wire Xd_0__inst_mult_1_400 ;
wire Xd_0__inst_mult_0_394 ;
wire Xd_0__inst_mult_0_395 ;
wire Xd_0__inst_mult_0_399 ;
wire Xd_0__inst_mult_0_400 ;
wire Xd_0__inst_mult_3_394 ;
wire Xd_0__inst_mult_3_395 ;
wire Xd_0__inst_mult_3_399 ;
wire Xd_0__inst_mult_3_400 ;
wire Xd_0__inst_mult_2_439 ;
wire Xd_0__inst_mult_2_440 ;
wire Xd_0__inst_mult_2_444 ;
wire Xd_0__inst_mult_2_445 ;
wire Xd_0__inst_mult_29_444 ;
wire Xd_0__inst_mult_29_445 ;
wire Xd_0__inst_mult_29_449 ;
wire Xd_0__inst_mult_29_450 ;
wire Xd_0__inst_mult_28_404 ;
wire Xd_0__inst_mult_28_405 ;
wire Xd_0__inst_mult_28_409 ;
wire Xd_0__inst_mult_28_410 ;
wire Xd_0__inst_mult_31_404 ;
wire Xd_0__inst_mult_31_405 ;
wire Xd_0__inst_mult_31_409 ;
wire Xd_0__inst_mult_31_410 ;
wire Xd_0__inst_mult_30_404 ;
wire Xd_0__inst_mult_30_405 ;
wire Xd_0__inst_mult_30_409 ;
wire Xd_0__inst_mult_30_410 ;
wire Xd_0__inst_mult_25_499 ;
wire Xd_0__inst_mult_25_500 ;
wire Xd_0__inst_mult_24_689 ;
wire Xd_0__inst_mult_24_690 ;
wire Xd_0__inst_mult_27_499 ;
wire Xd_0__inst_mult_27_500 ;
wire Xd_0__inst_mult_26_689 ;
wire Xd_0__inst_mult_26_690 ;
wire Xd_0__inst_mult_21_444 ;
wire Xd_0__inst_mult_21_445 ;
wire Xd_0__inst_mult_21_449 ;
wire Xd_0__inst_mult_21_450 ;
wire Xd_0__inst_mult_20_444 ;
wire Xd_0__inst_mult_20_445 ;
wire Xd_0__inst_mult_20_449 ;
wire Xd_0__inst_mult_20_450 ;
wire Xd_0__inst_mult_23_444 ;
wire Xd_0__inst_mult_23_445 ;
wire Xd_0__inst_mult_23_449 ;
wire Xd_0__inst_mult_23_450 ;
wire Xd_0__inst_mult_22_444 ;
wire Xd_0__inst_mult_22_445 ;
wire Xd_0__inst_mult_22_449 ;
wire Xd_0__inst_mult_22_450 ;
wire Xd_0__inst_mult_17_444 ;
wire Xd_0__inst_mult_17_445 ;
wire Xd_0__inst_mult_17_449 ;
wire Xd_0__inst_mult_17_450 ;
wire Xd_0__inst_mult_16_444 ;
wire Xd_0__inst_mult_16_445 ;
wire Xd_0__inst_mult_16_449 ;
wire Xd_0__inst_mult_16_450 ;
wire Xd_0__inst_mult_19_444 ;
wire Xd_0__inst_mult_19_445 ;
wire Xd_0__inst_mult_19_449 ;
wire Xd_0__inst_mult_19_450 ;
wire Xd_0__inst_mult_18_379 ;
wire Xd_0__inst_mult_18_380 ;
wire Xd_0__inst_mult_18_384 ;
wire Xd_0__inst_mult_18_385 ;
wire Xd_0__inst_mult_13_404 ;
wire Xd_0__inst_mult_13_405 ;
wire Xd_0__inst_mult_13_409 ;
wire Xd_0__inst_mult_13_410 ;
wire Xd_0__inst_mult_12_379 ;
wire Xd_0__inst_mult_12_380 ;
wire Xd_0__inst_mult_12_384 ;
wire Xd_0__inst_mult_12_385 ;
wire Xd_0__inst_mult_15_379 ;
wire Xd_0__inst_mult_15_380 ;
wire Xd_0__inst_mult_15_384 ;
wire Xd_0__inst_mult_15_385 ;
wire Xd_0__inst_mult_14_379 ;
wire Xd_0__inst_mult_14_380 ;
wire Xd_0__inst_mult_14_384 ;
wire Xd_0__inst_mult_14_385 ;
wire Xd_0__inst_mult_9_404 ;
wire Xd_0__inst_mult_9_405 ;
wire Xd_0__inst_mult_9_409 ;
wire Xd_0__inst_mult_9_410 ;
wire Xd_0__inst_mult_8_404 ;
wire Xd_0__inst_mult_8_405 ;
wire Xd_0__inst_mult_8_409 ;
wire Xd_0__inst_mult_8_410 ;
wire Xd_0__inst_mult_11_404 ;
wire Xd_0__inst_mult_11_405 ;
wire Xd_0__inst_mult_11_409 ;
wire Xd_0__inst_mult_11_410 ;
wire Xd_0__inst_mult_10_404 ;
wire Xd_0__inst_mult_10_405 ;
wire Xd_0__inst_mult_10_409 ;
wire Xd_0__inst_mult_10_410 ;
wire Xd_0__inst_mult_5_404 ;
wire Xd_0__inst_mult_5_405 ;
wire Xd_0__inst_mult_5_409 ;
wire Xd_0__inst_mult_5_410 ;
wire Xd_0__inst_mult_4_404 ;
wire Xd_0__inst_mult_4_405 ;
wire Xd_0__inst_mult_4_409 ;
wire Xd_0__inst_mult_4_410 ;
wire Xd_0__inst_mult_7_404 ;
wire Xd_0__inst_mult_7_405 ;
wire Xd_0__inst_mult_7_409 ;
wire Xd_0__inst_mult_7_410 ;
wire Xd_0__inst_mult_6_404 ;
wire Xd_0__inst_mult_6_405 ;
wire Xd_0__inst_mult_6_409 ;
wire Xd_0__inst_mult_6_410 ;
wire Xd_0__inst_mult_1_404 ;
wire Xd_0__inst_mult_1_405 ;
wire Xd_0__inst_mult_1_409 ;
wire Xd_0__inst_mult_1_410 ;
wire Xd_0__inst_mult_0_404 ;
wire Xd_0__inst_mult_0_405 ;
wire Xd_0__inst_mult_0_409 ;
wire Xd_0__inst_mult_0_410 ;
wire Xd_0__inst_mult_3_404 ;
wire Xd_0__inst_mult_3_405 ;
wire Xd_0__inst_mult_3_409 ;
wire Xd_0__inst_mult_3_410 ;
wire Xd_0__inst_mult_2_449 ;
wire Xd_0__inst_mult_2_450 ;
wire Xd_0__inst_mult_2_454 ;
wire Xd_0__inst_mult_2_455 ;
wire Xd_0__inst_mult_29_454 ;
wire Xd_0__inst_mult_29_455 ;
wire Xd_0__inst_mult_29_459 ;
wire Xd_0__inst_mult_29_460 ;
wire Xd_0__inst_mult_28_414 ;
wire Xd_0__inst_mult_28_415 ;
wire Xd_0__inst_mult_28_419 ;
wire Xd_0__inst_mult_28_420 ;
wire Xd_0__inst_mult_31_414 ;
wire Xd_0__inst_mult_31_415 ;
wire Xd_0__inst_mult_31_419 ;
wire Xd_0__inst_mult_31_420 ;
wire Xd_0__inst_mult_30_414 ;
wire Xd_0__inst_mult_30_415 ;
wire Xd_0__inst_mult_30_419 ;
wire Xd_0__inst_mult_30_420 ;
wire Xd_0__inst_mult_25_504 ;
wire Xd_0__inst_mult_25_505 ;
wire Xd_0__inst_mult_24_694 ;
wire Xd_0__inst_mult_24_695 ;
wire Xd_0__inst_mult_27_504 ;
wire Xd_0__inst_mult_27_505 ;
wire Xd_0__inst_mult_26_694 ;
wire Xd_0__inst_mult_26_695 ;
wire Xd_0__inst_mult_21_454 ;
wire Xd_0__inst_mult_21_455 ;
wire Xd_0__inst_mult_21_459 ;
wire Xd_0__inst_mult_21_460 ;
wire Xd_0__inst_mult_20_454 ;
wire Xd_0__inst_mult_20_455 ;
wire Xd_0__inst_mult_20_459 ;
wire Xd_0__inst_mult_20_460 ;
wire Xd_0__inst_mult_23_454 ;
wire Xd_0__inst_mult_23_455 ;
wire Xd_0__inst_mult_23_459 ;
wire Xd_0__inst_mult_23_460 ;
wire Xd_0__inst_mult_22_454 ;
wire Xd_0__inst_mult_22_455 ;
wire Xd_0__inst_mult_22_459 ;
wire Xd_0__inst_mult_22_460 ;
wire Xd_0__inst_mult_17_454 ;
wire Xd_0__inst_mult_17_455 ;
wire Xd_0__inst_mult_17_459 ;
wire Xd_0__inst_mult_17_460 ;
wire Xd_0__inst_mult_16_454 ;
wire Xd_0__inst_mult_16_455 ;
wire Xd_0__inst_mult_16_459 ;
wire Xd_0__inst_mult_16_460 ;
wire Xd_0__inst_mult_19_454 ;
wire Xd_0__inst_mult_19_455 ;
wire Xd_0__inst_mult_19_459 ;
wire Xd_0__inst_mult_19_460 ;
wire Xd_0__inst_mult_18_389 ;
wire Xd_0__inst_mult_18_390 ;
wire Xd_0__inst_mult_18_394 ;
wire Xd_0__inst_mult_18_395 ;
wire Xd_0__inst_mult_13_414 ;
wire Xd_0__inst_mult_13_415 ;
wire Xd_0__inst_mult_13_419 ;
wire Xd_0__inst_mult_13_420 ;
wire Xd_0__inst_mult_12_389 ;
wire Xd_0__inst_mult_12_390 ;
wire Xd_0__inst_mult_12_394 ;
wire Xd_0__inst_mult_12_395 ;
wire Xd_0__inst_mult_15_389 ;
wire Xd_0__inst_mult_15_390 ;
wire Xd_0__inst_mult_15_394 ;
wire Xd_0__inst_mult_15_395 ;
wire Xd_0__inst_mult_14_389 ;
wire Xd_0__inst_mult_14_390 ;
wire Xd_0__inst_mult_14_394 ;
wire Xd_0__inst_mult_14_395 ;
wire Xd_0__inst_mult_9_414 ;
wire Xd_0__inst_mult_9_415 ;
wire Xd_0__inst_mult_9_419 ;
wire Xd_0__inst_mult_9_420 ;
wire Xd_0__inst_mult_8_414 ;
wire Xd_0__inst_mult_8_415 ;
wire Xd_0__inst_mult_8_419 ;
wire Xd_0__inst_mult_8_420 ;
wire Xd_0__inst_mult_11_414 ;
wire Xd_0__inst_mult_11_415 ;
wire Xd_0__inst_mult_11_419 ;
wire Xd_0__inst_mult_11_420 ;
wire Xd_0__inst_mult_10_414 ;
wire Xd_0__inst_mult_10_415 ;
wire Xd_0__inst_mult_10_419 ;
wire Xd_0__inst_mult_10_420 ;
wire Xd_0__inst_mult_5_414 ;
wire Xd_0__inst_mult_5_415 ;
wire Xd_0__inst_mult_5_419 ;
wire Xd_0__inst_mult_5_420 ;
wire Xd_0__inst_mult_4_414 ;
wire Xd_0__inst_mult_4_415 ;
wire Xd_0__inst_mult_4_419 ;
wire Xd_0__inst_mult_4_420 ;
wire Xd_0__inst_mult_7_414 ;
wire Xd_0__inst_mult_7_415 ;
wire Xd_0__inst_mult_7_419 ;
wire Xd_0__inst_mult_7_420 ;
wire Xd_0__inst_mult_6_414 ;
wire Xd_0__inst_mult_6_415 ;
wire Xd_0__inst_mult_6_419 ;
wire Xd_0__inst_mult_6_420 ;
wire Xd_0__inst_mult_1_414 ;
wire Xd_0__inst_mult_1_415 ;
wire Xd_0__inst_mult_1_419 ;
wire Xd_0__inst_mult_1_420 ;
wire Xd_0__inst_mult_0_414 ;
wire Xd_0__inst_mult_0_415 ;
wire Xd_0__inst_mult_0_419 ;
wire Xd_0__inst_mult_0_420 ;
wire Xd_0__inst_mult_3_414 ;
wire Xd_0__inst_mult_3_415 ;
wire Xd_0__inst_mult_3_419 ;
wire Xd_0__inst_mult_3_420 ;
wire Xd_0__inst_mult_2_459 ;
wire Xd_0__inst_mult_2_460 ;
wire Xd_0__inst_mult_2_464 ;
wire Xd_0__inst_mult_2_465 ;
wire Xd_0__inst_mult_29_464 ;
wire Xd_0__inst_mult_29_465 ;
wire Xd_0__inst_mult_28_424 ;
wire Xd_0__inst_mult_28_425 ;
wire Xd_0__inst_mult_28_429 ;
wire Xd_0__inst_mult_28_430 ;
wire Xd_0__inst_mult_31_424 ;
wire Xd_0__inst_mult_31_425 ;
wire Xd_0__inst_mult_31_429 ;
wire Xd_0__inst_mult_31_430 ;
wire Xd_0__inst_mult_30_424 ;
wire Xd_0__inst_mult_30_425 ;
wire Xd_0__inst_mult_30_429 ;
wire Xd_0__inst_mult_30_430 ;
wire Xd_0__inst_mult_25_509 ;
wire Xd_0__inst_mult_25_510 ;
wire Xd_0__inst_mult_27_509 ;
wire Xd_0__inst_mult_27_510 ;
wire Xd_0__inst_mult_21_464 ;
wire Xd_0__inst_mult_21_465 ;
wire Xd_0__inst_mult_20_464 ;
wire Xd_0__inst_mult_20_465 ;
wire Xd_0__inst_mult_23_464 ;
wire Xd_0__inst_mult_23_465 ;
wire Xd_0__inst_mult_22_464 ;
wire Xd_0__inst_mult_22_465 ;
wire Xd_0__inst_mult_17_464 ;
wire Xd_0__inst_mult_17_465 ;
wire Xd_0__inst_mult_16_464 ;
wire Xd_0__inst_mult_16_465 ;
wire Xd_0__inst_mult_19_464 ;
wire Xd_0__inst_mult_19_465 ;
wire Xd_0__inst_mult_18_399 ;
wire Xd_0__inst_mult_18_400 ;
wire Xd_0__inst_mult_18_404 ;
wire Xd_0__inst_mult_18_405 ;
wire Xd_0__inst_mult_13_424 ;
wire Xd_0__inst_mult_13_425 ;
wire Xd_0__inst_mult_13_429 ;
wire Xd_0__inst_mult_13_430 ;
wire Xd_0__inst_mult_12_399 ;
wire Xd_0__inst_mult_12_400 ;
wire Xd_0__inst_mult_12_404 ;
wire Xd_0__inst_mult_12_405 ;
wire Xd_0__inst_mult_15_399 ;
wire Xd_0__inst_mult_15_400 ;
wire Xd_0__inst_mult_15_404 ;
wire Xd_0__inst_mult_15_405 ;
wire Xd_0__inst_mult_14_399 ;
wire Xd_0__inst_mult_14_400 ;
wire Xd_0__inst_mult_14_404 ;
wire Xd_0__inst_mult_14_405 ;
wire Xd_0__inst_mult_9_424 ;
wire Xd_0__inst_mult_9_425 ;
wire Xd_0__inst_mult_9_429 ;
wire Xd_0__inst_mult_9_430 ;
wire Xd_0__inst_mult_8_424 ;
wire Xd_0__inst_mult_8_425 ;
wire Xd_0__inst_mult_8_429 ;
wire Xd_0__inst_mult_8_430 ;
wire Xd_0__inst_mult_11_424 ;
wire Xd_0__inst_mult_11_425 ;
wire Xd_0__inst_mult_11_429 ;
wire Xd_0__inst_mult_11_430 ;
wire Xd_0__inst_mult_10_424 ;
wire Xd_0__inst_mult_10_425 ;
wire Xd_0__inst_mult_10_429 ;
wire Xd_0__inst_mult_10_430 ;
wire Xd_0__inst_mult_5_424 ;
wire Xd_0__inst_mult_5_425 ;
wire Xd_0__inst_mult_5_429 ;
wire Xd_0__inst_mult_5_430 ;
wire Xd_0__inst_mult_4_424 ;
wire Xd_0__inst_mult_4_425 ;
wire Xd_0__inst_mult_4_429 ;
wire Xd_0__inst_mult_4_430 ;
wire Xd_0__inst_mult_7_424 ;
wire Xd_0__inst_mult_7_425 ;
wire Xd_0__inst_mult_7_429 ;
wire Xd_0__inst_mult_7_430 ;
wire Xd_0__inst_mult_6_424 ;
wire Xd_0__inst_mult_6_425 ;
wire Xd_0__inst_mult_6_429 ;
wire Xd_0__inst_mult_6_430 ;
wire Xd_0__inst_mult_1_424 ;
wire Xd_0__inst_mult_1_425 ;
wire Xd_0__inst_mult_1_429 ;
wire Xd_0__inst_mult_1_430 ;
wire Xd_0__inst_mult_0_424 ;
wire Xd_0__inst_mult_0_425 ;
wire Xd_0__inst_mult_0_429 ;
wire Xd_0__inst_mult_0_430 ;
wire Xd_0__inst_mult_3_424 ;
wire Xd_0__inst_mult_3_425 ;
wire Xd_0__inst_mult_3_429 ;
wire Xd_0__inst_mult_3_430 ;
wire Xd_0__inst_mult_2_469 ;
wire Xd_0__inst_mult_2_470 ;
wire Xd_0__inst_mult_2_474 ;
wire Xd_0__inst_mult_2_475 ;
wire Xd_0__inst_mult_29_469 ;
wire Xd_0__inst_mult_29_470 ;
wire Xd_0__inst_mult_28_434 ;
wire Xd_0__inst_mult_28_435 ;
wire Xd_0__inst_mult_28_439 ;
wire Xd_0__inst_mult_28_440 ;
wire Xd_0__inst_mult_31_434 ;
wire Xd_0__inst_mult_31_435 ;
wire Xd_0__inst_mult_31_439 ;
wire Xd_0__inst_mult_31_440 ;
wire Xd_0__inst_mult_30_434 ;
wire Xd_0__inst_mult_30_435 ;
wire Xd_0__inst_mult_30_439 ;
wire Xd_0__inst_mult_30_440 ;
wire Xd_0__inst_mult_25_514 ;
wire Xd_0__inst_mult_25_515 ;
wire Xd_0__inst_mult_27_514 ;
wire Xd_0__inst_mult_27_515 ;
wire Xd_0__inst_mult_21_469 ;
wire Xd_0__inst_mult_21_470 ;
wire Xd_0__inst_mult_20_469 ;
wire Xd_0__inst_mult_20_470 ;
wire Xd_0__inst_mult_23_469 ;
wire Xd_0__inst_mult_23_470 ;
wire Xd_0__inst_mult_22_469 ;
wire Xd_0__inst_mult_22_470 ;
wire Xd_0__inst_mult_17_469 ;
wire Xd_0__inst_mult_17_470 ;
wire Xd_0__inst_mult_16_469 ;
wire Xd_0__inst_mult_16_470 ;
wire Xd_0__inst_mult_19_469 ;
wire Xd_0__inst_mult_19_470 ;
wire Xd_0__inst_mult_18_409 ;
wire Xd_0__inst_mult_18_410 ;
wire Xd_0__inst_mult_18_414 ;
wire Xd_0__inst_mult_18_415 ;
wire Xd_0__inst_mult_13_434 ;
wire Xd_0__inst_mult_13_435 ;
wire Xd_0__inst_mult_13_439 ;
wire Xd_0__inst_mult_13_440 ;
wire Xd_0__inst_mult_12_409 ;
wire Xd_0__inst_mult_12_410 ;
wire Xd_0__inst_mult_12_414 ;
wire Xd_0__inst_mult_12_415 ;
wire Xd_0__inst_mult_15_409 ;
wire Xd_0__inst_mult_15_410 ;
wire Xd_0__inst_mult_15_414 ;
wire Xd_0__inst_mult_15_415 ;
wire Xd_0__inst_mult_14_409 ;
wire Xd_0__inst_mult_14_410 ;
wire Xd_0__inst_mult_14_414 ;
wire Xd_0__inst_mult_14_415 ;
wire Xd_0__inst_mult_9_434 ;
wire Xd_0__inst_mult_9_435 ;
wire Xd_0__inst_mult_9_439 ;
wire Xd_0__inst_mult_9_440 ;
wire Xd_0__inst_mult_8_434 ;
wire Xd_0__inst_mult_8_435 ;
wire Xd_0__inst_mult_8_439 ;
wire Xd_0__inst_mult_8_440 ;
wire Xd_0__inst_mult_11_434 ;
wire Xd_0__inst_mult_11_435 ;
wire Xd_0__inst_mult_11_439 ;
wire Xd_0__inst_mult_11_440 ;
wire Xd_0__inst_mult_10_434 ;
wire Xd_0__inst_mult_10_435 ;
wire Xd_0__inst_mult_10_439 ;
wire Xd_0__inst_mult_10_440 ;
wire Xd_0__inst_mult_5_434 ;
wire Xd_0__inst_mult_5_435 ;
wire Xd_0__inst_mult_5_439 ;
wire Xd_0__inst_mult_5_440 ;
wire Xd_0__inst_mult_4_434 ;
wire Xd_0__inst_mult_4_435 ;
wire Xd_0__inst_mult_4_439 ;
wire Xd_0__inst_mult_4_440 ;
wire Xd_0__inst_mult_7_434 ;
wire Xd_0__inst_mult_7_435 ;
wire Xd_0__inst_mult_7_439 ;
wire Xd_0__inst_mult_7_440 ;
wire Xd_0__inst_mult_6_434 ;
wire Xd_0__inst_mult_6_435 ;
wire Xd_0__inst_mult_6_439 ;
wire Xd_0__inst_mult_6_440 ;
wire Xd_0__inst_mult_1_434 ;
wire Xd_0__inst_mult_1_435 ;
wire Xd_0__inst_mult_1_439 ;
wire Xd_0__inst_mult_1_440 ;
wire Xd_0__inst_mult_0_434 ;
wire Xd_0__inst_mult_0_435 ;
wire Xd_0__inst_mult_0_439 ;
wire Xd_0__inst_mult_0_440 ;
wire Xd_0__inst_mult_3_434 ;
wire Xd_0__inst_mult_3_435 ;
wire Xd_0__inst_mult_3_439 ;
wire Xd_0__inst_mult_3_440 ;
wire Xd_0__inst_mult_2_479 ;
wire Xd_0__inst_mult_2_480 ;
wire Xd_0__inst_mult_2_484 ;
wire Xd_0__inst_mult_2_485 ;
wire Xd_0__inst_mult_29_474 ;
wire Xd_0__inst_mult_29_475 ;
wire Xd_0__inst_mult_28_444 ;
wire Xd_0__inst_mult_28_445 ;
wire Xd_0__inst_mult_31_444 ;
wire Xd_0__inst_mult_31_445 ;
wire Xd_0__inst_mult_30_444 ;
wire Xd_0__inst_mult_30_445 ;
wire Xd_0__inst_mult_25_519 ;
wire Xd_0__inst_mult_25_520 ;
wire Xd_0__inst_mult_27_519 ;
wire Xd_0__inst_mult_27_520 ;
wire Xd_0__inst_mult_21_474 ;
wire Xd_0__inst_mult_21_475 ;
wire Xd_0__inst_mult_20_474 ;
wire Xd_0__inst_mult_20_475 ;
wire Xd_0__inst_mult_23_474 ;
wire Xd_0__inst_mult_23_475 ;
wire Xd_0__inst_mult_22_474 ;
wire Xd_0__inst_mult_22_475 ;
wire Xd_0__inst_mult_17_474 ;
wire Xd_0__inst_mult_17_475 ;
wire Xd_0__inst_mult_16_474 ;
wire Xd_0__inst_mult_16_475 ;
wire Xd_0__inst_mult_19_474 ;
wire Xd_0__inst_mult_19_475 ;
wire Xd_0__inst_mult_18_419 ;
wire Xd_0__inst_mult_18_420 ;
wire Xd_0__inst_mult_18_424 ;
wire Xd_0__inst_mult_18_425 ;
wire Xd_0__inst_mult_13_444 ;
wire Xd_0__inst_mult_13_445 ;
wire Xd_0__inst_mult_12_419 ;
wire Xd_0__inst_mult_12_420 ;
wire Xd_0__inst_mult_12_424 ;
wire Xd_0__inst_mult_12_425 ;
wire Xd_0__inst_mult_15_419 ;
wire Xd_0__inst_mult_15_420 ;
wire Xd_0__inst_mult_15_424 ;
wire Xd_0__inst_mult_15_425 ;
wire Xd_0__inst_mult_14_419 ;
wire Xd_0__inst_mult_14_420 ;
wire Xd_0__inst_mult_14_424 ;
wire Xd_0__inst_mult_14_425 ;
wire Xd_0__inst_mult_9_444 ;
wire Xd_0__inst_mult_9_445 ;
wire Xd_0__inst_mult_8_444 ;
wire Xd_0__inst_mult_8_445 ;
wire Xd_0__inst_mult_11_444 ;
wire Xd_0__inst_mult_11_445 ;
wire Xd_0__inst_mult_10_444 ;
wire Xd_0__inst_mult_10_445 ;
wire Xd_0__inst_mult_5_444 ;
wire Xd_0__inst_mult_5_445 ;
wire Xd_0__inst_mult_4_444 ;
wire Xd_0__inst_mult_4_445 ;
wire Xd_0__inst_mult_7_444 ;
wire Xd_0__inst_mult_7_445 ;
wire Xd_0__inst_mult_6_444 ;
wire Xd_0__inst_mult_6_445 ;
wire Xd_0__inst_mult_1_444 ;
wire Xd_0__inst_mult_1_445 ;
wire Xd_0__inst_mult_0_444 ;
wire Xd_0__inst_mult_0_445 ;
wire Xd_0__inst_mult_3_444 ;
wire Xd_0__inst_mult_3_445 ;
wire Xd_0__inst_mult_2_489 ;
wire Xd_0__inst_mult_2_490 ;
wire Xd_0__inst_mult_29_479 ;
wire Xd_0__inst_mult_29_480 ;
wire Xd_0__inst_mult_28_449 ;
wire Xd_0__inst_mult_28_450 ;
wire Xd_0__inst_mult_31_449 ;
wire Xd_0__inst_mult_31_450 ;
wire Xd_0__inst_mult_30_449 ;
wire Xd_0__inst_mult_30_450 ;
wire Xd_0__inst_mult_25_524 ;
wire Xd_0__inst_mult_25_525 ;
wire Xd_0__inst_mult_27_524 ;
wire Xd_0__inst_mult_27_525 ;
wire Xd_0__inst_mult_21_479 ;
wire Xd_0__inst_mult_21_480 ;
wire Xd_0__inst_mult_20_479 ;
wire Xd_0__inst_mult_20_480 ;
wire Xd_0__inst_mult_23_479 ;
wire Xd_0__inst_mult_23_480 ;
wire Xd_0__inst_mult_22_479 ;
wire Xd_0__inst_mult_22_480 ;
wire Xd_0__inst_mult_17_479 ;
wire Xd_0__inst_mult_17_480 ;
wire Xd_0__inst_mult_16_479 ;
wire Xd_0__inst_mult_16_480 ;
wire Xd_0__inst_mult_19_479 ;
wire Xd_0__inst_mult_19_480 ;
wire Xd_0__inst_mult_18_429 ;
wire Xd_0__inst_mult_18_430 ;
wire Xd_0__inst_mult_18_434 ;
wire Xd_0__inst_mult_18_435 ;
wire Xd_0__inst_mult_13_449 ;
wire Xd_0__inst_mult_13_450 ;
wire Xd_0__inst_mult_12_429 ;
wire Xd_0__inst_mult_12_430 ;
wire Xd_0__inst_mult_12_434 ;
wire Xd_0__inst_mult_12_435 ;
wire Xd_0__inst_mult_15_429 ;
wire Xd_0__inst_mult_15_430 ;
wire Xd_0__inst_mult_15_434 ;
wire Xd_0__inst_mult_15_435 ;
wire Xd_0__inst_mult_14_429 ;
wire Xd_0__inst_mult_14_430 ;
wire Xd_0__inst_mult_14_434 ;
wire Xd_0__inst_mult_14_435 ;
wire Xd_0__inst_mult_9_449 ;
wire Xd_0__inst_mult_9_450 ;
wire Xd_0__inst_mult_8_449 ;
wire Xd_0__inst_mult_8_450 ;
wire Xd_0__inst_mult_11_449 ;
wire Xd_0__inst_mult_11_450 ;
wire Xd_0__inst_mult_10_449 ;
wire Xd_0__inst_mult_10_450 ;
wire Xd_0__inst_mult_5_449 ;
wire Xd_0__inst_mult_5_450 ;
wire Xd_0__inst_mult_4_449 ;
wire Xd_0__inst_mult_4_450 ;
wire Xd_0__inst_mult_7_449 ;
wire Xd_0__inst_mult_7_450 ;
wire Xd_0__inst_mult_6_449 ;
wire Xd_0__inst_mult_6_450 ;
wire Xd_0__inst_mult_1_449 ;
wire Xd_0__inst_mult_1_450 ;
wire Xd_0__inst_mult_0_449 ;
wire Xd_0__inst_mult_0_450 ;
wire Xd_0__inst_mult_3_449 ;
wire Xd_0__inst_mult_3_450 ;
wire Xd_0__inst_mult_2_494 ;
wire Xd_0__inst_mult_2_495 ;
wire Xd_0__inst_mult_29_484 ;
wire Xd_0__inst_mult_29_485 ;
wire Xd_0__inst_mult_28_454 ;
wire Xd_0__inst_mult_28_455 ;
wire Xd_0__inst_mult_31_454 ;
wire Xd_0__inst_mult_31_455 ;
wire Xd_0__inst_mult_30_454 ;
wire Xd_0__inst_mult_30_455 ;
wire Xd_0__inst_mult_25_529 ;
wire Xd_0__inst_mult_25_530 ;
wire Xd_0__inst_mult_27_529 ;
wire Xd_0__inst_mult_27_530 ;
wire Xd_0__inst_mult_21_484 ;
wire Xd_0__inst_mult_21_485 ;
wire Xd_0__inst_mult_20_484 ;
wire Xd_0__inst_mult_20_485 ;
wire Xd_0__inst_mult_23_484 ;
wire Xd_0__inst_mult_23_485 ;
wire Xd_0__inst_mult_22_484 ;
wire Xd_0__inst_mult_22_485 ;
wire Xd_0__inst_mult_17_484 ;
wire Xd_0__inst_mult_17_485 ;
wire Xd_0__inst_mult_16_484 ;
wire Xd_0__inst_mult_16_485 ;
wire Xd_0__inst_mult_19_484 ;
wire Xd_0__inst_mult_19_485 ;
wire Xd_0__inst_mult_18_439 ;
wire Xd_0__inst_mult_18_444 ;
wire Xd_0__inst_mult_18_445 ;
wire Xd_0__inst_mult_13_454 ;
wire Xd_0__inst_mult_13_455 ;
wire Xd_0__inst_mult_12_439 ;
wire Xd_0__inst_mult_12_444 ;
wire Xd_0__inst_mult_12_445 ;
wire Xd_0__inst_mult_15_439 ;
wire Xd_0__inst_mult_15_444 ;
wire Xd_0__inst_mult_15_445 ;
wire Xd_0__inst_mult_14_439 ;
wire Xd_0__inst_mult_14_444 ;
wire Xd_0__inst_mult_14_445 ;
wire Xd_0__inst_mult_9_454 ;
wire Xd_0__inst_mult_9_455 ;
wire Xd_0__inst_mult_8_454 ;
wire Xd_0__inst_mult_8_455 ;
wire Xd_0__inst_mult_11_454 ;
wire Xd_0__inst_mult_11_455 ;
wire Xd_0__inst_mult_10_454 ;
wire Xd_0__inst_mult_10_455 ;
wire Xd_0__inst_mult_5_454 ;
wire Xd_0__inst_mult_5_455 ;
wire Xd_0__inst_mult_4_454 ;
wire Xd_0__inst_mult_4_455 ;
wire Xd_0__inst_mult_7_454 ;
wire Xd_0__inst_mult_7_455 ;
wire Xd_0__inst_mult_6_454 ;
wire Xd_0__inst_mult_6_455 ;
wire Xd_0__inst_mult_1_454 ;
wire Xd_0__inst_mult_1_455 ;
wire Xd_0__inst_mult_0_454 ;
wire Xd_0__inst_mult_0_455 ;
wire Xd_0__inst_mult_3_454 ;
wire Xd_0__inst_mult_3_455 ;
wire Xd_0__inst_mult_2_499 ;
wire Xd_0__inst_mult_2_500 ;
wire Xd_0__inst_mult_29_489 ;
wire Xd_0__inst_mult_29_490 ;
wire Xd_0__inst_mult_29_60_sumout ;
wire Xd_0__inst_mult_29_61 ;
wire Xd_0__inst_mult_28_459 ;
wire Xd_0__inst_mult_28_460 ;
wire Xd_0__inst_mult_31_459 ;
wire Xd_0__inst_mult_31_460 ;
wire Xd_0__inst_mult_30_459 ;
wire Xd_0__inst_mult_30_460 ;
wire Xd_0__inst_mult_30_60_sumout ;
wire Xd_0__inst_mult_30_61 ;
wire Xd_0__inst_mult_25_534 ;
wire Xd_0__inst_mult_25_535 ;
wire Xd_0__inst_mult_25_65_sumout ;
wire Xd_0__inst_mult_25_66 ;
wire Xd_0__inst_mult_24_60_sumout ;
wire Xd_0__inst_mult_24_61 ;
wire Xd_0__inst_mult_27_534 ;
wire Xd_0__inst_mult_27_535 ;
wire Xd_0__inst_mult_27_65_sumout ;
wire Xd_0__inst_mult_27_66 ;
wire Xd_0__inst_mult_26_60_sumout ;
wire Xd_0__inst_mult_26_61 ;
wire Xd_0__inst_mult_21_489 ;
wire Xd_0__inst_mult_21_490 ;
wire Xd_0__inst_mult_21_55_sumout ;
wire Xd_0__inst_mult_21_56 ;
wire Xd_0__inst_mult_20_489 ;
wire Xd_0__inst_mult_20_490 ;
wire Xd_0__inst_mult_20_65_sumout ;
wire Xd_0__inst_mult_20_66 ;
wire Xd_0__inst_mult_23_489 ;
wire Xd_0__inst_mult_23_490 ;
wire Xd_0__inst_mult_23_50_sumout ;
wire Xd_0__inst_mult_23_51 ;
wire Xd_0__inst_mult_22_489 ;
wire Xd_0__inst_mult_22_490 ;
wire Xd_0__inst_mult_22_55_sumout ;
wire Xd_0__inst_mult_22_56 ;
wire Xd_0__inst_mult_17_489 ;
wire Xd_0__inst_mult_17_490 ;
wire Xd_0__inst_mult_16_489 ;
wire Xd_0__inst_mult_16_490 ;
wire Xd_0__inst_mult_19_489 ;
wire Xd_0__inst_mult_19_490 ;
wire Xd_0__inst_mult_19_55_sumout ;
wire Xd_0__inst_mult_19_56 ;
wire Xd_0__inst_mult_18_449 ;
wire Xd_0__inst_mult_18_450 ;
wire Xd_0__inst_mult_18_60_sumout ;
wire Xd_0__inst_mult_18_61 ;
wire Xd_0__inst_mult_13_459 ;
wire Xd_0__inst_mult_13_460 ;
wire Xd_0__inst_mult_13_55_sumout ;
wire Xd_0__inst_mult_13_56 ;
wire Xd_0__inst_mult_12_449 ;
wire Xd_0__inst_mult_12_450 ;
wire Xd_0__inst_mult_12_50_sumout ;
wire Xd_0__inst_mult_12_51 ;
wire Xd_0__inst_mult_15_449 ;
wire Xd_0__inst_mult_15_450 ;
wire Xd_0__inst_mult_15_70_sumout ;
wire Xd_0__inst_mult_15_71 ;
wire Xd_0__inst_mult_14_449 ;
wire Xd_0__inst_mult_14_450 ;
wire Xd_0__inst_mult_14_50_sumout ;
wire Xd_0__inst_mult_14_51 ;
wire Xd_0__inst_mult_9_459 ;
wire Xd_0__inst_mult_9_460 ;
wire Xd_0__inst_mult_9_60_sumout ;
wire Xd_0__inst_mult_9_61 ;
wire Xd_0__inst_mult_8_459 ;
wire Xd_0__inst_mult_8_460 ;
wire Xd_0__inst_mult_8_70_sumout ;
wire Xd_0__inst_mult_8_71 ;
wire Xd_0__inst_mult_11_459 ;
wire Xd_0__inst_mult_11_460 ;
wire Xd_0__inst_mult_11_50_sumout ;
wire Xd_0__inst_mult_11_51 ;
wire Xd_0__inst_mult_10_459 ;
wire Xd_0__inst_mult_10_460 ;
wire Xd_0__inst_mult_10_65_sumout ;
wire Xd_0__inst_mult_10_66 ;
wire Xd_0__inst_mult_5_459 ;
wire Xd_0__inst_mult_5_460 ;
wire Xd_0__inst_mult_4_459 ;
wire Xd_0__inst_mult_4_460 ;
wire Xd_0__inst_mult_4_50_sumout ;
wire Xd_0__inst_mult_4_51 ;
wire Xd_0__inst_mult_7_459 ;
wire Xd_0__inst_mult_7_460 ;
wire Xd_0__inst_mult_7_65_sumout ;
wire Xd_0__inst_mult_7_66 ;
wire Xd_0__inst_mult_6_459 ;
wire Xd_0__inst_mult_6_460 ;
wire Xd_0__inst_mult_6_65_sumout ;
wire Xd_0__inst_mult_6_66 ;
wire Xd_0__inst_mult_1_459 ;
wire Xd_0__inst_mult_1_460 ;
wire Xd_0__inst_mult_1_50_sumout ;
wire Xd_0__inst_mult_1_51 ;
wire Xd_0__inst_mult_0_459 ;
wire Xd_0__inst_mult_0_460 ;
wire Xd_0__inst_mult_0_60_sumout ;
wire Xd_0__inst_mult_0_61 ;
wire Xd_0__inst_mult_3_459 ;
wire Xd_0__inst_mult_3_460 ;
wire Xd_0__inst_mult_3_70_sumout ;
wire Xd_0__inst_mult_3_71 ;
wire Xd_0__inst_mult_2_504 ;
wire Xd_0__inst_mult_2_505 ;
wire Xd_0__inst_mult_2_60_sumout ;
wire Xd_0__inst_mult_2_61 ;
wire Xd_0__inst_mult_29_494 ;
wire Xd_0__inst_mult_29_495 ;
wire Xd_0__inst_mult_29_65_sumout ;
wire Xd_0__inst_mult_29_66 ;
wire Xd_0__inst_mult_28_464 ;
wire Xd_0__inst_mult_28_465 ;
wire Xd_0__inst_mult_28_65_sumout ;
wire Xd_0__inst_mult_28_66 ;
wire Xd_0__inst_mult_31_464 ;
wire Xd_0__inst_mult_31_465 ;
wire Xd_0__inst_mult_31_55_sumout ;
wire Xd_0__inst_mult_31_56 ;
wire Xd_0__inst_mult_30_464 ;
wire Xd_0__inst_mult_30_465 ;
wire Xd_0__inst_mult_30_65_sumout ;
wire Xd_0__inst_mult_30_66 ;
wire Xd_0__inst_mult_25_539 ;
wire Xd_0__inst_mult_25_540 ;
wire Xd_0__inst_mult_25_70_sumout ;
wire Xd_0__inst_mult_25_71 ;
wire Xd_0__inst_mult_24_65_sumout ;
wire Xd_0__inst_mult_24_66 ;
wire Xd_0__inst_mult_27_539 ;
wire Xd_0__inst_mult_27_540 ;
wire Xd_0__inst_mult_27_70_sumout ;
wire Xd_0__inst_mult_27_71 ;
wire Xd_0__inst_mult_26_65_sumout ;
wire Xd_0__inst_mult_26_66 ;
wire Xd_0__inst_mult_21_494 ;
wire Xd_0__inst_mult_21_495 ;
wire Xd_0__inst_mult_21_60_sumout ;
wire Xd_0__inst_mult_21_61 ;
wire Xd_0__inst_mult_20_494 ;
wire Xd_0__inst_mult_20_495 ;
wire Xd_0__inst_mult_20_70_sumout ;
wire Xd_0__inst_mult_20_71 ;
wire Xd_0__inst_mult_23_494 ;
wire Xd_0__inst_mult_23_495 ;
wire Xd_0__inst_mult_23_55_sumout ;
wire Xd_0__inst_mult_23_56 ;
wire Xd_0__inst_mult_22_494 ;
wire Xd_0__inst_mult_22_495 ;
wire Xd_0__inst_mult_22_60_sumout ;
wire Xd_0__inst_mult_22_61 ;
wire Xd_0__inst_mult_17_494 ;
wire Xd_0__inst_mult_17_495 ;
wire Xd_0__inst_mult_17_65_sumout ;
wire Xd_0__inst_mult_17_66 ;
wire Xd_0__inst_mult_16_494 ;
wire Xd_0__inst_mult_16_495 ;
wire Xd_0__inst_mult_16_55_sumout ;
wire Xd_0__inst_mult_16_56 ;
wire Xd_0__inst_mult_19_494 ;
wire Xd_0__inst_mult_19_495 ;
wire Xd_0__inst_mult_19_60_sumout ;
wire Xd_0__inst_mult_19_61 ;
wire Xd_0__inst_mult_18_454 ;
wire Xd_0__inst_mult_18_455 ;
wire Xd_0__inst_mult_18_65_sumout ;
wire Xd_0__inst_mult_18_66 ;
wire Xd_0__inst_mult_13_464 ;
wire Xd_0__inst_mult_13_465 ;
wire Xd_0__inst_mult_13_60_sumout ;
wire Xd_0__inst_mult_13_61 ;
wire Xd_0__inst_mult_12_454 ;
wire Xd_0__inst_mult_12_455 ;
wire Xd_0__inst_mult_12_55_sumout ;
wire Xd_0__inst_mult_12_56 ;
wire Xd_0__inst_mult_15_454 ;
wire Xd_0__inst_mult_15_455 ;
wire Xd_0__inst_mult_15_75_sumout ;
wire Xd_0__inst_mult_15_76 ;
wire Xd_0__inst_mult_14_454 ;
wire Xd_0__inst_mult_14_455 ;
wire Xd_0__inst_mult_14_55_sumout ;
wire Xd_0__inst_mult_14_56 ;
wire Xd_0__inst_mult_9_464 ;
wire Xd_0__inst_mult_9_465 ;
wire Xd_0__inst_mult_9_65_sumout ;
wire Xd_0__inst_mult_9_66 ;
wire Xd_0__inst_mult_8_464 ;
wire Xd_0__inst_mult_8_465 ;
wire Xd_0__inst_mult_8_75_sumout ;
wire Xd_0__inst_mult_8_76 ;
wire Xd_0__inst_mult_11_464 ;
wire Xd_0__inst_mult_11_465 ;
wire Xd_0__inst_mult_11_55_sumout ;
wire Xd_0__inst_mult_11_56 ;
wire Xd_0__inst_mult_10_464 ;
wire Xd_0__inst_mult_10_465 ;
wire Xd_0__inst_mult_10_70_sumout ;
wire Xd_0__inst_mult_10_71 ;
wire Xd_0__inst_mult_5_464 ;
wire Xd_0__inst_mult_5_465 ;
wire Xd_0__inst_mult_4_464 ;
wire Xd_0__inst_mult_4_465 ;
wire Xd_0__inst_mult_4_55_sumout ;
wire Xd_0__inst_mult_4_56 ;
wire Xd_0__inst_mult_7_464 ;
wire Xd_0__inst_mult_7_465 ;
wire Xd_0__inst_mult_7_70_sumout ;
wire Xd_0__inst_mult_7_71 ;
wire Xd_0__inst_mult_6_464 ;
wire Xd_0__inst_mult_6_465 ;
wire Xd_0__inst_mult_6_70_sumout ;
wire Xd_0__inst_mult_6_71 ;
wire Xd_0__inst_mult_1_464 ;
wire Xd_0__inst_mult_1_465 ;
wire Xd_0__inst_mult_1_55_sumout ;
wire Xd_0__inst_mult_1_56 ;
wire Xd_0__inst_mult_0_464 ;
wire Xd_0__inst_mult_0_465 ;
wire Xd_0__inst_mult_0_65_sumout ;
wire Xd_0__inst_mult_0_66 ;
wire Xd_0__inst_mult_3_464 ;
wire Xd_0__inst_mult_3_465 ;
wire Xd_0__inst_mult_3_75_sumout ;
wire Xd_0__inst_mult_3_76 ;
wire Xd_0__inst_mult_2_509 ;
wire Xd_0__inst_mult_2_510 ;
wire Xd_0__inst_mult_2_65_sumout ;
wire Xd_0__inst_mult_2_66 ;
wire Xd_0__inst_mult_29_499 ;
wire Xd_0__inst_mult_29_500 ;
wire Xd_0__inst_mult_29_70_sumout ;
wire Xd_0__inst_mult_29_71 ;
wire Xd_0__inst_mult_28_469 ;
wire Xd_0__inst_mult_28_470 ;
wire Xd_0__inst_mult_28_70_sumout ;
wire Xd_0__inst_mult_28_71 ;
wire Xd_0__inst_mult_31_469 ;
wire Xd_0__inst_mult_31_470 ;
wire Xd_0__inst_mult_31_60_sumout ;
wire Xd_0__inst_mult_31_61 ;
wire Xd_0__inst_mult_30_469 ;
wire Xd_0__inst_mult_30_470 ;
wire Xd_0__inst_mult_30_70_sumout ;
wire Xd_0__inst_mult_30_71 ;
wire Xd_0__inst_mult_25_544 ;
wire Xd_0__inst_mult_25_545 ;
wire Xd_0__inst_mult_25_75_sumout ;
wire Xd_0__inst_mult_25_76 ;
wire Xd_0__inst_mult_24_70_sumout ;
wire Xd_0__inst_mult_24_71 ;
wire Xd_0__inst_mult_27_544 ;
wire Xd_0__inst_mult_27_545 ;
wire Xd_0__inst_mult_27_75_sumout ;
wire Xd_0__inst_mult_27_76 ;
wire Xd_0__inst_mult_26_70_sumout ;
wire Xd_0__inst_mult_26_71 ;
wire Xd_0__inst_mult_21_499 ;
wire Xd_0__inst_mult_21_500 ;
wire Xd_0__inst_mult_21_65_sumout ;
wire Xd_0__inst_mult_21_66 ;
wire Xd_0__inst_mult_20_499 ;
wire Xd_0__inst_mult_20_500 ;
wire Xd_0__inst_mult_20_75_sumout ;
wire Xd_0__inst_mult_20_76 ;
wire Xd_0__inst_mult_23_499 ;
wire Xd_0__inst_mult_23_500 ;
wire Xd_0__inst_mult_23_60_sumout ;
wire Xd_0__inst_mult_23_61 ;
wire Xd_0__inst_mult_22_499 ;
wire Xd_0__inst_mult_22_500 ;
wire Xd_0__inst_mult_22_65_sumout ;
wire Xd_0__inst_mult_22_66 ;
wire Xd_0__inst_mult_17_499 ;
wire Xd_0__inst_mult_17_500 ;
wire Xd_0__inst_mult_17_70_sumout ;
wire Xd_0__inst_mult_17_71 ;
wire Xd_0__inst_mult_16_499 ;
wire Xd_0__inst_mult_16_500 ;
wire Xd_0__inst_mult_16_60_sumout ;
wire Xd_0__inst_mult_16_61 ;
wire Xd_0__inst_mult_19_499 ;
wire Xd_0__inst_mult_19_500 ;
wire Xd_0__inst_mult_19_65_sumout ;
wire Xd_0__inst_mult_19_66 ;
wire Xd_0__inst_mult_18_459 ;
wire Xd_0__inst_mult_18_460 ;
wire Xd_0__inst_mult_13_469 ;
wire Xd_0__inst_mult_13_470 ;
wire Xd_0__inst_mult_13_65_sumout ;
wire Xd_0__inst_mult_13_66 ;
wire Xd_0__inst_mult_12_459 ;
wire Xd_0__inst_mult_12_460 ;
wire Xd_0__inst_mult_12_60_sumout ;
wire Xd_0__inst_mult_12_61 ;
wire Xd_0__inst_mult_15_459 ;
wire Xd_0__inst_mult_15_460 ;
wire Xd_0__inst_mult_15_80_sumout ;
wire Xd_0__inst_mult_15_81 ;
wire Xd_0__inst_mult_14_459 ;
wire Xd_0__inst_mult_14_460 ;
wire Xd_0__inst_mult_14_60_sumout ;
wire Xd_0__inst_mult_14_61 ;
wire Xd_0__inst_mult_9_469 ;
wire Xd_0__inst_mult_9_470 ;
wire Xd_0__inst_mult_9_70_sumout ;
wire Xd_0__inst_mult_9_71 ;
wire Xd_0__inst_mult_8_469 ;
wire Xd_0__inst_mult_8_470 ;
wire Xd_0__inst_mult_8_80_sumout ;
wire Xd_0__inst_mult_8_81 ;
wire Xd_0__inst_mult_11_469 ;
wire Xd_0__inst_mult_11_470 ;
wire Xd_0__inst_mult_11_60_sumout ;
wire Xd_0__inst_mult_11_61 ;
wire Xd_0__inst_mult_10_469 ;
wire Xd_0__inst_mult_10_470 ;
wire Xd_0__inst_mult_10_75_sumout ;
wire Xd_0__inst_mult_10_76 ;
wire Xd_0__inst_mult_5_469 ;
wire Xd_0__inst_mult_5_470 ;
wire Xd_0__inst_mult_5_80_sumout ;
wire Xd_0__inst_mult_5_81 ;
wire Xd_0__inst_mult_4_469 ;
wire Xd_0__inst_mult_4_470 ;
wire Xd_0__inst_mult_4_60_sumout ;
wire Xd_0__inst_mult_4_61 ;
wire Xd_0__inst_mult_7_469 ;
wire Xd_0__inst_mult_7_470 ;
wire Xd_0__inst_mult_7_75_sumout ;
wire Xd_0__inst_mult_7_76 ;
wire Xd_0__inst_mult_6_469 ;
wire Xd_0__inst_mult_6_470 ;
wire Xd_0__inst_mult_6_75_sumout ;
wire Xd_0__inst_mult_6_76 ;
wire Xd_0__inst_mult_1_469 ;
wire Xd_0__inst_mult_1_470 ;
wire Xd_0__inst_mult_1_60_sumout ;
wire Xd_0__inst_mult_1_61 ;
wire Xd_0__inst_mult_0_469 ;
wire Xd_0__inst_mult_0_470 ;
wire Xd_0__inst_mult_0_70_sumout ;
wire Xd_0__inst_mult_0_71 ;
wire Xd_0__inst_mult_3_469 ;
wire Xd_0__inst_mult_3_470 ;
wire Xd_0__inst_mult_3_80_sumout ;
wire Xd_0__inst_mult_3_81 ;
wire Xd_0__inst_mult_2_514 ;
wire Xd_0__inst_mult_2_515 ;
wire Xd_0__inst_mult_2_70_sumout ;
wire Xd_0__inst_mult_2_71 ;
wire Xd_0__inst_mult_29_504 ;
wire Xd_0__inst_mult_29_505 ;
wire Xd_0__inst_mult_29_75_sumout ;
wire Xd_0__inst_mult_29_76 ;
wire Xd_0__inst_mult_28_474 ;
wire Xd_0__inst_mult_28_475 ;
wire Xd_0__inst_mult_28_75_sumout ;
wire Xd_0__inst_mult_28_76 ;
wire Xd_0__inst_mult_31_474 ;
wire Xd_0__inst_mult_31_475 ;
wire Xd_0__inst_mult_31_65_sumout ;
wire Xd_0__inst_mult_31_66 ;
wire Xd_0__inst_mult_30_474 ;
wire Xd_0__inst_mult_30_475 ;
wire Xd_0__inst_mult_30_75_sumout ;
wire Xd_0__inst_mult_30_76 ;
wire Xd_0__inst_mult_25_549 ;
wire Xd_0__inst_mult_25_550 ;
wire Xd_0__inst_mult_25_80_sumout ;
wire Xd_0__inst_mult_25_81 ;
wire Xd_0__inst_mult_24_75_sumout ;
wire Xd_0__inst_mult_24_76 ;
wire Xd_0__inst_mult_27_549 ;
wire Xd_0__inst_mult_27_550 ;
wire Xd_0__inst_mult_27_80_sumout ;
wire Xd_0__inst_mult_27_81 ;
wire Xd_0__inst_mult_26_75_sumout ;
wire Xd_0__inst_mult_26_76 ;
wire Xd_0__inst_mult_21_504 ;
wire Xd_0__inst_mult_21_505 ;
wire Xd_0__inst_mult_21_70_sumout ;
wire Xd_0__inst_mult_21_71 ;
wire Xd_0__inst_mult_20_504 ;
wire Xd_0__inst_mult_20_505 ;
wire Xd_0__inst_mult_20_80_sumout ;
wire Xd_0__inst_mult_20_81 ;
wire Xd_0__inst_mult_23_504 ;
wire Xd_0__inst_mult_23_505 ;
wire Xd_0__inst_mult_23_65_sumout ;
wire Xd_0__inst_mult_23_66 ;
wire Xd_0__inst_mult_22_504 ;
wire Xd_0__inst_mult_22_505 ;
wire Xd_0__inst_mult_22_70_sumout ;
wire Xd_0__inst_mult_22_71 ;
wire Xd_0__inst_mult_17_504 ;
wire Xd_0__inst_mult_17_505 ;
wire Xd_0__inst_mult_17_75_sumout ;
wire Xd_0__inst_mult_17_76 ;
wire Xd_0__inst_mult_16_504 ;
wire Xd_0__inst_mult_16_505 ;
wire Xd_0__inst_mult_16_65_sumout ;
wire Xd_0__inst_mult_16_66 ;
wire Xd_0__inst_mult_19_504 ;
wire Xd_0__inst_mult_19_505 ;
wire Xd_0__inst_mult_19_70_sumout ;
wire Xd_0__inst_mult_19_71 ;
wire Xd_0__inst_mult_18_464 ;
wire Xd_0__inst_mult_18_465 ;
wire Xd_0__inst_mult_18_70_sumout ;
wire Xd_0__inst_mult_18_71 ;
wire Xd_0__inst_mult_13_474 ;
wire Xd_0__inst_mult_13_475 ;
wire Xd_0__inst_mult_13_70_sumout ;
wire Xd_0__inst_mult_13_71 ;
wire Xd_0__inst_mult_12_464 ;
wire Xd_0__inst_mult_12_465 ;
wire Xd_0__inst_mult_15_464 ;
wire Xd_0__inst_mult_15_465 ;
wire Xd_0__inst_mult_14_464 ;
wire Xd_0__inst_mult_14_465 ;
wire Xd_0__inst_mult_14_65_sumout ;
wire Xd_0__inst_mult_14_66 ;
wire Xd_0__inst_mult_9_474 ;
wire Xd_0__inst_mult_9_475 ;
wire Xd_0__inst_mult_8_474 ;
wire Xd_0__inst_mult_8_475 ;
wire Xd_0__inst_mult_11_474 ;
wire Xd_0__inst_mult_11_475 ;
wire Xd_0__inst_mult_11_65_sumout ;
wire Xd_0__inst_mult_11_66 ;
wire Xd_0__inst_mult_10_474 ;
wire Xd_0__inst_mult_10_475 ;
wire Xd_0__inst_mult_5_474 ;
wire Xd_0__inst_mult_5_475 ;
wire Xd_0__inst_mult_4_474 ;
wire Xd_0__inst_mult_4_475 ;
wire Xd_0__inst_mult_4_65_sumout ;
wire Xd_0__inst_mult_4_66 ;
wire Xd_0__inst_mult_7_474 ;
wire Xd_0__inst_mult_7_475 ;
wire Xd_0__inst_mult_6_474 ;
wire Xd_0__inst_mult_6_475 ;
wire Xd_0__inst_mult_1_474 ;
wire Xd_0__inst_mult_1_475 ;
wire Xd_0__inst_mult_1_65_sumout ;
wire Xd_0__inst_mult_1_66 ;
wire Xd_0__inst_mult_0_474 ;
wire Xd_0__inst_mult_0_475 ;
wire Xd_0__inst_mult_3_474 ;
wire Xd_0__inst_mult_3_475 ;
wire Xd_0__inst_mult_2_519 ;
wire Xd_0__inst_mult_2_520 ;
wire Xd_0__inst_mult_2_75_sumout ;
wire Xd_0__inst_mult_2_76 ;
wire Xd_0__inst_mult_29_509 ;
wire Xd_0__inst_mult_28_479 ;
wire Xd_0__inst_mult_31_479 ;
wire Xd_0__inst_mult_31_70_sumout ;
wire Xd_0__inst_mult_31_71 ;
wire Xd_0__inst_mult_30_479 ;
wire Xd_0__inst_mult_25_554 ;
wire Xd_0__inst_mult_24_80_sumout ;
wire Xd_0__inst_mult_24_81 ;
wire Xd_0__inst_mult_27_554 ;
wire Xd_0__inst_mult_26_80_sumout ;
wire Xd_0__inst_mult_26_81 ;
wire Xd_0__inst_mult_21_509 ;
wire Xd_0__inst_mult_20_509 ;
wire Xd_0__inst_mult_23_509 ;
wire Xd_0__inst_mult_23_70_sumout ;
wire Xd_0__inst_mult_23_71 ;
wire Xd_0__inst_mult_22_509 ;
wire Xd_0__inst_mult_17_509 ;
wire Xd_0__inst_mult_16_509 ;
wire Xd_0__inst_mult_16_70_sumout ;
wire Xd_0__inst_mult_16_71 ;
wire Xd_0__inst_mult_19_509 ;
wire Xd_0__inst_mult_18_469 ;
wire Xd_0__inst_mult_13_479 ;
wire Xd_0__inst_mult_12_469 ;
wire Xd_0__inst_mult_12_65_sumout ;
wire Xd_0__inst_mult_12_66 ;
wire Xd_0__inst_mult_15_469 ;
wire Xd_0__inst_mult_14_469 ;
wire Xd_0__inst_mult_14_70_sumout ;
wire Xd_0__inst_mult_14_71 ;
wire Xd_0__inst_mult_9_479 ;
wire Xd_0__inst_mult_8_479 ;
wire Xd_0__inst_mult_11_479 ;
wire Xd_0__inst_mult_11_70_sumout ;
wire Xd_0__inst_mult_11_71 ;
wire Xd_0__inst_mult_10_479 ;
wire Xd_0__inst_mult_5_479 ;
wire Xd_0__inst_mult_4_479 ;
wire Xd_0__inst_mult_4_70_sumout ;
wire Xd_0__inst_mult_4_71 ;
wire Xd_0__inst_mult_7_479 ;
wire Xd_0__inst_mult_6_479 ;
wire Xd_0__inst_mult_1_479 ;
wire Xd_0__inst_mult_1_70_sumout ;
wire Xd_0__inst_mult_1_71 ;
wire Xd_0__inst_mult_0_479 ;
wire Xd_0__inst_mult_0_75_sumout ;
wire Xd_0__inst_mult_0_76 ;
wire Xd_0__inst_mult_3_479 ;
wire Xd_0__inst_mult_2_524 ;
wire Xd_0__inst_mult_9_484 ;
wire Xd_0__inst_mult_9_489 ;
wire Xd_0__inst_mult_9_490 ;
wire Xd_0__inst_mult_9_494 ;
wire Xd_0__inst_mult_8_484 ;
wire Xd_0__inst_mult_8_489 ;
wire Xd_0__inst_mult_8_490 ;
wire Xd_0__inst_mult_8_494 ;
wire Xd_0__inst_mult_21_514 ;
wire Xd_0__inst_mult_21_515 ;
wire Xd_0__inst_mult_21_519 ;
wire Xd_0__inst_mult_21_520 ;
wire Xd_0__inst_mult_21_524 ;
wire Xd_0__inst_mult_21_525 ;
wire Xd_0__inst_mult_11_484 ;
wire Xd_0__inst_mult_11_489 ;
wire Xd_0__inst_mult_11_490 ;
wire Xd_0__inst_mult_11_494 ;
wire Xd_0__inst_mult_10_484 ;
wire Xd_0__inst_mult_10_489 ;
wire Xd_0__inst_mult_10_490 ;
wire Xd_0__inst_mult_10_494 ;
wire Xd_0__inst_mult_20_514 ;
wire Xd_0__inst_mult_20_515 ;
wire Xd_0__inst_mult_20_519 ;
wire Xd_0__inst_mult_20_520 ;
wire Xd_0__inst_mult_20_524 ;
wire Xd_0__inst_mult_20_525 ;
wire Xd_0__inst_mult_25_559 ;
wire Xd_0__inst_mult_25_560 ;
wire Xd_0__inst_mult_25_564 ;
wire Xd_0__inst_mult_25_565 ;
wire Xd_0__inst_mult_25_569 ;
wire Xd_0__inst_mult_25_570 ;
wire Xd_0__inst_mult_3_484 ;
wire Xd_0__inst_mult_3_489 ;
wire Xd_0__inst_mult_3_490 ;
wire Xd_0__inst_mult_12_70_sumout ;
wire Xd_0__inst_mult_12_71 ;
wire Xd_0__inst_mult_3_494 ;
wire Xd_0__inst_mult_0_484 ;
wire Xd_0__inst_mult_0_489 ;
wire Xd_0__inst_mult_0_490 ;
wire Xd_0__inst_mult_0_494 ;
wire Xd_0__inst_mult_23_514 ;
wire Xd_0__inst_mult_23_515 ;
wire Xd_0__inst_mult_23_519 ;
wire Xd_0__inst_mult_23_520 ;
wire Xd_0__inst_mult_23_524 ;
wire Xd_0__inst_mult_23_525 ;
wire Xd_0__inst_mult_6_484 ;
wire Xd_0__inst_mult_6_489 ;
wire Xd_0__inst_mult_6_490 ;
wire Xd_0__inst_mult_6_494 ;
wire Xd_0__inst_mult_1_484 ;
wire Xd_0__inst_mult_1_489 ;
wire Xd_0__inst_mult_1_490 ;
wire Xd_0__inst_mult_1_494 ;
wire Xd_0__inst_mult_22_514 ;
wire Xd_0__inst_mult_22_515 ;
wire Xd_0__inst_mult_22_519 ;
wire Xd_0__inst_mult_22_520 ;
wire Xd_0__inst_mult_22_524 ;
wire Xd_0__inst_mult_22_525 ;
wire Xd_0__inst_mult_24_699 ;
wire Xd_0__inst_mult_24_700 ;
wire Xd_0__inst_mult_24_704 ;
wire Xd_0__inst_mult_24_705 ;
wire Xd_0__inst_mult_24_709 ;
wire Xd_0__inst_mult_24_710 ;
wire Xd_0__inst_mult_26_699 ;
wire Xd_0__inst_mult_26_700 ;
wire Xd_0__inst_mult_26_704 ;
wire Xd_0__inst_mult_26_705 ;
wire Xd_0__inst_mult_26_709 ;
wire Xd_0__inst_mult_26_710 ;
wire Xd_0__inst_mult_7_484 ;
wire Xd_0__inst_mult_7_489 ;
wire Xd_0__inst_mult_7_490 ;
wire Xd_0__inst_mult_7_494 ;
wire Xd_0__inst_mult_4_484 ;
wire Xd_0__inst_mult_4_489 ;
wire Xd_0__inst_mult_4_490 ;
wire Xd_0__inst_mult_4_494 ;
wire Xd_0__inst_mult_19_514 ;
wire Xd_0__inst_mult_19_515 ;
wire Xd_0__inst_mult_19_519 ;
wire Xd_0__inst_mult_19_520 ;
wire Xd_0__inst_mult_19_524 ;
wire Xd_0__inst_mult_19_525 ;
wire Xd_0__inst_mult_30_484 ;
wire Xd_0__inst_mult_30_489 ;
wire Xd_0__inst_mult_30_490 ;
wire Xd_0__inst_mult_30_494 ;
wire Xd_0__inst_mult_5_484 ;
wire Xd_0__inst_mult_5_489 ;
wire Xd_0__inst_mult_5_490 ;
wire Xd_0__inst_mult_5_494 ;
wire Xd_0__inst_mult_17_514 ;
wire Xd_0__inst_mult_17_515 ;
wire Xd_0__inst_mult_17_519 ;
wire Xd_0__inst_mult_17_520 ;
wire Xd_0__inst_mult_17_524 ;
wire Xd_0__inst_mult_17_525 ;
wire Xd_0__inst_mult_27_559 ;
wire Xd_0__inst_mult_27_560 ;
wire Xd_0__inst_mult_27_564 ;
wire Xd_0__inst_mult_27_565 ;
wire Xd_0__inst_mult_27_569 ;
wire Xd_0__inst_mult_27_570 ;
wire Xd_0__inst_mult_13_484 ;
wire Xd_0__inst_mult_13_489 ;
wire Xd_0__inst_mult_13_490 ;
wire Xd_0__inst_mult_13_494 ;
wire Xd_0__inst_mult_2_529 ;
wire Xd_0__inst_mult_2_534 ;
wire Xd_0__inst_mult_2_535 ;
wire Xd_0__inst_mult_2_539 ;
wire Xd_0__inst_mult_16_514 ;
wire Xd_0__inst_mult_16_515 ;
wire Xd_0__inst_mult_16_519 ;
wire Xd_0__inst_mult_16_520 ;
wire Xd_0__inst_mult_16_524 ;
wire Xd_0__inst_mult_16_525 ;
wire Xd_0__inst_mult_28_484 ;
wire Xd_0__inst_mult_28_489 ;
wire Xd_0__inst_mult_28_490 ;
wire Xd_0__inst_mult_28_494 ;
wire Xd_0__inst_mult_31_484 ;
wire Xd_0__inst_mult_31_489 ;
wire Xd_0__inst_mult_31_490 ;
wire Xd_0__inst_mult_31_494 ;
wire Xd_0__inst_mult_29_514 ;
wire Xd_0__inst_mult_29_515 ;
wire Xd_0__inst_mult_29_519 ;
wire Xd_0__inst_mult_29_520 ;
wire Xd_0__inst_mult_29_524 ;
wire Xd_0__inst_mult_29_525 ;
wire Xd_0__inst_mult_26_714 ;
wire Xd_0__inst_mult_26_715 ;
wire Xd_0__inst_mult_26_719 ;
wire Xd_0__inst_mult_26_720 ;
wire Xd_0__inst_mult_26_724 ;
wire Xd_0__inst_mult_26_725 ;
wire Xd_0__inst_mult_24_714 ;
wire Xd_0__inst_mult_24_715 ;
wire Xd_0__inst_mult_24_719 ;
wire Xd_0__inst_mult_24_720 ;
wire Xd_0__inst_mult_24_724 ;
wire Xd_0__inst_mult_24_725 ;
wire Xd_0__inst_mult_22_75_sumout ;
wire Xd_0__inst_mult_22_76 ;
wire Xd_0__inst_mult_12_75_sumout ;
wire Xd_0__inst_mult_12_76 ;
wire Xd_0__inst_mult_10_80_sumout ;
wire Xd_0__inst_mult_10_81 ;
wire Xd_0__inst_mult_0_80_sumout ;
wire Xd_0__inst_mult_0_81 ;
wire Xd_0__inst_mult_29_529 ;
wire Xd_0__inst_mult_29_530 ;
wire Xd_0__inst_mult_29_534 ;
wire Xd_0__inst_mult_29_535 ;
wire Xd_0__inst_mult_28_499 ;
wire Xd_0__inst_mult_28_500 ;
wire Xd_0__inst_mult_28_504 ;
wire Xd_0__inst_mult_28_505 ;
wire Xd_0__inst_mult_31_499 ;
wire Xd_0__inst_mult_31_500 ;
wire Xd_0__inst_mult_31_504 ;
wire Xd_0__inst_mult_31_505 ;
wire Xd_0__inst_mult_30_499 ;
wire Xd_0__inst_mult_30_500 ;
wire Xd_0__inst_mult_30_504 ;
wire Xd_0__inst_mult_30_505 ;
wire Xd_0__inst_mult_21_75_sumout ;
wire Xd_0__inst_mult_21_76 ;
wire Xd_0__inst_mult_25_574 ;
wire Xd_0__inst_mult_25_575 ;
wire Xd_0__inst_mult_25_579 ;
wire Xd_0__inst_mult_25_580 ;
wire Xd_0__inst_mult_24_729 ;
wire Xd_0__inst_mult_24_730 ;
wire Xd_0__inst_mult_24_734 ;
wire Xd_0__inst_mult_24_735 ;
wire Xd_0__inst_mult_31_75_sumout ;
wire Xd_0__inst_mult_31_76 ;
wire Xd_0__inst_mult_27_574 ;
wire Xd_0__inst_mult_27_575 ;
wire Xd_0__inst_mult_27_579 ;
wire Xd_0__inst_mult_27_580 ;
wire Xd_0__inst_mult_23_75_sumout ;
wire Xd_0__inst_mult_23_76 ;
wire Xd_0__inst_mult_26_729 ;
wire Xd_0__inst_mult_26_730 ;
wire Xd_0__inst_mult_26_734 ;
wire Xd_0__inst_mult_26_735 ;
wire Xd_0__inst_mult_1_75_sumout ;
wire Xd_0__inst_mult_1_76 ;
wire Xd_0__inst_mult_21_529 ;
wire Xd_0__inst_mult_21_530 ;
wire Xd_0__inst_mult_21_534 ;
wire Xd_0__inst_mult_21_535 ;
wire Xd_0__inst_mult_4_75_sumout ;
wire Xd_0__inst_mult_4_76 ;
wire Xd_0__inst_mult_20_529 ;
wire Xd_0__inst_mult_20_530 ;
wire Xd_0__inst_mult_20_534 ;
wire Xd_0__inst_mult_20_535 ;
wire Xd_0__inst_mult_23_529 ;
wire Xd_0__inst_mult_23_530 ;
wire Xd_0__inst_mult_23_534 ;
wire Xd_0__inst_mult_23_535 ;
wire Xd_0__inst_mult_2_80_sumout ;
wire Xd_0__inst_mult_2_81 ;
wire Xd_0__inst_mult_22_529 ;
wire Xd_0__inst_mult_22_530 ;
wire Xd_0__inst_mult_22_534 ;
wire Xd_0__inst_mult_22_535 ;
wire Xd_0__inst_mult_17_529 ;
wire Xd_0__inst_mult_17_530 ;
wire Xd_0__inst_mult_17_534 ;
wire Xd_0__inst_mult_17_535 ;
wire Xd_0__inst_mult_11_75_sumout ;
wire Xd_0__inst_mult_11_76 ;
wire Xd_0__inst_mult_16_529 ;
wire Xd_0__inst_mult_16_530 ;
wire Xd_0__inst_mult_16_534 ;
wire Xd_0__inst_mult_16_535 ;
wire Xd_0__inst_mult_19_529 ;
wire Xd_0__inst_mult_19_530 ;
wire Xd_0__inst_mult_19_534 ;
wire Xd_0__inst_mult_19_535 ;
wire Xd_0__inst_mult_18_474 ;
wire Xd_0__inst_mult_18_475 ;
wire Xd_0__inst_mult_18_479 ;
wire Xd_0__inst_mult_18_480 ;
wire Xd_0__inst_mult_13_499 ;
wire Xd_0__inst_mult_13_500 ;
wire Xd_0__inst_mult_13_504 ;
wire Xd_0__inst_mult_13_505 ;
wire Xd_0__inst_mult_12_474 ;
wire Xd_0__inst_mult_12_475 ;
wire Xd_0__inst_mult_12_479 ;
wire Xd_0__inst_mult_12_480 ;
wire Xd_0__inst_mult_15_474 ;
wire Xd_0__inst_mult_15_475 ;
wire Xd_0__inst_mult_15_479 ;
wire Xd_0__inst_mult_15_480 ;
wire Xd_0__inst_mult_14_474 ;
wire Xd_0__inst_mult_14_475 ;
wire Xd_0__inst_mult_14_479 ;
wire Xd_0__inst_mult_14_480 ;
wire Xd_0__inst_mult_9_499 ;
wire Xd_0__inst_mult_9_500 ;
wire Xd_0__inst_mult_9_504 ;
wire Xd_0__inst_mult_9_505 ;
wire Xd_0__inst_mult_8_499 ;
wire Xd_0__inst_mult_8_500 ;
wire Xd_0__inst_mult_8_504 ;
wire Xd_0__inst_mult_8_505 ;
wire Xd_0__inst_mult_11_499 ;
wire Xd_0__inst_mult_11_500 ;
wire Xd_0__inst_mult_11_504 ;
wire Xd_0__inst_mult_11_505 ;
wire Xd_0__inst_mult_10_499 ;
wire Xd_0__inst_mult_10_500 ;
wire Xd_0__inst_mult_10_504 ;
wire Xd_0__inst_mult_10_505 ;
wire Xd_0__inst_mult_5_499 ;
wire Xd_0__inst_mult_5_500 ;
wire Xd_0__inst_mult_5_504 ;
wire Xd_0__inst_mult_5_505 ;
wire Xd_0__inst_mult_4_499 ;
wire Xd_0__inst_mult_4_500 ;
wire Xd_0__inst_mult_4_504 ;
wire Xd_0__inst_mult_4_505 ;
wire Xd_0__inst_mult_7_499 ;
wire Xd_0__inst_mult_7_500 ;
wire Xd_0__inst_mult_7_504 ;
wire Xd_0__inst_mult_7_505 ;
wire Xd_0__inst_mult_6_499 ;
wire Xd_0__inst_mult_6_500 ;
wire Xd_0__inst_mult_6_504 ;
wire Xd_0__inst_mult_6_505 ;
wire Xd_0__inst_mult_1_499 ;
wire Xd_0__inst_mult_1_500 ;
wire Xd_0__inst_mult_1_504 ;
wire Xd_0__inst_mult_1_505 ;
wire Xd_0__inst_mult_0_499 ;
wire Xd_0__inst_mult_0_500 ;
wire Xd_0__inst_mult_0_504 ;
wire Xd_0__inst_mult_0_505 ;
wire Xd_0__inst_mult_3_499 ;
wire Xd_0__inst_mult_3_500 ;
wire Xd_0__inst_mult_3_504 ;
wire Xd_0__inst_mult_3_505 ;
wire Xd_0__inst_mult_2_544 ;
wire Xd_0__inst_mult_2_545 ;
wire Xd_0__inst_mult_2_549 ;
wire Xd_0__inst_mult_2_550 ;
wire Xd_0__inst_mult_29_539 ;
wire Xd_0__inst_mult_29_540 ;
wire Xd_0__inst_mult_29_544 ;
wire Xd_0__inst_mult_29_545 ;
wire Xd_0__inst_mult_28_509 ;
wire Xd_0__inst_mult_28_510 ;
wire Xd_0__inst_mult_28_514 ;
wire Xd_0__inst_mult_28_515 ;
wire Xd_0__inst_mult_31_509 ;
wire Xd_0__inst_mult_31_510 ;
wire Xd_0__inst_mult_31_514 ;
wire Xd_0__inst_mult_31_515 ;
wire Xd_0__inst_mult_30_509 ;
wire Xd_0__inst_mult_30_510 ;
wire Xd_0__inst_mult_30_514 ;
wire Xd_0__inst_mult_30_515 ;
wire Xd_0__inst_mult_25_584 ;
wire Xd_0__inst_mult_25_585 ;
wire Xd_0__inst_mult_25_589 ;
wire Xd_0__inst_mult_25_590 ;
wire Xd_0__inst_mult_24_739 ;
wire Xd_0__inst_mult_24_740 ;
wire Xd_0__inst_mult_24_744 ;
wire Xd_0__inst_mult_24_745 ;
wire Xd_0__inst_mult_27_584 ;
wire Xd_0__inst_mult_27_585 ;
wire Xd_0__inst_mult_27_589 ;
wire Xd_0__inst_mult_27_590 ;
wire Xd_0__inst_mult_26_739 ;
wire Xd_0__inst_mult_26_740 ;
wire Xd_0__inst_mult_26_744 ;
wire Xd_0__inst_mult_26_745 ;
wire Xd_0__inst_mult_21_539 ;
wire Xd_0__inst_mult_21_540 ;
wire Xd_0__inst_mult_21_544 ;
wire Xd_0__inst_mult_21_545 ;
wire Xd_0__inst_mult_20_539 ;
wire Xd_0__inst_mult_20_540 ;
wire Xd_0__inst_mult_20_544 ;
wire Xd_0__inst_mult_20_545 ;
wire Xd_0__inst_mult_23_539 ;
wire Xd_0__inst_mult_23_540 ;
wire Xd_0__inst_mult_23_544 ;
wire Xd_0__inst_mult_23_545 ;
wire Xd_0__inst_mult_22_539 ;
wire Xd_0__inst_mult_22_540 ;
wire Xd_0__inst_mult_22_544 ;
wire Xd_0__inst_mult_22_545 ;
wire Xd_0__inst_mult_17_539 ;
wire Xd_0__inst_mult_17_540 ;
wire Xd_0__inst_mult_17_544 ;
wire Xd_0__inst_mult_17_545 ;
wire Xd_0__inst_mult_16_539 ;
wire Xd_0__inst_mult_16_540 ;
wire Xd_0__inst_mult_16_544 ;
wire Xd_0__inst_mult_16_545 ;
wire Xd_0__inst_mult_19_539 ;
wire Xd_0__inst_mult_19_540 ;
wire Xd_0__inst_mult_19_544 ;
wire Xd_0__inst_mult_19_545 ;
wire Xd_0__inst_mult_18_484 ;
wire Xd_0__inst_mult_18_485 ;
wire Xd_0__inst_mult_18_489 ;
wire Xd_0__inst_mult_18_490 ;
wire Xd_0__inst_mult_13_509 ;
wire Xd_0__inst_mult_13_510 ;
wire Xd_0__inst_mult_13_514 ;
wire Xd_0__inst_mult_13_515 ;
wire Xd_0__inst_mult_12_484 ;
wire Xd_0__inst_mult_12_485 ;
wire Xd_0__inst_mult_12_489 ;
wire Xd_0__inst_mult_12_490 ;
wire Xd_0__inst_mult_15_484 ;
wire Xd_0__inst_mult_15_485 ;
wire Xd_0__inst_mult_15_489 ;
wire Xd_0__inst_mult_15_490 ;
wire Xd_0__inst_mult_14_484 ;
wire Xd_0__inst_mult_14_485 ;
wire Xd_0__inst_mult_14_489 ;
wire Xd_0__inst_mult_14_490 ;
wire Xd_0__inst_mult_9_509 ;
wire Xd_0__inst_mult_9_510 ;
wire Xd_0__inst_mult_9_514 ;
wire Xd_0__inst_mult_9_515 ;
wire Xd_0__inst_mult_8_509 ;
wire Xd_0__inst_mult_8_510 ;
wire Xd_0__inst_mult_8_514 ;
wire Xd_0__inst_mult_8_515 ;
wire Xd_0__inst_mult_11_509 ;
wire Xd_0__inst_mult_11_510 ;
wire Xd_0__inst_mult_11_514 ;
wire Xd_0__inst_mult_11_515 ;
wire Xd_0__inst_mult_10_509 ;
wire Xd_0__inst_mult_10_510 ;
wire Xd_0__inst_mult_10_514 ;
wire Xd_0__inst_mult_10_515 ;
wire Xd_0__inst_mult_5_509 ;
wire Xd_0__inst_mult_5_510 ;
wire Xd_0__inst_mult_5_514 ;
wire Xd_0__inst_mult_5_515 ;
wire Xd_0__inst_mult_4_509 ;
wire Xd_0__inst_mult_4_510 ;
wire Xd_0__inst_mult_4_514 ;
wire Xd_0__inst_mult_4_515 ;
wire Xd_0__inst_mult_7_509 ;
wire Xd_0__inst_mult_7_510 ;
wire Xd_0__inst_mult_7_514 ;
wire Xd_0__inst_mult_7_515 ;
wire Xd_0__inst_mult_6_509 ;
wire Xd_0__inst_mult_6_510 ;
wire Xd_0__inst_mult_6_514 ;
wire Xd_0__inst_mult_6_515 ;
wire Xd_0__inst_mult_1_509 ;
wire Xd_0__inst_mult_1_510 ;
wire Xd_0__inst_mult_1_514 ;
wire Xd_0__inst_mult_1_515 ;
wire Xd_0__inst_mult_0_509 ;
wire Xd_0__inst_mult_0_510 ;
wire Xd_0__inst_mult_0_514 ;
wire Xd_0__inst_mult_0_515 ;
wire Xd_0__inst_mult_3_509 ;
wire Xd_0__inst_mult_3_510 ;
wire Xd_0__inst_mult_3_514 ;
wire Xd_0__inst_mult_3_515 ;
wire Xd_0__inst_mult_2_554 ;
wire Xd_0__inst_mult_2_555 ;
wire Xd_0__inst_mult_2_559 ;
wire Xd_0__inst_mult_2_560 ;
wire Xd_0__inst_mult_29_549 ;
wire Xd_0__inst_mult_29_550 ;
wire Xd_0__inst_mult_29_554 ;
wire Xd_0__inst_mult_29_555 ;
wire Xd_0__inst_mult_28_519 ;
wire Xd_0__inst_mult_28_520 ;
wire Xd_0__inst_mult_28_524 ;
wire Xd_0__inst_mult_28_525 ;
wire Xd_0__inst_mult_31_519 ;
wire Xd_0__inst_mult_31_520 ;
wire Xd_0__inst_mult_31_524 ;
wire Xd_0__inst_mult_31_525 ;
wire Xd_0__inst_mult_30_519 ;
wire Xd_0__inst_mult_30_520 ;
wire Xd_0__inst_mult_30_524 ;
wire Xd_0__inst_mult_30_525 ;
wire Xd_0__inst_mult_21_549 ;
wire Xd_0__inst_mult_21_550 ;
wire Xd_0__inst_mult_21_554 ;
wire Xd_0__inst_mult_21_555 ;
wire Xd_0__inst_mult_20_549 ;
wire Xd_0__inst_mult_20_550 ;
wire Xd_0__inst_mult_20_554 ;
wire Xd_0__inst_mult_20_555 ;
wire Xd_0__inst_mult_23_549 ;
wire Xd_0__inst_mult_23_550 ;
wire Xd_0__inst_mult_23_554 ;
wire Xd_0__inst_mult_23_555 ;
wire Xd_0__inst_mult_22_549 ;
wire Xd_0__inst_mult_22_550 ;
wire Xd_0__inst_mult_22_554 ;
wire Xd_0__inst_mult_22_555 ;
wire Xd_0__inst_mult_17_549 ;
wire Xd_0__inst_mult_17_550 ;
wire Xd_0__inst_mult_17_554 ;
wire Xd_0__inst_mult_17_555 ;
wire Xd_0__inst_mult_16_549 ;
wire Xd_0__inst_mult_16_550 ;
wire Xd_0__inst_mult_16_554 ;
wire Xd_0__inst_mult_16_555 ;
wire Xd_0__inst_mult_19_549 ;
wire Xd_0__inst_mult_19_550 ;
wire Xd_0__inst_mult_19_554 ;
wire Xd_0__inst_mult_19_555 ;
wire Xd_0__inst_mult_18_494 ;
wire Xd_0__inst_mult_18_495 ;
wire Xd_0__inst_mult_18_499 ;
wire Xd_0__inst_mult_18_500 ;
wire Xd_0__inst_mult_13_519 ;
wire Xd_0__inst_mult_13_520 ;
wire Xd_0__inst_mult_13_524 ;
wire Xd_0__inst_mult_13_525 ;
wire Xd_0__inst_mult_12_494 ;
wire Xd_0__inst_mult_12_495 ;
wire Xd_0__inst_mult_12_499 ;
wire Xd_0__inst_mult_12_500 ;
wire Xd_0__inst_mult_15_494 ;
wire Xd_0__inst_mult_15_495 ;
wire Xd_0__inst_mult_15_499 ;
wire Xd_0__inst_mult_15_500 ;
wire Xd_0__inst_mult_14_494 ;
wire Xd_0__inst_mult_14_495 ;
wire Xd_0__inst_mult_14_499 ;
wire Xd_0__inst_mult_14_500 ;
wire Xd_0__inst_mult_9_519 ;
wire Xd_0__inst_mult_9_520 ;
wire Xd_0__inst_mult_9_524 ;
wire Xd_0__inst_mult_9_525 ;
wire Xd_0__inst_mult_8_519 ;
wire Xd_0__inst_mult_8_520 ;
wire Xd_0__inst_mult_8_524 ;
wire Xd_0__inst_mult_8_525 ;
wire Xd_0__inst_mult_11_519 ;
wire Xd_0__inst_mult_11_520 ;
wire Xd_0__inst_mult_11_524 ;
wire Xd_0__inst_mult_11_525 ;
wire Xd_0__inst_mult_10_519 ;
wire Xd_0__inst_mult_10_520 ;
wire Xd_0__inst_mult_10_524 ;
wire Xd_0__inst_mult_10_525 ;
wire Xd_0__inst_mult_5_519 ;
wire Xd_0__inst_mult_5_520 ;
wire Xd_0__inst_mult_5_524 ;
wire Xd_0__inst_mult_5_525 ;
wire Xd_0__inst_mult_4_519 ;
wire Xd_0__inst_mult_4_520 ;
wire Xd_0__inst_mult_4_524 ;
wire Xd_0__inst_mult_4_525 ;
wire Xd_0__inst_mult_7_519 ;
wire Xd_0__inst_mult_7_520 ;
wire Xd_0__inst_mult_7_524 ;
wire Xd_0__inst_mult_7_525 ;
wire Xd_0__inst_mult_6_519 ;
wire Xd_0__inst_mult_6_520 ;
wire Xd_0__inst_mult_6_524 ;
wire Xd_0__inst_mult_6_525 ;
wire Xd_0__inst_mult_1_519 ;
wire Xd_0__inst_mult_1_520 ;
wire Xd_0__inst_mult_1_524 ;
wire Xd_0__inst_mult_1_525 ;
wire Xd_0__inst_mult_0_519 ;
wire Xd_0__inst_mult_0_520 ;
wire Xd_0__inst_mult_0_524 ;
wire Xd_0__inst_mult_0_525 ;
wire Xd_0__inst_mult_3_519 ;
wire Xd_0__inst_mult_3_520 ;
wire Xd_0__inst_mult_3_524 ;
wire Xd_0__inst_mult_3_525 ;
wire Xd_0__inst_mult_2_564 ;
wire Xd_0__inst_mult_2_565 ;
wire Xd_0__inst_mult_2_569 ;
wire Xd_0__inst_mult_2_570 ;
wire Xd_0__inst_mult_29_559 ;
wire Xd_0__inst_mult_29_560 ;
wire Xd_0__inst_mult_29_564 ;
wire Xd_0__inst_mult_29_565 ;
wire Xd_0__inst_mult_29_569 ;
wire Xd_0__inst_mult_29_570 ;
wire Xd_0__inst_mult_29_574 ;
wire Xd_0__inst_mult_29_575 ;
wire Xd_0__inst_mult_28_529 ;
wire Xd_0__inst_mult_28_530 ;
wire Xd_0__inst_mult_28_534 ;
wire Xd_0__inst_mult_28_535 ;
wire Xd_0__inst_mult_28_539 ;
wire Xd_0__inst_mult_28_540 ;
wire Xd_0__inst_mult_28_544 ;
wire Xd_0__inst_mult_28_545 ;
wire Xd_0__inst_mult_31_529 ;
wire Xd_0__inst_mult_31_530 ;
wire Xd_0__inst_mult_31_534 ;
wire Xd_0__inst_mult_31_535 ;
wire Xd_0__inst_mult_31_539 ;
wire Xd_0__inst_mult_31_540 ;
wire Xd_0__inst_mult_31_544 ;
wire Xd_0__inst_mult_31_545 ;
wire Xd_0__inst_mult_30_529 ;
wire Xd_0__inst_mult_30_530 ;
wire Xd_0__inst_mult_30_534 ;
wire Xd_0__inst_mult_30_535 ;
wire Xd_0__inst_mult_30_539 ;
wire Xd_0__inst_mult_30_540 ;
wire Xd_0__inst_mult_30_544 ;
wire Xd_0__inst_mult_30_545 ;
wire Xd_0__inst_mult_25_594 ;
wire Xd_0__inst_mult_25_595 ;
wire Xd_0__inst_mult_25_599 ;
wire Xd_0__inst_mult_25_600 ;
wire Xd_0__inst_mult_24_749 ;
wire Xd_0__inst_mult_24_750 ;
wire Xd_0__inst_mult_24_754 ;
wire Xd_0__inst_mult_24_755 ;
wire Xd_0__inst_mult_27_594 ;
wire Xd_0__inst_mult_27_595 ;
wire Xd_0__inst_mult_27_599 ;
wire Xd_0__inst_mult_27_600 ;
wire Xd_0__inst_mult_26_749 ;
wire Xd_0__inst_mult_26_750 ;
wire Xd_0__inst_mult_26_754 ;
wire Xd_0__inst_mult_26_755 ;
wire Xd_0__inst_mult_21_559 ;
wire Xd_0__inst_mult_21_560 ;
wire Xd_0__inst_mult_21_564 ;
wire Xd_0__inst_mult_21_565 ;
wire Xd_0__inst_mult_21_569 ;
wire Xd_0__inst_mult_21_570 ;
wire Xd_0__inst_mult_21_574 ;
wire Xd_0__inst_mult_21_575 ;
wire Xd_0__inst_mult_20_559 ;
wire Xd_0__inst_mult_20_560 ;
wire Xd_0__inst_mult_20_564 ;
wire Xd_0__inst_mult_20_565 ;
wire Xd_0__inst_mult_20_569 ;
wire Xd_0__inst_mult_20_570 ;
wire Xd_0__inst_mult_20_574 ;
wire Xd_0__inst_mult_20_575 ;
wire Xd_0__inst_mult_23_559 ;
wire Xd_0__inst_mult_23_560 ;
wire Xd_0__inst_mult_23_564 ;
wire Xd_0__inst_mult_23_565 ;
wire Xd_0__inst_mult_23_569 ;
wire Xd_0__inst_mult_23_570 ;
wire Xd_0__inst_mult_23_574 ;
wire Xd_0__inst_mult_23_575 ;
wire Xd_0__inst_mult_22_559 ;
wire Xd_0__inst_mult_22_560 ;
wire Xd_0__inst_mult_22_564 ;
wire Xd_0__inst_mult_22_565 ;
wire Xd_0__inst_mult_22_569 ;
wire Xd_0__inst_mult_22_570 ;
wire Xd_0__inst_mult_22_574 ;
wire Xd_0__inst_mult_22_575 ;
wire Xd_0__inst_mult_17_559 ;
wire Xd_0__inst_mult_17_560 ;
wire Xd_0__inst_mult_17_564 ;
wire Xd_0__inst_mult_17_565 ;
wire Xd_0__inst_mult_17_569 ;
wire Xd_0__inst_mult_17_570 ;
wire Xd_0__inst_mult_17_574 ;
wire Xd_0__inst_mult_17_575 ;
wire Xd_0__inst_mult_16_559 ;
wire Xd_0__inst_mult_16_560 ;
wire Xd_0__inst_mult_16_564 ;
wire Xd_0__inst_mult_16_565 ;
wire Xd_0__inst_mult_16_569 ;
wire Xd_0__inst_mult_16_570 ;
wire Xd_0__inst_mult_16_574 ;
wire Xd_0__inst_mult_16_575 ;
wire Xd_0__inst_mult_19_559 ;
wire Xd_0__inst_mult_19_560 ;
wire Xd_0__inst_mult_19_564 ;
wire Xd_0__inst_mult_19_565 ;
wire Xd_0__inst_mult_19_569 ;
wire Xd_0__inst_mult_19_570 ;
wire Xd_0__inst_mult_19_574 ;
wire Xd_0__inst_mult_19_575 ;
wire Xd_0__inst_mult_18_504 ;
wire Xd_0__inst_mult_18_505 ;
wire Xd_0__inst_mult_18_509 ;
wire Xd_0__inst_mult_18_510 ;
wire Xd_0__inst_mult_18_514 ;
wire Xd_0__inst_mult_18_515 ;
wire Xd_0__inst_mult_18_519 ;
wire Xd_0__inst_mult_18_520 ;
wire Xd_0__inst_mult_13_529 ;
wire Xd_0__inst_mult_13_530 ;
wire Xd_0__inst_mult_13_534 ;
wire Xd_0__inst_mult_13_535 ;
wire Xd_0__inst_mult_13_539 ;
wire Xd_0__inst_mult_13_540 ;
wire Xd_0__inst_mult_13_544 ;
wire Xd_0__inst_mult_13_545 ;
wire Xd_0__inst_mult_12_504 ;
wire Xd_0__inst_mult_12_505 ;
wire Xd_0__inst_mult_12_509 ;
wire Xd_0__inst_mult_12_510 ;
wire Xd_0__inst_mult_12_514 ;
wire Xd_0__inst_mult_12_515 ;
wire Xd_0__inst_mult_12_519 ;
wire Xd_0__inst_mult_12_520 ;
wire Xd_0__inst_mult_15_504 ;
wire Xd_0__inst_mult_15_505 ;
wire Xd_0__inst_mult_15_509 ;
wire Xd_0__inst_mult_15_510 ;
wire Xd_0__inst_mult_15_514 ;
wire Xd_0__inst_mult_15_515 ;
wire Xd_0__inst_mult_15_519 ;
wire Xd_0__inst_mult_15_520 ;
wire Xd_0__inst_mult_30_80_sumout ;
wire Xd_0__inst_mult_30_81 ;
wire Xd_0__inst_mult_14_504 ;
wire Xd_0__inst_mult_14_505 ;
wire Xd_0__inst_mult_14_509 ;
wire Xd_0__inst_mult_14_510 ;
wire Xd_0__inst_mult_14_514 ;
wire Xd_0__inst_mult_14_515 ;
wire Xd_0__inst_mult_14_519 ;
wire Xd_0__inst_mult_14_520 ;
wire Xd_0__inst_mult_23_80_sumout ;
wire Xd_0__inst_mult_23_81 ;
wire Xd_0__inst_mult_9_529 ;
wire Xd_0__inst_mult_9_530 ;
wire Xd_0__inst_mult_9_534 ;
wire Xd_0__inst_mult_9_535 ;
wire Xd_0__inst_mult_9_539 ;
wire Xd_0__inst_mult_9_540 ;
wire Xd_0__inst_mult_9_544 ;
wire Xd_0__inst_mult_9_545 ;
wire Xd_0__inst_mult_12_80_sumout ;
wire Xd_0__inst_mult_12_81 ;
wire Xd_0__inst_mult_8_529 ;
wire Xd_0__inst_mult_8_530 ;
wire Xd_0__inst_mult_8_534 ;
wire Xd_0__inst_mult_8_535 ;
wire Xd_0__inst_mult_8_539 ;
wire Xd_0__inst_mult_8_540 ;
wire Xd_0__inst_mult_8_544 ;
wire Xd_0__inst_mult_8_545 ;
wire Xd_0__inst_mult_11_529 ;
wire Xd_0__inst_mult_11_530 ;
wire Xd_0__inst_mult_11_534 ;
wire Xd_0__inst_mult_11_535 ;
wire Xd_0__inst_mult_11_539 ;
wire Xd_0__inst_mult_11_540 ;
wire Xd_0__inst_mult_11_544 ;
wire Xd_0__inst_mult_11_545 ;
wire Xd_0__inst_mult_10_529 ;
wire Xd_0__inst_mult_10_530 ;
wire Xd_0__inst_mult_10_534 ;
wire Xd_0__inst_mult_10_535 ;
wire Xd_0__inst_mult_10_539 ;
wire Xd_0__inst_mult_10_540 ;
wire Xd_0__inst_mult_10_544 ;
wire Xd_0__inst_mult_10_545 ;
wire Xd_0__inst_mult_5_529 ;
wire Xd_0__inst_mult_5_530 ;
wire Xd_0__inst_mult_5_534 ;
wire Xd_0__inst_mult_5_535 ;
wire Xd_0__inst_mult_5_539 ;
wire Xd_0__inst_mult_5_540 ;
wire Xd_0__inst_mult_5_544 ;
wire Xd_0__inst_mult_5_545 ;
wire Xd_0__inst_mult_4_529 ;
wire Xd_0__inst_mult_4_530 ;
wire Xd_0__inst_mult_4_534 ;
wire Xd_0__inst_mult_4_535 ;
wire Xd_0__inst_mult_4_539 ;
wire Xd_0__inst_mult_4_540 ;
wire Xd_0__inst_mult_4_544 ;
wire Xd_0__inst_mult_4_545 ;
wire Xd_0__inst_mult_7_529 ;
wire Xd_0__inst_mult_7_530 ;
wire Xd_0__inst_mult_7_534 ;
wire Xd_0__inst_mult_7_535 ;
wire Xd_0__inst_mult_7_539 ;
wire Xd_0__inst_mult_7_540 ;
wire Xd_0__inst_mult_7_544 ;
wire Xd_0__inst_mult_7_545 ;
wire Xd_0__inst_mult_6_529 ;
wire Xd_0__inst_mult_6_530 ;
wire Xd_0__inst_mult_6_534 ;
wire Xd_0__inst_mult_6_535 ;
wire Xd_0__inst_mult_6_539 ;
wire Xd_0__inst_mult_6_540 ;
wire Xd_0__inst_mult_6_544 ;
wire Xd_0__inst_mult_6_545 ;
wire Xd_0__inst_mult_1_529 ;
wire Xd_0__inst_mult_1_530 ;
wire Xd_0__inst_mult_1_534 ;
wire Xd_0__inst_mult_1_535 ;
wire Xd_0__inst_mult_1_539 ;
wire Xd_0__inst_mult_1_540 ;
wire Xd_0__inst_mult_1_544 ;
wire Xd_0__inst_mult_1_545 ;
wire Xd_0__inst_mult_0_529 ;
wire Xd_0__inst_mult_0_530 ;
wire Xd_0__inst_mult_0_534 ;
wire Xd_0__inst_mult_0_535 ;
wire Xd_0__inst_mult_0_539 ;
wire Xd_0__inst_mult_0_540 ;
wire Xd_0__inst_mult_0_544 ;
wire Xd_0__inst_mult_0_545 ;
wire Xd_0__inst_mult_3_529 ;
wire Xd_0__inst_mult_3_530 ;
wire Xd_0__inst_mult_3_534 ;
wire Xd_0__inst_mult_3_535 ;
wire Xd_0__inst_mult_3_539 ;
wire Xd_0__inst_mult_3_540 ;
wire Xd_0__inst_mult_3_544 ;
wire Xd_0__inst_mult_3_545 ;
wire Xd_0__inst_mult_2_574 ;
wire Xd_0__inst_mult_2_575 ;
wire Xd_0__inst_mult_2_579 ;
wire Xd_0__inst_mult_2_580 ;
wire Xd_0__inst_mult_2_584 ;
wire Xd_0__inst_mult_2_585 ;
wire Xd_0__inst_mult_2_589 ;
wire Xd_0__inst_mult_2_590 ;
wire Xd_0__inst_mult_29_579 ;
wire Xd_0__inst_mult_29_580 ;
wire Xd_0__inst_mult_29_584 ;
wire Xd_0__inst_mult_29_585 ;
wire Xd_0__inst_mult_29_589 ;
wire Xd_0__inst_mult_29_590 ;
wire Xd_0__inst_mult_29_594 ;
wire Xd_0__inst_mult_29_595 ;
wire Xd_0__inst_mult_28_549 ;
wire Xd_0__inst_mult_28_550 ;
wire Xd_0__inst_mult_28_554 ;
wire Xd_0__inst_mult_28_555 ;
wire Xd_0__inst_mult_28_559 ;
wire Xd_0__inst_mult_28_560 ;
wire Xd_0__inst_mult_28_564 ;
wire Xd_0__inst_mult_28_565 ;
wire Xd_0__inst_mult_31_549 ;
wire Xd_0__inst_mult_31_550 ;
wire Xd_0__inst_mult_31_554 ;
wire Xd_0__inst_mult_31_555 ;
wire Xd_0__inst_mult_31_559 ;
wire Xd_0__inst_mult_31_560 ;
wire Xd_0__inst_mult_31_564 ;
wire Xd_0__inst_mult_31_565 ;
wire Xd_0__inst_mult_30_549 ;
wire Xd_0__inst_mult_30_550 ;
wire Xd_0__inst_mult_30_554 ;
wire Xd_0__inst_mult_30_555 ;
wire Xd_0__inst_mult_30_559 ;
wire Xd_0__inst_mult_30_560 ;
wire Xd_0__inst_mult_30_564 ;
wire Xd_0__inst_mult_30_565 ;
wire Xd_0__inst_mult_25_604 ;
wire Xd_0__inst_mult_25_605 ;
wire Xd_0__inst_mult_25_609 ;
wire Xd_0__inst_mult_25_610 ;
wire Xd_0__inst_mult_24_759 ;
wire Xd_0__inst_mult_24_760 ;
wire Xd_0__inst_mult_24_764 ;
wire Xd_0__inst_mult_24_765 ;
wire Xd_0__inst_mult_27_604 ;
wire Xd_0__inst_mult_27_605 ;
wire Xd_0__inst_mult_27_609 ;
wire Xd_0__inst_mult_27_610 ;
wire Xd_0__inst_mult_26_759 ;
wire Xd_0__inst_mult_26_760 ;
wire Xd_0__inst_mult_26_764 ;
wire Xd_0__inst_mult_26_765 ;
wire Xd_0__inst_mult_21_579 ;
wire Xd_0__inst_mult_21_580 ;
wire Xd_0__inst_mult_21_584 ;
wire Xd_0__inst_mult_21_585 ;
wire Xd_0__inst_mult_21_589 ;
wire Xd_0__inst_mult_21_590 ;
wire Xd_0__inst_mult_21_594 ;
wire Xd_0__inst_mult_21_595 ;
wire Xd_0__inst_mult_20_579 ;
wire Xd_0__inst_mult_20_580 ;
wire Xd_0__inst_mult_20_584 ;
wire Xd_0__inst_mult_20_585 ;
wire Xd_0__inst_mult_20_589 ;
wire Xd_0__inst_mult_20_590 ;
wire Xd_0__inst_mult_20_594 ;
wire Xd_0__inst_mult_20_595 ;
wire Xd_0__inst_mult_23_579 ;
wire Xd_0__inst_mult_23_580 ;
wire Xd_0__inst_mult_23_584 ;
wire Xd_0__inst_mult_23_585 ;
wire Xd_0__inst_mult_23_589 ;
wire Xd_0__inst_mult_23_590 ;
wire Xd_0__inst_mult_23_594 ;
wire Xd_0__inst_mult_23_595 ;
wire Xd_0__inst_mult_22_579 ;
wire Xd_0__inst_mult_22_580 ;
wire Xd_0__inst_mult_22_584 ;
wire Xd_0__inst_mult_22_585 ;
wire Xd_0__inst_mult_22_589 ;
wire Xd_0__inst_mult_22_590 ;
wire Xd_0__inst_mult_22_594 ;
wire Xd_0__inst_mult_22_595 ;
wire Xd_0__inst_mult_17_579 ;
wire Xd_0__inst_mult_17_580 ;
wire Xd_0__inst_mult_17_584 ;
wire Xd_0__inst_mult_17_585 ;
wire Xd_0__inst_mult_17_589 ;
wire Xd_0__inst_mult_17_590 ;
wire Xd_0__inst_mult_17_594 ;
wire Xd_0__inst_mult_17_595 ;
wire Xd_0__inst_mult_16_579 ;
wire Xd_0__inst_mult_16_580 ;
wire Xd_0__inst_mult_16_584 ;
wire Xd_0__inst_mult_16_585 ;
wire Xd_0__inst_mult_16_589 ;
wire Xd_0__inst_mult_16_590 ;
wire Xd_0__inst_mult_16_594 ;
wire Xd_0__inst_mult_16_595 ;
wire Xd_0__inst_mult_19_579 ;
wire Xd_0__inst_mult_19_580 ;
wire Xd_0__inst_mult_19_584 ;
wire Xd_0__inst_mult_19_585 ;
wire Xd_0__inst_mult_19_589 ;
wire Xd_0__inst_mult_19_590 ;
wire Xd_0__inst_mult_19_594 ;
wire Xd_0__inst_mult_19_595 ;
wire Xd_0__inst_mult_18_524 ;
wire Xd_0__inst_mult_18_525 ;
wire Xd_0__inst_mult_18_529 ;
wire Xd_0__inst_mult_18_530 ;
wire Xd_0__inst_mult_18_534 ;
wire Xd_0__inst_mult_18_535 ;
wire Xd_0__inst_mult_18_539 ;
wire Xd_0__inst_mult_18_540 ;
wire Xd_0__inst_mult_13_549 ;
wire Xd_0__inst_mult_13_550 ;
wire Xd_0__inst_mult_13_554 ;
wire Xd_0__inst_mult_13_555 ;
wire Xd_0__inst_mult_13_559 ;
wire Xd_0__inst_mult_13_560 ;
wire Xd_0__inst_mult_13_564 ;
wire Xd_0__inst_mult_13_565 ;
wire Xd_0__inst_mult_12_524 ;
wire Xd_0__inst_mult_12_525 ;
wire Xd_0__inst_mult_12_529 ;
wire Xd_0__inst_mult_12_530 ;
wire Xd_0__inst_mult_12_534 ;
wire Xd_0__inst_mult_12_535 ;
wire Xd_0__inst_mult_12_539 ;
wire Xd_0__inst_mult_12_540 ;
wire Xd_0__inst_mult_15_524 ;
wire Xd_0__inst_mult_15_525 ;
wire Xd_0__inst_mult_15_529 ;
wire Xd_0__inst_mult_15_530 ;
wire Xd_0__inst_mult_15_534 ;
wire Xd_0__inst_mult_15_535 ;
wire Xd_0__inst_mult_15_539 ;
wire Xd_0__inst_mult_15_540 ;
wire Xd_0__inst_mult_14_524 ;
wire Xd_0__inst_mult_14_525 ;
wire Xd_0__inst_mult_14_529 ;
wire Xd_0__inst_mult_14_530 ;
wire Xd_0__inst_mult_14_534 ;
wire Xd_0__inst_mult_14_535 ;
wire Xd_0__inst_mult_14_539 ;
wire Xd_0__inst_mult_14_540 ;
wire Xd_0__inst_mult_9_549 ;
wire Xd_0__inst_mult_9_550 ;
wire Xd_0__inst_mult_9_554 ;
wire Xd_0__inst_mult_9_555 ;
wire Xd_0__inst_mult_9_559 ;
wire Xd_0__inst_mult_9_560 ;
wire Xd_0__inst_mult_9_564 ;
wire Xd_0__inst_mult_9_565 ;
wire Xd_0__inst_mult_8_549 ;
wire Xd_0__inst_mult_8_550 ;
wire Xd_0__inst_mult_8_554 ;
wire Xd_0__inst_mult_8_555 ;
wire Xd_0__inst_mult_8_559 ;
wire Xd_0__inst_mult_8_560 ;
wire Xd_0__inst_mult_8_564 ;
wire Xd_0__inst_mult_8_565 ;
wire Xd_0__inst_mult_11_549 ;
wire Xd_0__inst_mult_11_550 ;
wire Xd_0__inst_mult_11_554 ;
wire Xd_0__inst_mult_11_555 ;
wire Xd_0__inst_mult_11_559 ;
wire Xd_0__inst_mult_11_560 ;
wire Xd_0__inst_mult_11_564 ;
wire Xd_0__inst_mult_11_565 ;
wire Xd_0__inst_mult_10_549 ;
wire Xd_0__inst_mult_10_550 ;
wire Xd_0__inst_mult_10_554 ;
wire Xd_0__inst_mult_10_555 ;
wire Xd_0__inst_mult_10_559 ;
wire Xd_0__inst_mult_10_560 ;
wire Xd_0__inst_mult_10_564 ;
wire Xd_0__inst_mult_10_565 ;
wire Xd_0__inst_mult_5_549 ;
wire Xd_0__inst_mult_5_550 ;
wire Xd_0__inst_mult_5_554 ;
wire Xd_0__inst_mult_5_555 ;
wire Xd_0__inst_mult_5_559 ;
wire Xd_0__inst_mult_5_560 ;
wire Xd_0__inst_mult_5_564 ;
wire Xd_0__inst_mult_5_565 ;
wire Xd_0__inst_mult_4_549 ;
wire Xd_0__inst_mult_4_550 ;
wire Xd_0__inst_mult_4_554 ;
wire Xd_0__inst_mult_4_555 ;
wire Xd_0__inst_mult_4_559 ;
wire Xd_0__inst_mult_4_560 ;
wire Xd_0__inst_mult_4_564 ;
wire Xd_0__inst_mult_4_565 ;
wire Xd_0__inst_mult_7_549 ;
wire Xd_0__inst_mult_7_550 ;
wire Xd_0__inst_mult_7_554 ;
wire Xd_0__inst_mult_7_555 ;
wire Xd_0__inst_mult_7_559 ;
wire Xd_0__inst_mult_7_560 ;
wire Xd_0__inst_mult_7_564 ;
wire Xd_0__inst_mult_7_565 ;
wire Xd_0__inst_mult_6_549 ;
wire Xd_0__inst_mult_6_550 ;
wire Xd_0__inst_mult_6_554 ;
wire Xd_0__inst_mult_6_555 ;
wire Xd_0__inst_mult_6_559 ;
wire Xd_0__inst_mult_6_560 ;
wire Xd_0__inst_mult_6_564 ;
wire Xd_0__inst_mult_6_565 ;
wire Xd_0__inst_mult_1_549 ;
wire Xd_0__inst_mult_1_550 ;
wire Xd_0__inst_mult_1_554 ;
wire Xd_0__inst_mult_1_555 ;
wire Xd_0__inst_mult_1_559 ;
wire Xd_0__inst_mult_1_560 ;
wire Xd_0__inst_mult_1_564 ;
wire Xd_0__inst_mult_1_565 ;
wire Xd_0__inst_mult_0_549 ;
wire Xd_0__inst_mult_0_550 ;
wire Xd_0__inst_mult_0_554 ;
wire Xd_0__inst_mult_0_555 ;
wire Xd_0__inst_mult_0_559 ;
wire Xd_0__inst_mult_0_560 ;
wire Xd_0__inst_mult_0_564 ;
wire Xd_0__inst_mult_0_565 ;
wire Xd_0__inst_mult_3_549 ;
wire Xd_0__inst_mult_3_550 ;
wire Xd_0__inst_mult_3_554 ;
wire Xd_0__inst_mult_3_555 ;
wire Xd_0__inst_mult_3_559 ;
wire Xd_0__inst_mult_3_560 ;
wire Xd_0__inst_mult_3_564 ;
wire Xd_0__inst_mult_3_565 ;
wire Xd_0__inst_mult_2_594 ;
wire Xd_0__inst_mult_2_595 ;
wire Xd_0__inst_mult_2_599 ;
wire Xd_0__inst_mult_2_600 ;
wire Xd_0__inst_mult_2_604 ;
wire Xd_0__inst_mult_2_605 ;
wire Xd_0__inst_mult_2_609 ;
wire Xd_0__inst_mult_2_610 ;
wire Xd_0__inst_mult_29_599 ;
wire Xd_0__inst_mult_29_600 ;
wire Xd_0__inst_mult_29_604 ;
wire Xd_0__inst_mult_29_605 ;
wire Xd_0__inst_mult_28_569 ;
wire Xd_0__inst_mult_28_570 ;
wire Xd_0__inst_mult_28_574 ;
wire Xd_0__inst_mult_28_575 ;
wire Xd_0__inst_mult_28_579 ;
wire Xd_0__inst_mult_28_580 ;
wire Xd_0__inst_mult_28_584 ;
wire Xd_0__inst_mult_28_585 ;
wire Xd_0__inst_mult_31_569 ;
wire Xd_0__inst_mult_31_570 ;
wire Xd_0__inst_mult_31_574 ;
wire Xd_0__inst_mult_31_575 ;
wire Xd_0__inst_mult_31_579 ;
wire Xd_0__inst_mult_31_580 ;
wire Xd_0__inst_mult_31_584 ;
wire Xd_0__inst_mult_31_585 ;
wire Xd_0__inst_mult_30_569 ;
wire Xd_0__inst_mult_30_570 ;
wire Xd_0__inst_mult_30_574 ;
wire Xd_0__inst_mult_30_575 ;
wire Xd_0__inst_mult_30_579 ;
wire Xd_0__inst_mult_30_580 ;
wire Xd_0__inst_mult_30_584 ;
wire Xd_0__inst_mult_30_585 ;
wire Xd_0__inst_mult_25_614 ;
wire Xd_0__inst_mult_25_615 ;
wire Xd_0__inst_mult_25_619 ;
wire Xd_0__inst_mult_25_620 ;
wire Xd_0__inst_mult_24_769 ;
wire Xd_0__inst_mult_24_770 ;
wire Xd_0__inst_mult_27_614 ;
wire Xd_0__inst_mult_27_615 ;
wire Xd_0__inst_mult_27_619 ;
wire Xd_0__inst_mult_27_620 ;
wire Xd_0__inst_mult_26_769 ;
wire Xd_0__inst_mult_26_770 ;
wire Xd_0__inst_mult_21_599 ;
wire Xd_0__inst_mult_21_600 ;
wire Xd_0__inst_mult_21_604 ;
wire Xd_0__inst_mult_21_605 ;
wire Xd_0__inst_mult_20_599 ;
wire Xd_0__inst_mult_20_600 ;
wire Xd_0__inst_mult_20_604 ;
wire Xd_0__inst_mult_20_605 ;
wire Xd_0__inst_mult_23_599 ;
wire Xd_0__inst_mult_23_600 ;
wire Xd_0__inst_mult_23_604 ;
wire Xd_0__inst_mult_23_605 ;
wire Xd_0__inst_mult_22_599 ;
wire Xd_0__inst_mult_22_600 ;
wire Xd_0__inst_mult_22_604 ;
wire Xd_0__inst_mult_22_605 ;
wire Xd_0__inst_mult_17_599 ;
wire Xd_0__inst_mult_17_600 ;
wire Xd_0__inst_mult_17_604 ;
wire Xd_0__inst_mult_17_605 ;
wire Xd_0__inst_mult_16_599 ;
wire Xd_0__inst_mult_16_600 ;
wire Xd_0__inst_mult_16_604 ;
wire Xd_0__inst_mult_16_605 ;
wire Xd_0__inst_mult_19_599 ;
wire Xd_0__inst_mult_19_600 ;
wire Xd_0__inst_mult_19_604 ;
wire Xd_0__inst_mult_19_605 ;
wire Xd_0__inst_mult_18_544 ;
wire Xd_0__inst_mult_18_545 ;
wire Xd_0__inst_mult_18_549 ;
wire Xd_0__inst_mult_18_550 ;
wire Xd_0__inst_mult_18_554 ;
wire Xd_0__inst_mult_18_555 ;
wire Xd_0__inst_mult_18_559 ;
wire Xd_0__inst_mult_18_560 ;
wire Xd_0__inst_mult_13_569 ;
wire Xd_0__inst_mult_13_570 ;
wire Xd_0__inst_mult_13_574 ;
wire Xd_0__inst_mult_13_575 ;
wire Xd_0__inst_mult_13_579 ;
wire Xd_0__inst_mult_13_580 ;
wire Xd_0__inst_mult_13_584 ;
wire Xd_0__inst_mult_13_585 ;
wire Xd_0__inst_mult_12_544 ;
wire Xd_0__inst_mult_12_545 ;
wire Xd_0__inst_mult_12_549 ;
wire Xd_0__inst_mult_12_550 ;
wire Xd_0__inst_mult_12_554 ;
wire Xd_0__inst_mult_12_555 ;
wire Xd_0__inst_mult_12_559 ;
wire Xd_0__inst_mult_12_560 ;
wire Xd_0__inst_mult_15_544 ;
wire Xd_0__inst_mult_15_545 ;
wire Xd_0__inst_mult_15_549 ;
wire Xd_0__inst_mult_15_550 ;
wire Xd_0__inst_mult_15_554 ;
wire Xd_0__inst_mult_15_555 ;
wire Xd_0__inst_mult_15_559 ;
wire Xd_0__inst_mult_15_560 ;
wire Xd_0__inst_mult_14_544 ;
wire Xd_0__inst_mult_14_545 ;
wire Xd_0__inst_mult_14_549 ;
wire Xd_0__inst_mult_14_550 ;
wire Xd_0__inst_mult_14_554 ;
wire Xd_0__inst_mult_14_555 ;
wire Xd_0__inst_mult_14_559 ;
wire Xd_0__inst_mult_14_560 ;
wire Xd_0__inst_mult_9_569 ;
wire Xd_0__inst_mult_9_570 ;
wire Xd_0__inst_mult_9_574 ;
wire Xd_0__inst_mult_9_575 ;
wire Xd_0__inst_mult_9_579 ;
wire Xd_0__inst_mult_9_580 ;
wire Xd_0__inst_mult_9_584 ;
wire Xd_0__inst_mult_9_585 ;
wire Xd_0__inst_mult_8_569 ;
wire Xd_0__inst_mult_8_570 ;
wire Xd_0__inst_mult_8_574 ;
wire Xd_0__inst_mult_8_575 ;
wire Xd_0__inst_mult_8_579 ;
wire Xd_0__inst_mult_8_580 ;
wire Xd_0__inst_mult_8_584 ;
wire Xd_0__inst_mult_8_585 ;
wire Xd_0__inst_mult_11_569 ;
wire Xd_0__inst_mult_11_570 ;
wire Xd_0__inst_mult_11_574 ;
wire Xd_0__inst_mult_11_575 ;
wire Xd_0__inst_mult_11_579 ;
wire Xd_0__inst_mult_11_580 ;
wire Xd_0__inst_mult_11_584 ;
wire Xd_0__inst_mult_11_585 ;
wire Xd_0__inst_mult_10_569 ;
wire Xd_0__inst_mult_10_570 ;
wire Xd_0__inst_mult_10_574 ;
wire Xd_0__inst_mult_10_575 ;
wire Xd_0__inst_mult_10_579 ;
wire Xd_0__inst_mult_10_580 ;
wire Xd_0__inst_mult_10_584 ;
wire Xd_0__inst_mult_10_585 ;
wire Xd_0__inst_mult_5_569 ;
wire Xd_0__inst_mult_5_570 ;
wire Xd_0__inst_mult_5_574 ;
wire Xd_0__inst_mult_5_575 ;
wire Xd_0__inst_mult_5_579 ;
wire Xd_0__inst_mult_5_580 ;
wire Xd_0__inst_mult_5_584 ;
wire Xd_0__inst_mult_5_585 ;
wire Xd_0__inst_mult_4_569 ;
wire Xd_0__inst_mult_4_570 ;
wire Xd_0__inst_mult_4_574 ;
wire Xd_0__inst_mult_4_575 ;
wire Xd_0__inst_mult_4_579 ;
wire Xd_0__inst_mult_4_580 ;
wire Xd_0__inst_mult_4_584 ;
wire Xd_0__inst_mult_4_585 ;
wire Xd_0__inst_mult_7_569 ;
wire Xd_0__inst_mult_7_570 ;
wire Xd_0__inst_mult_7_574 ;
wire Xd_0__inst_mult_7_575 ;
wire Xd_0__inst_mult_7_579 ;
wire Xd_0__inst_mult_7_580 ;
wire Xd_0__inst_mult_7_584 ;
wire Xd_0__inst_mult_7_585 ;
wire Xd_0__inst_mult_6_569 ;
wire Xd_0__inst_mult_6_570 ;
wire Xd_0__inst_mult_6_574 ;
wire Xd_0__inst_mult_6_575 ;
wire Xd_0__inst_mult_6_579 ;
wire Xd_0__inst_mult_6_580 ;
wire Xd_0__inst_mult_6_584 ;
wire Xd_0__inst_mult_6_585 ;
wire Xd_0__inst_mult_1_569 ;
wire Xd_0__inst_mult_1_570 ;
wire Xd_0__inst_mult_1_574 ;
wire Xd_0__inst_mult_1_575 ;
wire Xd_0__inst_mult_1_579 ;
wire Xd_0__inst_mult_1_580 ;
wire Xd_0__inst_mult_1_584 ;
wire Xd_0__inst_mult_1_585 ;
wire Xd_0__inst_mult_0_569 ;
wire Xd_0__inst_mult_0_570 ;
wire Xd_0__inst_mult_0_574 ;
wire Xd_0__inst_mult_0_575 ;
wire Xd_0__inst_mult_0_579 ;
wire Xd_0__inst_mult_0_580 ;
wire Xd_0__inst_mult_0_584 ;
wire Xd_0__inst_mult_0_585 ;
wire Xd_0__inst_mult_3_569 ;
wire Xd_0__inst_mult_3_570 ;
wire Xd_0__inst_mult_3_574 ;
wire Xd_0__inst_mult_3_575 ;
wire Xd_0__inst_mult_3_579 ;
wire Xd_0__inst_mult_3_580 ;
wire Xd_0__inst_mult_3_584 ;
wire Xd_0__inst_mult_3_585 ;
wire Xd_0__inst_mult_2_614 ;
wire Xd_0__inst_mult_2_615 ;
wire Xd_0__inst_mult_2_619 ;
wire Xd_0__inst_mult_2_620 ;
wire Xd_0__inst_mult_2_624 ;
wire Xd_0__inst_mult_2_625 ;
wire Xd_0__inst_mult_2_629 ;
wire Xd_0__inst_mult_2_630 ;
wire Xd_0__inst_mult_29_609 ;
wire Xd_0__inst_mult_29_610 ;
wire Xd_0__inst_mult_29_614 ;
wire Xd_0__inst_mult_29_615 ;
wire Xd_0__inst_mult_28_589 ;
wire Xd_0__inst_mult_28_590 ;
wire Xd_0__inst_mult_28_594 ;
wire Xd_0__inst_mult_28_595 ;
wire Xd_0__inst_mult_28_599 ;
wire Xd_0__inst_mult_28_600 ;
wire Xd_0__inst_mult_28_604 ;
wire Xd_0__inst_mult_28_605 ;
wire Xd_0__inst_mult_31_589 ;
wire Xd_0__inst_mult_31_590 ;
wire Xd_0__inst_mult_31_594 ;
wire Xd_0__inst_mult_31_595 ;
wire Xd_0__inst_mult_31_599 ;
wire Xd_0__inst_mult_31_600 ;
wire Xd_0__inst_mult_31_604 ;
wire Xd_0__inst_mult_31_605 ;
wire Xd_0__inst_mult_30_589 ;
wire Xd_0__inst_mult_30_590 ;
wire Xd_0__inst_mult_30_594 ;
wire Xd_0__inst_mult_30_595 ;
wire Xd_0__inst_mult_30_599 ;
wire Xd_0__inst_mult_30_600 ;
wire Xd_0__inst_mult_30_604 ;
wire Xd_0__inst_mult_30_605 ;
wire Xd_0__inst_mult_25_624 ;
wire Xd_0__inst_mult_25_625 ;
wire Xd_0__inst_mult_25_629 ;
wire Xd_0__inst_mult_25_630 ;
wire Xd_0__inst_mult_27_624 ;
wire Xd_0__inst_mult_27_625 ;
wire Xd_0__inst_mult_27_629 ;
wire Xd_0__inst_mult_27_630 ;
wire Xd_0__inst_mult_21_609 ;
wire Xd_0__inst_mult_21_610 ;
wire Xd_0__inst_mult_21_614 ;
wire Xd_0__inst_mult_21_615 ;
wire Xd_0__inst_mult_20_609 ;
wire Xd_0__inst_mult_20_610 ;
wire Xd_0__inst_mult_20_614 ;
wire Xd_0__inst_mult_20_615 ;
wire Xd_0__inst_mult_23_609 ;
wire Xd_0__inst_mult_23_610 ;
wire Xd_0__inst_mult_23_614 ;
wire Xd_0__inst_mult_23_615 ;
wire Xd_0__inst_mult_22_609 ;
wire Xd_0__inst_mult_22_610 ;
wire Xd_0__inst_mult_22_614 ;
wire Xd_0__inst_mult_22_615 ;
wire Xd_0__inst_mult_17_609 ;
wire Xd_0__inst_mult_17_610 ;
wire Xd_0__inst_mult_17_614 ;
wire Xd_0__inst_mult_17_615 ;
wire Xd_0__inst_mult_16_609 ;
wire Xd_0__inst_mult_16_610 ;
wire Xd_0__inst_mult_16_614 ;
wire Xd_0__inst_mult_16_615 ;
wire Xd_0__inst_mult_19_609 ;
wire Xd_0__inst_mult_19_610 ;
wire Xd_0__inst_mult_19_614 ;
wire Xd_0__inst_mult_19_615 ;
wire Xd_0__inst_mult_18_564 ;
wire Xd_0__inst_mult_18_565 ;
wire Xd_0__inst_mult_18_569 ;
wire Xd_0__inst_mult_18_570 ;
wire Xd_0__inst_mult_18_574 ;
wire Xd_0__inst_mult_18_575 ;
wire Xd_0__inst_mult_18_579 ;
wire Xd_0__inst_mult_18_580 ;
wire Xd_0__inst_mult_13_589 ;
wire Xd_0__inst_mult_13_590 ;
wire Xd_0__inst_mult_13_594 ;
wire Xd_0__inst_mult_13_595 ;
wire Xd_0__inst_mult_13_599 ;
wire Xd_0__inst_mult_13_600 ;
wire Xd_0__inst_mult_13_604 ;
wire Xd_0__inst_mult_13_605 ;
wire Xd_0__inst_mult_12_564 ;
wire Xd_0__inst_mult_12_565 ;
wire Xd_0__inst_mult_12_569 ;
wire Xd_0__inst_mult_12_570 ;
wire Xd_0__inst_mult_12_574 ;
wire Xd_0__inst_mult_12_575 ;
wire Xd_0__inst_mult_12_579 ;
wire Xd_0__inst_mult_12_580 ;
wire Xd_0__inst_mult_15_564 ;
wire Xd_0__inst_mult_15_565 ;
wire Xd_0__inst_mult_15_569 ;
wire Xd_0__inst_mult_15_570 ;
wire Xd_0__inst_mult_15_574 ;
wire Xd_0__inst_mult_15_575 ;
wire Xd_0__inst_mult_15_579 ;
wire Xd_0__inst_mult_15_580 ;
wire Xd_0__inst_mult_14_564 ;
wire Xd_0__inst_mult_14_565 ;
wire Xd_0__inst_mult_14_569 ;
wire Xd_0__inst_mult_14_570 ;
wire Xd_0__inst_mult_14_574 ;
wire Xd_0__inst_mult_14_575 ;
wire Xd_0__inst_mult_14_579 ;
wire Xd_0__inst_mult_14_580 ;
wire Xd_0__inst_mult_9_589 ;
wire Xd_0__inst_mult_9_590 ;
wire Xd_0__inst_mult_9_594 ;
wire Xd_0__inst_mult_9_595 ;
wire Xd_0__inst_mult_9_599 ;
wire Xd_0__inst_mult_9_600 ;
wire Xd_0__inst_mult_9_604 ;
wire Xd_0__inst_mult_9_605 ;
wire Xd_0__inst_mult_8_589 ;
wire Xd_0__inst_mult_8_590 ;
wire Xd_0__inst_mult_8_594 ;
wire Xd_0__inst_mult_8_595 ;
wire Xd_0__inst_mult_8_599 ;
wire Xd_0__inst_mult_8_600 ;
wire Xd_0__inst_mult_8_604 ;
wire Xd_0__inst_mult_8_605 ;
wire Xd_0__inst_mult_11_589 ;
wire Xd_0__inst_mult_11_590 ;
wire Xd_0__inst_mult_11_594 ;
wire Xd_0__inst_mult_11_595 ;
wire Xd_0__inst_mult_11_599 ;
wire Xd_0__inst_mult_11_600 ;
wire Xd_0__inst_mult_11_604 ;
wire Xd_0__inst_mult_11_605 ;
wire Xd_0__inst_mult_10_589 ;
wire Xd_0__inst_mult_10_590 ;
wire Xd_0__inst_mult_10_594 ;
wire Xd_0__inst_mult_10_595 ;
wire Xd_0__inst_mult_10_599 ;
wire Xd_0__inst_mult_10_600 ;
wire Xd_0__inst_mult_10_604 ;
wire Xd_0__inst_mult_10_605 ;
wire Xd_0__inst_mult_5_589 ;
wire Xd_0__inst_mult_5_590 ;
wire Xd_0__inst_mult_5_594 ;
wire Xd_0__inst_mult_5_595 ;
wire Xd_0__inst_mult_5_599 ;
wire Xd_0__inst_mult_5_600 ;
wire Xd_0__inst_mult_5_604 ;
wire Xd_0__inst_mult_5_605 ;
wire Xd_0__inst_mult_4_589 ;
wire Xd_0__inst_mult_4_590 ;
wire Xd_0__inst_mult_4_594 ;
wire Xd_0__inst_mult_4_595 ;
wire Xd_0__inst_mult_4_599 ;
wire Xd_0__inst_mult_4_600 ;
wire Xd_0__inst_mult_4_604 ;
wire Xd_0__inst_mult_4_605 ;
wire Xd_0__inst_mult_7_589 ;
wire Xd_0__inst_mult_7_590 ;
wire Xd_0__inst_mult_7_594 ;
wire Xd_0__inst_mult_7_595 ;
wire Xd_0__inst_mult_7_599 ;
wire Xd_0__inst_mult_7_600 ;
wire Xd_0__inst_mult_7_604 ;
wire Xd_0__inst_mult_7_605 ;
wire Xd_0__inst_mult_6_589 ;
wire Xd_0__inst_mult_6_590 ;
wire Xd_0__inst_mult_6_594 ;
wire Xd_0__inst_mult_6_595 ;
wire Xd_0__inst_mult_6_599 ;
wire Xd_0__inst_mult_6_600 ;
wire Xd_0__inst_mult_6_604 ;
wire Xd_0__inst_mult_6_605 ;
wire Xd_0__inst_mult_1_589 ;
wire Xd_0__inst_mult_1_590 ;
wire Xd_0__inst_mult_1_594 ;
wire Xd_0__inst_mult_1_595 ;
wire Xd_0__inst_mult_1_599 ;
wire Xd_0__inst_mult_1_600 ;
wire Xd_0__inst_mult_1_604 ;
wire Xd_0__inst_mult_1_605 ;
wire Xd_0__inst_mult_0_589 ;
wire Xd_0__inst_mult_0_590 ;
wire Xd_0__inst_mult_0_594 ;
wire Xd_0__inst_mult_0_595 ;
wire Xd_0__inst_mult_0_599 ;
wire Xd_0__inst_mult_0_600 ;
wire Xd_0__inst_mult_0_604 ;
wire Xd_0__inst_mult_0_605 ;
wire Xd_0__inst_mult_3_589 ;
wire Xd_0__inst_mult_3_590 ;
wire Xd_0__inst_mult_3_594 ;
wire Xd_0__inst_mult_3_595 ;
wire Xd_0__inst_mult_3_599 ;
wire Xd_0__inst_mult_3_600 ;
wire Xd_0__inst_mult_3_604 ;
wire Xd_0__inst_mult_3_605 ;
wire Xd_0__inst_mult_2_634 ;
wire Xd_0__inst_mult_2_635 ;
wire Xd_0__inst_mult_2_639 ;
wire Xd_0__inst_mult_2_640 ;
wire Xd_0__inst_mult_2_644 ;
wire Xd_0__inst_mult_2_645 ;
wire Xd_0__inst_mult_2_649 ;
wire Xd_0__inst_mult_2_650 ;
wire Xd_0__inst_mult_29_619 ;
wire Xd_0__inst_mult_29_620 ;
wire Xd_0__inst_mult_29_624 ;
wire Xd_0__inst_mult_29_625 ;
wire Xd_0__inst_mult_28_609 ;
wire Xd_0__inst_mult_28_610 ;
wire Xd_0__inst_mult_28_614 ;
wire Xd_0__inst_mult_28_615 ;
wire Xd_0__inst_mult_31_609 ;
wire Xd_0__inst_mult_31_610 ;
wire Xd_0__inst_mult_31_614 ;
wire Xd_0__inst_mult_31_615 ;
wire Xd_0__inst_mult_30_609 ;
wire Xd_0__inst_mult_30_610 ;
wire Xd_0__inst_mult_30_614 ;
wire Xd_0__inst_mult_30_615 ;
wire Xd_0__inst_mult_25_634 ;
wire Xd_0__inst_mult_25_635 ;
wire Xd_0__inst_mult_25_639 ;
wire Xd_0__inst_mult_25_640 ;
wire Xd_0__inst_mult_27_634 ;
wire Xd_0__inst_mult_27_635 ;
wire Xd_0__inst_mult_27_639 ;
wire Xd_0__inst_mult_27_640 ;
wire Xd_0__inst_mult_21_619 ;
wire Xd_0__inst_mult_21_620 ;
wire Xd_0__inst_mult_21_624 ;
wire Xd_0__inst_mult_21_625 ;
wire Xd_0__inst_mult_20_619 ;
wire Xd_0__inst_mult_20_620 ;
wire Xd_0__inst_mult_20_624 ;
wire Xd_0__inst_mult_20_625 ;
wire Xd_0__inst_mult_23_619 ;
wire Xd_0__inst_mult_23_620 ;
wire Xd_0__inst_mult_23_624 ;
wire Xd_0__inst_mult_23_625 ;
wire Xd_0__inst_mult_22_619 ;
wire Xd_0__inst_mult_22_620 ;
wire Xd_0__inst_mult_22_624 ;
wire Xd_0__inst_mult_22_625 ;
wire Xd_0__inst_mult_17_619 ;
wire Xd_0__inst_mult_17_620 ;
wire Xd_0__inst_mult_17_624 ;
wire Xd_0__inst_mult_17_625 ;
wire Xd_0__inst_mult_16_619 ;
wire Xd_0__inst_mult_16_620 ;
wire Xd_0__inst_mult_16_624 ;
wire Xd_0__inst_mult_16_625 ;
wire Xd_0__inst_mult_19_619 ;
wire Xd_0__inst_mult_19_620 ;
wire Xd_0__inst_mult_19_624 ;
wire Xd_0__inst_mult_19_625 ;
wire Xd_0__inst_mult_18_584 ;
wire Xd_0__inst_mult_18_589 ;
wire Xd_0__inst_mult_18_590 ;
wire Xd_0__inst_mult_18_594 ;
wire Xd_0__inst_mult_18_595 ;
wire Xd_0__inst_mult_18_599 ;
wire Xd_0__inst_mult_18_600 ;
wire Xd_0__inst_mult_13_609 ;
wire Xd_0__inst_mult_13_610 ;
wire Xd_0__inst_mult_13_614 ;
wire Xd_0__inst_mult_13_615 ;
wire Xd_0__inst_mult_12_584 ;
wire Xd_0__inst_mult_12_589 ;
wire Xd_0__inst_mult_12_590 ;
wire Xd_0__inst_mult_12_594 ;
wire Xd_0__inst_mult_12_595 ;
wire Xd_0__inst_mult_12_599 ;
wire Xd_0__inst_mult_12_600 ;
wire Xd_0__inst_mult_15_584 ;
wire Xd_0__inst_mult_15_589 ;
wire Xd_0__inst_mult_15_590 ;
wire Xd_0__inst_mult_15_594 ;
wire Xd_0__inst_mult_15_595 ;
wire Xd_0__inst_mult_15_599 ;
wire Xd_0__inst_mult_15_600 ;
wire Xd_0__inst_mult_14_584 ;
wire Xd_0__inst_mult_14_589 ;
wire Xd_0__inst_mult_14_590 ;
wire Xd_0__inst_mult_14_594 ;
wire Xd_0__inst_mult_14_595 ;
wire Xd_0__inst_mult_14_599 ;
wire Xd_0__inst_mult_14_600 ;
wire Xd_0__inst_mult_9_609 ;
wire Xd_0__inst_mult_9_610 ;
wire Xd_0__inst_mult_9_614 ;
wire Xd_0__inst_mult_9_615 ;
wire Xd_0__inst_mult_8_609 ;
wire Xd_0__inst_mult_8_610 ;
wire Xd_0__inst_mult_8_614 ;
wire Xd_0__inst_mult_8_615 ;
wire Xd_0__inst_mult_11_609 ;
wire Xd_0__inst_mult_11_610 ;
wire Xd_0__inst_mult_11_614 ;
wire Xd_0__inst_mult_11_615 ;
wire Xd_0__inst_mult_10_609 ;
wire Xd_0__inst_mult_10_610 ;
wire Xd_0__inst_mult_10_614 ;
wire Xd_0__inst_mult_10_615 ;
wire Xd_0__inst_mult_5_609 ;
wire Xd_0__inst_mult_5_610 ;
wire Xd_0__inst_mult_5_614 ;
wire Xd_0__inst_mult_5_615 ;
wire Xd_0__inst_mult_4_609 ;
wire Xd_0__inst_mult_4_610 ;
wire Xd_0__inst_mult_4_614 ;
wire Xd_0__inst_mult_4_615 ;
wire Xd_0__inst_mult_7_609 ;
wire Xd_0__inst_mult_7_610 ;
wire Xd_0__inst_mult_7_614 ;
wire Xd_0__inst_mult_7_615 ;
wire Xd_0__inst_mult_6_609 ;
wire Xd_0__inst_mult_6_610 ;
wire Xd_0__inst_mult_6_614 ;
wire Xd_0__inst_mult_6_615 ;
wire Xd_0__inst_mult_1_609 ;
wire Xd_0__inst_mult_1_610 ;
wire Xd_0__inst_mult_1_614 ;
wire Xd_0__inst_mult_1_615 ;
wire Xd_0__inst_mult_0_609 ;
wire Xd_0__inst_mult_0_610 ;
wire Xd_0__inst_mult_0_614 ;
wire Xd_0__inst_mult_0_615 ;
wire Xd_0__inst_mult_3_609 ;
wire Xd_0__inst_mult_3_610 ;
wire Xd_0__inst_mult_3_614 ;
wire Xd_0__inst_mult_3_615 ;
wire Xd_0__inst_mult_2_654 ;
wire Xd_0__inst_mult_2_655 ;
wire Xd_0__inst_mult_2_659 ;
wire Xd_0__inst_mult_2_660 ;
wire Xd_0__inst_mult_29_629 ;
wire Xd_0__inst_mult_29_630 ;
wire Xd_0__inst_mult_29_634 ;
wire Xd_0__inst_mult_29_635 ;
wire Xd_0__inst_mult_28_619 ;
wire Xd_0__inst_mult_28_620 ;
wire Xd_0__inst_mult_28_624 ;
wire Xd_0__inst_mult_28_625 ;
wire Xd_0__inst_mult_31_619 ;
wire Xd_0__inst_mult_31_620 ;
wire Xd_0__inst_mult_31_624 ;
wire Xd_0__inst_mult_31_625 ;
wire Xd_0__inst_mult_30_619 ;
wire Xd_0__inst_mult_30_620 ;
wire Xd_0__inst_mult_30_624 ;
wire Xd_0__inst_mult_30_625 ;
wire Xd_0__inst_mult_25_644 ;
wire Xd_0__inst_mult_25_645 ;
wire Xd_0__inst_mult_25_649 ;
wire Xd_0__inst_mult_25_650 ;
wire Xd_0__inst_mult_27_644 ;
wire Xd_0__inst_mult_27_645 ;
wire Xd_0__inst_mult_27_649 ;
wire Xd_0__inst_mult_27_650 ;
wire Xd_0__inst_mult_21_629 ;
wire Xd_0__inst_mult_21_630 ;
wire Xd_0__inst_mult_21_634 ;
wire Xd_0__inst_mult_21_635 ;
wire Xd_0__inst_mult_20_629 ;
wire Xd_0__inst_mult_20_630 ;
wire Xd_0__inst_mult_20_634 ;
wire Xd_0__inst_mult_20_635 ;
wire Xd_0__inst_mult_23_629 ;
wire Xd_0__inst_mult_23_630 ;
wire Xd_0__inst_mult_23_634 ;
wire Xd_0__inst_mult_23_635 ;
wire Xd_0__inst_mult_22_629 ;
wire Xd_0__inst_mult_22_630 ;
wire Xd_0__inst_mult_22_634 ;
wire Xd_0__inst_mult_22_635 ;
wire Xd_0__inst_mult_17_629 ;
wire Xd_0__inst_mult_17_630 ;
wire Xd_0__inst_mult_17_634 ;
wire Xd_0__inst_mult_17_635 ;
wire Xd_0__inst_mult_16_629 ;
wire Xd_0__inst_mult_16_630 ;
wire Xd_0__inst_mult_16_634 ;
wire Xd_0__inst_mult_16_635 ;
wire Xd_0__inst_mult_19_629 ;
wire Xd_0__inst_mult_19_630 ;
wire Xd_0__inst_mult_19_634 ;
wire Xd_0__inst_mult_19_635 ;
wire Xd_0__inst_mult_18_604 ;
wire Xd_0__inst_mult_18_605 ;
wire Xd_0__inst_mult_18_609 ;
wire Xd_0__inst_mult_18_610 ;
wire Xd_0__inst_mult_18_614 ;
wire Xd_0__inst_mult_18_615 ;
wire Xd_0__inst_mult_13_619 ;
wire Xd_0__inst_mult_13_620 ;
wire Xd_0__inst_mult_13_624 ;
wire Xd_0__inst_mult_13_625 ;
wire Xd_0__inst_mult_12_604 ;
wire Xd_0__inst_mult_12_605 ;
wire Xd_0__inst_mult_12_609 ;
wire Xd_0__inst_mult_12_610 ;
wire Xd_0__inst_mult_12_614 ;
wire Xd_0__inst_mult_12_615 ;
wire Xd_0__inst_mult_15_604 ;
wire Xd_0__inst_mult_15_605 ;
wire Xd_0__inst_mult_15_609 ;
wire Xd_0__inst_mult_15_610 ;
wire Xd_0__inst_mult_15_614 ;
wire Xd_0__inst_mult_15_615 ;
wire Xd_0__inst_mult_14_604 ;
wire Xd_0__inst_mult_14_605 ;
wire Xd_0__inst_mult_14_609 ;
wire Xd_0__inst_mult_14_610 ;
wire Xd_0__inst_mult_14_614 ;
wire Xd_0__inst_mult_14_615 ;
wire Xd_0__inst_mult_9_619 ;
wire Xd_0__inst_mult_9_620 ;
wire Xd_0__inst_mult_9_624 ;
wire Xd_0__inst_mult_9_625 ;
wire Xd_0__inst_mult_8_619 ;
wire Xd_0__inst_mult_8_620 ;
wire Xd_0__inst_mult_8_624 ;
wire Xd_0__inst_mult_8_625 ;
wire Xd_0__inst_mult_11_619 ;
wire Xd_0__inst_mult_11_620 ;
wire Xd_0__inst_mult_11_624 ;
wire Xd_0__inst_mult_11_625 ;
wire Xd_0__inst_mult_10_619 ;
wire Xd_0__inst_mult_10_620 ;
wire Xd_0__inst_mult_10_624 ;
wire Xd_0__inst_mult_10_625 ;
wire Xd_0__inst_mult_5_619 ;
wire Xd_0__inst_mult_5_620 ;
wire Xd_0__inst_mult_5_624 ;
wire Xd_0__inst_mult_5_625 ;
wire Xd_0__inst_mult_4_619 ;
wire Xd_0__inst_mult_4_620 ;
wire Xd_0__inst_mult_4_624 ;
wire Xd_0__inst_mult_4_625 ;
wire Xd_0__inst_mult_7_619 ;
wire Xd_0__inst_mult_7_620 ;
wire Xd_0__inst_mult_7_624 ;
wire Xd_0__inst_mult_7_625 ;
wire Xd_0__inst_mult_6_619 ;
wire Xd_0__inst_mult_6_620 ;
wire Xd_0__inst_mult_6_624 ;
wire Xd_0__inst_mult_6_625 ;
wire Xd_0__inst_mult_1_619 ;
wire Xd_0__inst_mult_1_620 ;
wire Xd_0__inst_mult_1_624 ;
wire Xd_0__inst_mult_1_625 ;
wire Xd_0__inst_mult_0_619 ;
wire Xd_0__inst_mult_0_620 ;
wire Xd_0__inst_mult_0_624 ;
wire Xd_0__inst_mult_0_625 ;
wire Xd_0__inst_mult_3_619 ;
wire Xd_0__inst_mult_3_620 ;
wire Xd_0__inst_mult_3_624 ;
wire Xd_0__inst_mult_3_625 ;
wire Xd_0__inst_mult_2_664 ;
wire Xd_0__inst_mult_2_665 ;
wire Xd_0__inst_mult_2_669 ;
wire Xd_0__inst_mult_2_670 ;
wire Xd_0__inst_mult_29_639 ;
wire Xd_0__inst_mult_29_640 ;
wire Xd_0__inst_mult_29_644 ;
wire Xd_0__inst_mult_29_645 ;
wire Xd_0__inst_mult_28_629 ;
wire Xd_0__inst_mult_28_630 ;
wire Xd_0__inst_mult_28_634 ;
wire Xd_0__inst_mult_28_635 ;
wire Xd_0__inst_mult_31_629 ;
wire Xd_0__inst_mult_31_630 ;
wire Xd_0__inst_mult_31_634 ;
wire Xd_0__inst_mult_31_635 ;
wire Xd_0__inst_mult_30_629 ;
wire Xd_0__inst_mult_30_630 ;
wire Xd_0__inst_mult_30_634 ;
wire Xd_0__inst_mult_30_635 ;
wire Xd_0__inst_mult_25_654 ;
wire Xd_0__inst_mult_25_655 ;
wire Xd_0__inst_mult_25_659 ;
wire Xd_0__inst_mult_25_660 ;
wire Xd_0__inst_mult_27_654 ;
wire Xd_0__inst_mult_27_655 ;
wire Xd_0__inst_mult_27_659 ;
wire Xd_0__inst_mult_27_660 ;
wire Xd_0__inst_mult_21_639 ;
wire Xd_0__inst_mult_21_640 ;
wire Xd_0__inst_mult_21_644 ;
wire Xd_0__inst_mult_21_645 ;
wire Xd_0__inst_mult_20_639 ;
wire Xd_0__inst_mult_20_640 ;
wire Xd_0__inst_mult_20_644 ;
wire Xd_0__inst_mult_20_645 ;
wire Xd_0__inst_mult_23_639 ;
wire Xd_0__inst_mult_23_640 ;
wire Xd_0__inst_mult_23_644 ;
wire Xd_0__inst_mult_23_645 ;
wire Xd_0__inst_mult_22_639 ;
wire Xd_0__inst_mult_22_640 ;
wire Xd_0__inst_mult_22_644 ;
wire Xd_0__inst_mult_22_645 ;
wire Xd_0__inst_mult_17_639 ;
wire Xd_0__inst_mult_17_640 ;
wire Xd_0__inst_mult_17_644 ;
wire Xd_0__inst_mult_17_645 ;
wire Xd_0__inst_mult_16_639 ;
wire Xd_0__inst_mult_16_640 ;
wire Xd_0__inst_mult_16_644 ;
wire Xd_0__inst_mult_16_645 ;
wire Xd_0__inst_mult_19_639 ;
wire Xd_0__inst_mult_19_640 ;
wire Xd_0__inst_mult_19_644 ;
wire Xd_0__inst_mult_19_645 ;
wire Xd_0__inst_mult_18_619 ;
wire Xd_0__inst_mult_18_624 ;
wire Xd_0__inst_mult_18_625 ;
wire Xd_0__inst_mult_18_629 ;
wire Xd_0__inst_mult_18_630 ;
wire Xd_0__inst_mult_13_629 ;
wire Xd_0__inst_mult_13_630 ;
wire Xd_0__inst_mult_13_634 ;
wire Xd_0__inst_mult_13_635 ;
wire Xd_0__inst_mult_12_619 ;
wire Xd_0__inst_mult_12_624 ;
wire Xd_0__inst_mult_12_625 ;
wire Xd_0__inst_mult_12_629 ;
wire Xd_0__inst_mult_12_630 ;
wire Xd_0__inst_mult_15_619 ;
wire Xd_0__inst_mult_15_624 ;
wire Xd_0__inst_mult_15_625 ;
wire Xd_0__inst_mult_15_629 ;
wire Xd_0__inst_mult_15_630 ;
wire Xd_0__inst_mult_14_619 ;
wire Xd_0__inst_mult_14_75_sumout ;
wire Xd_0__inst_mult_14_76 ;
wire Xd_0__inst_mult_14_624 ;
wire Xd_0__inst_mult_14_625 ;
wire Xd_0__inst_mult_14_629 ;
wire Xd_0__inst_mult_14_630 ;
wire Xd_0__inst_mult_9_629 ;
wire Xd_0__inst_mult_9_630 ;
wire Xd_0__inst_mult_9_634 ;
wire Xd_0__inst_mult_9_635 ;
wire Xd_0__inst_mult_8_629 ;
wire Xd_0__inst_mult_8_630 ;
wire Xd_0__inst_mult_8_634 ;
wire Xd_0__inst_mult_8_635 ;
wire Xd_0__inst_mult_11_629 ;
wire Xd_0__inst_mult_11_630 ;
wire Xd_0__inst_mult_11_634 ;
wire Xd_0__inst_mult_11_635 ;
wire Xd_0__inst_mult_10_629 ;
wire Xd_0__inst_mult_10_630 ;
wire Xd_0__inst_mult_10_634 ;
wire Xd_0__inst_mult_10_635 ;
wire Xd_0__inst_mult_5_629 ;
wire Xd_0__inst_mult_5_630 ;
wire Xd_0__inst_mult_5_634 ;
wire Xd_0__inst_mult_5_635 ;
wire Xd_0__inst_mult_4_629 ;
wire Xd_0__inst_mult_4_630 ;
wire Xd_0__inst_mult_4_634 ;
wire Xd_0__inst_mult_4_635 ;
wire Xd_0__inst_mult_7_629 ;
wire Xd_0__inst_mult_7_630 ;
wire Xd_0__inst_mult_7_634 ;
wire Xd_0__inst_mult_7_635 ;
wire Xd_0__inst_mult_6_629 ;
wire Xd_0__inst_mult_6_630 ;
wire Xd_0__inst_mult_6_634 ;
wire Xd_0__inst_mult_6_635 ;
wire Xd_0__inst_mult_1_629 ;
wire Xd_0__inst_mult_1_630 ;
wire Xd_0__inst_mult_1_634 ;
wire Xd_0__inst_mult_1_635 ;
wire Xd_0__inst_mult_0_629 ;
wire Xd_0__inst_mult_0_630 ;
wire Xd_0__inst_mult_0_634 ;
wire Xd_0__inst_mult_0_635 ;
wire Xd_0__inst_mult_3_629 ;
wire Xd_0__inst_mult_3_630 ;
wire Xd_0__inst_mult_3_634 ;
wire Xd_0__inst_mult_3_635 ;
wire Xd_0__inst_mult_2_674 ;
wire Xd_0__inst_mult_2_675 ;
wire Xd_0__inst_mult_2_679 ;
wire Xd_0__inst_mult_2_680 ;
wire Xd_0__inst_mult_29_649 ;
wire Xd_0__inst_mult_29_650 ;
wire Xd_0__inst_mult_29_654 ;
wire Xd_0__inst_mult_29_655 ;
wire Xd_0__inst_mult_28_639 ;
wire Xd_0__inst_mult_28_640 ;
wire Xd_0__inst_mult_28_644 ;
wire Xd_0__inst_mult_28_645 ;
wire Xd_0__inst_mult_31_639 ;
wire Xd_0__inst_mult_31_640 ;
wire Xd_0__inst_mult_31_644 ;
wire Xd_0__inst_mult_31_645 ;
wire Xd_0__inst_mult_30_639 ;
wire Xd_0__inst_mult_30_640 ;
wire Xd_0__inst_mult_30_644 ;
wire Xd_0__inst_mult_30_645 ;
wire Xd_0__inst_mult_25_664 ;
wire Xd_0__inst_mult_25_665 ;
wire Xd_0__inst_mult_25_669 ;
wire Xd_0__inst_mult_25_670 ;
wire Xd_0__inst_mult_27_664 ;
wire Xd_0__inst_mult_27_665 ;
wire Xd_0__inst_mult_27_669 ;
wire Xd_0__inst_mult_27_670 ;
wire Xd_0__inst_mult_21_649 ;
wire Xd_0__inst_mult_21_650 ;
wire Xd_0__inst_mult_21_654 ;
wire Xd_0__inst_mult_21_655 ;
wire Xd_0__inst_mult_20_649 ;
wire Xd_0__inst_mult_20_650 ;
wire Xd_0__inst_mult_20_654 ;
wire Xd_0__inst_mult_20_655 ;
wire Xd_0__inst_mult_23_649 ;
wire Xd_0__inst_mult_23_650 ;
wire Xd_0__inst_mult_23_654 ;
wire Xd_0__inst_mult_23_655 ;
wire Xd_0__inst_mult_22_649 ;
wire Xd_0__inst_mult_22_650 ;
wire Xd_0__inst_mult_22_654 ;
wire Xd_0__inst_mult_22_655 ;
wire Xd_0__inst_mult_17_649 ;
wire Xd_0__inst_mult_17_650 ;
wire Xd_0__inst_mult_17_654 ;
wire Xd_0__inst_mult_17_655 ;
wire Xd_0__inst_mult_16_649 ;
wire Xd_0__inst_mult_16_650 ;
wire Xd_0__inst_mult_16_654 ;
wire Xd_0__inst_mult_16_655 ;
wire Xd_0__inst_mult_19_649 ;
wire Xd_0__inst_mult_19_650 ;
wire Xd_0__inst_mult_19_654 ;
wire Xd_0__inst_mult_19_655 ;
wire Xd_0__inst_mult_18_634 ;
wire Xd_0__inst_mult_18_635 ;
wire Xd_0__inst_mult_18_639 ;
wire Xd_0__inst_mult_18_640 ;
wire Xd_0__inst_mult_13_639 ;
wire Xd_0__inst_mult_13_640 ;
wire Xd_0__inst_mult_13_644 ;
wire Xd_0__inst_mult_13_645 ;
wire Xd_0__inst_mult_12_634 ;
wire Xd_0__inst_mult_12_635 ;
wire Xd_0__inst_mult_12_639 ;
wire Xd_0__inst_mult_12_640 ;
wire Xd_0__inst_mult_15_634 ;
wire Xd_0__inst_mult_15_635 ;
wire Xd_0__inst_mult_15_639 ;
wire Xd_0__inst_mult_15_640 ;
wire Xd_0__inst_mult_14_634 ;
wire Xd_0__inst_mult_14_635 ;
wire Xd_0__inst_mult_14_639 ;
wire Xd_0__inst_mult_14_640 ;
wire Xd_0__inst_mult_9_639 ;
wire Xd_0__inst_mult_9_640 ;
wire Xd_0__inst_mult_9_644 ;
wire Xd_0__inst_mult_9_645 ;
wire Xd_0__inst_mult_8_639 ;
wire Xd_0__inst_mult_8_640 ;
wire Xd_0__inst_mult_8_644 ;
wire Xd_0__inst_mult_8_645 ;
wire Xd_0__inst_mult_11_639 ;
wire Xd_0__inst_mult_11_640 ;
wire Xd_0__inst_mult_11_644 ;
wire Xd_0__inst_mult_11_645 ;
wire Xd_0__inst_mult_10_639 ;
wire Xd_0__inst_mult_10_640 ;
wire Xd_0__inst_mult_10_644 ;
wire Xd_0__inst_mult_10_645 ;
wire Xd_0__inst_mult_5_639 ;
wire Xd_0__inst_mult_5_640 ;
wire Xd_0__inst_mult_5_644 ;
wire Xd_0__inst_mult_5_645 ;
wire Xd_0__inst_mult_4_639 ;
wire Xd_0__inst_mult_4_640 ;
wire Xd_0__inst_mult_4_644 ;
wire Xd_0__inst_mult_4_645 ;
wire Xd_0__inst_mult_7_639 ;
wire Xd_0__inst_mult_7_640 ;
wire Xd_0__inst_mult_7_644 ;
wire Xd_0__inst_mult_7_645 ;
wire Xd_0__inst_mult_6_639 ;
wire Xd_0__inst_mult_6_640 ;
wire Xd_0__inst_mult_6_644 ;
wire Xd_0__inst_mult_6_645 ;
wire Xd_0__inst_mult_1_639 ;
wire Xd_0__inst_mult_1_640 ;
wire Xd_0__inst_mult_1_644 ;
wire Xd_0__inst_mult_1_645 ;
wire Xd_0__inst_mult_0_639 ;
wire Xd_0__inst_mult_0_640 ;
wire Xd_0__inst_mult_0_644 ;
wire Xd_0__inst_mult_0_645 ;
wire Xd_0__inst_mult_3_639 ;
wire Xd_0__inst_mult_3_640 ;
wire Xd_0__inst_mult_3_644 ;
wire Xd_0__inst_mult_3_645 ;
wire Xd_0__inst_mult_2_684 ;
wire Xd_0__inst_mult_2_685 ;
wire Xd_0__inst_mult_2_689 ;
wire Xd_0__inst_mult_2_690 ;
wire Xd_0__inst_mult_29_659 ;
wire Xd_0__inst_mult_29_660 ;
wire Xd_0__inst_mult_29_664 ;
wire Xd_0__inst_mult_29_665 ;
wire Xd_0__inst_mult_28_649 ;
wire Xd_0__inst_mult_28_650 ;
wire Xd_0__inst_mult_28_654 ;
wire Xd_0__inst_mult_28_655 ;
wire Xd_0__inst_mult_31_649 ;
wire Xd_0__inst_mult_31_650 ;
wire Xd_0__inst_mult_31_654 ;
wire Xd_0__inst_mult_31_655 ;
wire Xd_0__inst_mult_30_649 ;
wire Xd_0__inst_mult_30_650 ;
wire Xd_0__inst_mult_30_654 ;
wire Xd_0__inst_mult_30_655 ;
wire Xd_0__inst_mult_25_674 ;
wire Xd_0__inst_mult_25_675 ;
wire Xd_0__inst_mult_25_679 ;
wire Xd_0__inst_mult_25_680 ;
wire Xd_0__inst_mult_27_674 ;
wire Xd_0__inst_mult_27_675 ;
wire Xd_0__inst_mult_27_679 ;
wire Xd_0__inst_mult_27_680 ;
wire Xd_0__inst_mult_21_659 ;
wire Xd_0__inst_mult_21_660 ;
wire Xd_0__inst_mult_21_664 ;
wire Xd_0__inst_mult_21_665 ;
wire Xd_0__inst_mult_20_659 ;
wire Xd_0__inst_mult_20_660 ;
wire Xd_0__inst_mult_20_664 ;
wire Xd_0__inst_mult_20_665 ;
wire Xd_0__inst_mult_23_659 ;
wire Xd_0__inst_mult_23_660 ;
wire Xd_0__inst_mult_23_664 ;
wire Xd_0__inst_mult_23_665 ;
wire Xd_0__inst_mult_22_659 ;
wire Xd_0__inst_mult_22_660 ;
wire Xd_0__inst_mult_22_664 ;
wire Xd_0__inst_mult_22_665 ;
wire Xd_0__inst_mult_17_659 ;
wire Xd_0__inst_mult_17_660 ;
wire Xd_0__inst_mult_17_664 ;
wire Xd_0__inst_mult_17_665 ;
wire Xd_0__inst_mult_16_659 ;
wire Xd_0__inst_mult_16_660 ;
wire Xd_0__inst_mult_16_664 ;
wire Xd_0__inst_mult_16_665 ;
wire Xd_0__inst_mult_19_659 ;
wire Xd_0__inst_mult_19_660 ;
wire Xd_0__inst_mult_19_664 ;
wire Xd_0__inst_mult_19_665 ;
wire Xd_0__inst_mult_18_644 ;
wire Xd_0__inst_mult_18_645 ;
wire Xd_0__inst_mult_18_649 ;
wire Xd_0__inst_mult_18_650 ;
wire Xd_0__inst_mult_13_649 ;
wire Xd_0__inst_mult_13_650 ;
wire Xd_0__inst_mult_13_654 ;
wire Xd_0__inst_mult_13_655 ;
wire Xd_0__inst_mult_12_644 ;
wire Xd_0__inst_mult_12_645 ;
wire Xd_0__inst_mult_12_649 ;
wire Xd_0__inst_mult_12_650 ;
wire Xd_0__inst_mult_15_644 ;
wire Xd_0__inst_mult_15_645 ;
wire Xd_0__inst_mult_15_649 ;
wire Xd_0__inst_mult_15_650 ;
wire Xd_0__inst_mult_14_644 ;
wire Xd_0__inst_mult_14_645 ;
wire Xd_0__inst_mult_14_649 ;
wire Xd_0__inst_mult_14_650 ;
wire Xd_0__inst_mult_9_649 ;
wire Xd_0__inst_mult_9_650 ;
wire Xd_0__inst_mult_9_654 ;
wire Xd_0__inst_mult_9_655 ;
wire Xd_0__inst_mult_8_649 ;
wire Xd_0__inst_mult_8_650 ;
wire Xd_0__inst_mult_8_654 ;
wire Xd_0__inst_mult_8_655 ;
wire Xd_0__inst_mult_11_649 ;
wire Xd_0__inst_mult_11_650 ;
wire Xd_0__inst_mult_11_654 ;
wire Xd_0__inst_mult_11_655 ;
wire Xd_0__inst_mult_10_649 ;
wire Xd_0__inst_mult_10_650 ;
wire Xd_0__inst_mult_10_654 ;
wire Xd_0__inst_mult_10_655 ;
wire Xd_0__inst_mult_5_649 ;
wire Xd_0__inst_mult_5_650 ;
wire Xd_0__inst_mult_5_654 ;
wire Xd_0__inst_mult_5_655 ;
wire Xd_0__inst_mult_4_649 ;
wire Xd_0__inst_mult_4_650 ;
wire Xd_0__inst_mult_4_654 ;
wire Xd_0__inst_mult_4_655 ;
wire Xd_0__inst_mult_7_649 ;
wire Xd_0__inst_mult_7_650 ;
wire Xd_0__inst_mult_7_654 ;
wire Xd_0__inst_mult_7_655 ;
wire Xd_0__inst_mult_6_649 ;
wire Xd_0__inst_mult_6_650 ;
wire Xd_0__inst_mult_6_654 ;
wire Xd_0__inst_mult_6_655 ;
wire Xd_0__inst_mult_1_649 ;
wire Xd_0__inst_mult_1_650 ;
wire Xd_0__inst_mult_1_654 ;
wire Xd_0__inst_mult_1_655 ;
wire Xd_0__inst_mult_0_649 ;
wire Xd_0__inst_mult_0_650 ;
wire Xd_0__inst_mult_0_654 ;
wire Xd_0__inst_mult_0_655 ;
wire Xd_0__inst_mult_3_649 ;
wire Xd_0__inst_mult_3_650 ;
wire Xd_0__inst_mult_3_654 ;
wire Xd_0__inst_mult_3_655 ;
wire Xd_0__inst_mult_2_694 ;
wire Xd_0__inst_mult_2_695 ;
wire Xd_0__inst_mult_2_699 ;
wire Xd_0__inst_mult_2_700 ;
wire Xd_0__inst_mult_29_669 ;
wire Xd_0__inst_mult_29_674 ;
wire Xd_0__inst_mult_29_675 ;
wire Xd_0__inst_mult_28_659 ;
wire Xd_0__inst_mult_28_664 ;
wire Xd_0__inst_mult_28_665 ;
wire Xd_0__inst_mult_31_659 ;
wire Xd_0__inst_mult_31_664 ;
wire Xd_0__inst_mult_31_665 ;
wire Xd_0__inst_mult_30_659 ;
wire Xd_0__inst_mult_30_664 ;
wire Xd_0__inst_mult_30_665 ;
wire Xd_0__inst_mult_25_684 ;
wire Xd_0__inst_mult_25_689 ;
wire Xd_0__inst_mult_25_690 ;
wire Xd_0__inst_mult_27_684 ;
wire Xd_0__inst_mult_27_689 ;
wire Xd_0__inst_mult_27_690 ;
wire Xd_0__inst_mult_21_669 ;
wire Xd_0__inst_mult_21_674 ;
wire Xd_0__inst_mult_21_675 ;
wire Xd_0__inst_mult_20_669 ;
wire Xd_0__inst_mult_20_674 ;
wire Xd_0__inst_mult_20_675 ;
wire Xd_0__inst_mult_23_669 ;
wire Xd_0__inst_mult_23_674 ;
wire Xd_0__inst_mult_23_675 ;
wire Xd_0__inst_mult_22_669 ;
wire Xd_0__inst_mult_22_674 ;
wire Xd_0__inst_mult_22_675 ;
wire Xd_0__inst_mult_17_669 ;
wire Xd_0__inst_mult_17_674 ;
wire Xd_0__inst_mult_17_675 ;
wire Xd_0__inst_mult_16_669 ;
wire Xd_0__inst_mult_16_674 ;
wire Xd_0__inst_mult_16_675 ;
wire Xd_0__inst_mult_19_669 ;
wire Xd_0__inst_mult_19_674 ;
wire Xd_0__inst_mult_19_675 ;
wire Xd_0__inst_mult_18_654 ;
wire Xd_0__inst_mult_18_659 ;
wire Xd_0__inst_mult_18_660 ;
wire Xd_0__inst_mult_13_659 ;
wire Xd_0__inst_mult_13_664 ;
wire Xd_0__inst_mult_13_665 ;
wire Xd_0__inst_mult_12_654 ;
wire Xd_0__inst_mult_12_659 ;
wire Xd_0__inst_mult_12_660 ;
wire Xd_0__inst_mult_15_654 ;
wire Xd_0__inst_mult_15_659 ;
wire Xd_0__inst_mult_15_660 ;
wire Xd_0__inst_mult_14_654 ;
wire Xd_0__inst_mult_14_659 ;
wire Xd_0__inst_mult_14_660 ;
wire Xd_0__inst_mult_9_659 ;
wire Xd_0__inst_mult_9_664 ;
wire Xd_0__inst_mult_9_665 ;
wire Xd_0__inst_mult_8_659 ;
wire Xd_0__inst_mult_8_664 ;
wire Xd_0__inst_mult_8_665 ;
wire Xd_0__inst_mult_11_659 ;
wire Xd_0__inst_mult_11_664 ;
wire Xd_0__inst_mult_11_665 ;
wire Xd_0__inst_mult_10_659 ;
wire Xd_0__inst_mult_10_664 ;
wire Xd_0__inst_mult_10_665 ;
wire Xd_0__inst_mult_5_659 ;
wire Xd_0__inst_mult_5_664 ;
wire Xd_0__inst_mult_5_665 ;
wire Xd_0__inst_mult_4_659 ;
wire Xd_0__inst_mult_4_664 ;
wire Xd_0__inst_mult_4_665 ;
wire Xd_0__inst_mult_7_659 ;
wire Xd_0__inst_mult_7_664 ;
wire Xd_0__inst_mult_7_665 ;
wire Xd_0__inst_mult_6_659 ;
wire Xd_0__inst_mult_6_664 ;
wire Xd_0__inst_mult_6_665 ;
wire Xd_0__inst_mult_1_659 ;
wire Xd_0__inst_mult_1_664 ;
wire Xd_0__inst_mult_1_665 ;
wire Xd_0__inst_mult_0_659 ;
wire Xd_0__inst_mult_0_664 ;
wire Xd_0__inst_mult_0_665 ;
wire Xd_0__inst_mult_3_659 ;
wire Xd_0__inst_mult_3_664 ;
wire Xd_0__inst_mult_3_665 ;
wire Xd_0__inst_mult_2_704 ;
wire Xd_0__inst_mult_2_709 ;
wire Xd_0__inst_mult_2_710 ;
wire Xd_0__inst_mult_29_679 ;
wire Xd_0__inst_mult_29_680 ;
wire Xd_0__inst_mult_29_80_sumout ;
wire Xd_0__inst_mult_29_81 ;
wire Xd_0__inst_mult_28_669 ;
wire Xd_0__inst_mult_28_670 ;
wire Xd_0__inst_mult_28_80_sumout ;
wire Xd_0__inst_mult_28_81 ;
wire Xd_0__inst_mult_31_669 ;
wire Xd_0__inst_mult_31_670 ;
wire Xd_0__inst_mult_31_80_sumout ;
wire Xd_0__inst_mult_31_81 ;
wire Xd_0__inst_mult_30_669 ;
wire Xd_0__inst_mult_30_670 ;
wire Xd_0__inst_mult_25_694 ;
wire Xd_0__inst_mult_25_695 ;
wire Xd_0__inst_mult_27_694 ;
wire Xd_0__inst_mult_27_695 ;
wire Xd_0__inst_mult_21_679 ;
wire Xd_0__inst_mult_21_680 ;
wire Xd_0__inst_mult_21_80_sumout ;
wire Xd_0__inst_mult_21_81 ;
wire Xd_0__inst_mult_20_679 ;
wire Xd_0__inst_mult_20_680 ;
wire Xd_0__inst_mult_23_679 ;
wire Xd_0__inst_mult_23_680 ;
wire Xd_0__inst_mult_22_679 ;
wire Xd_0__inst_mult_22_680 ;
wire Xd_0__inst_mult_22_80_sumout ;
wire Xd_0__inst_mult_22_81 ;
wire Xd_0__inst_mult_17_679 ;
wire Xd_0__inst_mult_17_680 ;
wire Xd_0__inst_mult_17_80_sumout ;
wire Xd_0__inst_mult_17_81 ;
wire Xd_0__inst_mult_16_679 ;
wire Xd_0__inst_mult_16_680 ;
wire Xd_0__inst_mult_16_75_sumout ;
wire Xd_0__inst_mult_16_76 ;
wire Xd_0__inst_mult_19_679 ;
wire Xd_0__inst_mult_19_680 ;
wire Xd_0__inst_mult_19_75_sumout ;
wire Xd_0__inst_mult_19_76 ;
wire Xd_0__inst_mult_18_664 ;
wire Xd_0__inst_mult_18_665 ;
wire Xd_0__inst_mult_18_75_sumout ;
wire Xd_0__inst_mult_18_76 ;
wire Xd_0__inst_mult_13_669 ;
wire Xd_0__inst_mult_13_670 ;
wire Xd_0__inst_mult_13_75_sumout ;
wire Xd_0__inst_mult_13_76 ;
wire Xd_0__inst_mult_12_664 ;
wire Xd_0__inst_mult_12_665 ;
wire Xd_0__inst_mult_15_664 ;
wire Xd_0__inst_mult_15_665 ;
wire Xd_0__inst_mult_14_664 ;
wire Xd_0__inst_mult_14_665 ;
wire Xd_0__inst_mult_9_669 ;
wire Xd_0__inst_mult_9_670 ;
wire Xd_0__inst_mult_9_75_sumout ;
wire Xd_0__inst_mult_9_76 ;
wire Xd_0__inst_mult_8_669 ;
wire Xd_0__inst_mult_8_670 ;
wire Xd_0__inst_mult_11_669 ;
wire Xd_0__inst_mult_11_670 ;
wire Xd_0__inst_mult_10_669 ;
wire Xd_0__inst_mult_10_670 ;
wire Xd_0__inst_mult_5_669 ;
wire Xd_0__inst_mult_5_670 ;
wire Xd_0__inst_mult_4_669 ;
wire Xd_0__inst_mult_4_670 ;
wire Xd_0__inst_mult_7_669 ;
wire Xd_0__inst_mult_7_670 ;
wire Xd_0__inst_mult_6_669 ;
wire Xd_0__inst_mult_6_670 ;
wire Xd_0__inst_mult_1_669 ;
wire Xd_0__inst_mult_1_670 ;
wire Xd_0__inst_mult_0_669 ;
wire Xd_0__inst_mult_0_670 ;
wire Xd_0__inst_mult_3_669 ;
wire Xd_0__inst_mult_3_670 ;
wire Xd_0__inst_mult_2_714 ;
wire Xd_0__inst_mult_2_715 ;
wire Xd_0__inst_mult_29_684 ;
wire Xd_0__inst_mult_28_674 ;
wire Xd_0__inst_mult_31_674 ;
wire Xd_0__inst_mult_30_674 ;
wire Xd_0__inst_mult_25_699 ;
wire Xd_0__inst_mult_27_699 ;
wire Xd_0__inst_mult_21_684 ;
wire Xd_0__inst_mult_20_684 ;
wire Xd_0__inst_mult_23_684 ;
wire Xd_0__inst_mult_22_684 ;
wire Xd_0__inst_mult_17_684 ;
wire Xd_0__inst_mult_16_684 ;
wire Xd_0__inst_mult_16_80_sumout ;
wire Xd_0__inst_mult_16_81 ;
wire Xd_0__inst_mult_19_684 ;
wire Xd_0__inst_mult_19_80_sumout ;
wire Xd_0__inst_mult_19_81 ;
wire Xd_0__inst_mult_18_669 ;
wire Xd_0__inst_mult_18_80_sumout ;
wire Xd_0__inst_mult_18_81 ;
wire Xd_0__inst_mult_13_674 ;
wire Xd_0__inst_mult_13_80_sumout ;
wire Xd_0__inst_mult_13_81 ;
wire Xd_0__inst_mult_12_669 ;
wire Xd_0__inst_mult_15_669 ;
wire Xd_0__inst_mult_14_669 ;
wire Xd_0__inst_mult_14_80_sumout ;
wire Xd_0__inst_mult_14_81 ;
wire Xd_0__inst_mult_9_674 ;
wire Xd_0__inst_mult_9_80_sumout ;
wire Xd_0__inst_mult_9_81 ;
wire Xd_0__inst_mult_8_674 ;
wire Xd_0__inst_mult_11_674 ;
wire Xd_0__inst_mult_11_80_sumout ;
wire Xd_0__inst_mult_11_81 ;
wire Xd_0__inst_mult_10_674 ;
wire Xd_0__inst_mult_5_674 ;
wire Xd_0__inst_mult_4_674 ;
wire Xd_0__inst_mult_4_80_sumout ;
wire Xd_0__inst_mult_4_81 ;
wire Xd_0__inst_mult_7_674 ;
wire Xd_0__inst_mult_7_80_sumout ;
wire Xd_0__inst_mult_7_81 ;
wire Xd_0__inst_mult_6_674 ;
wire Xd_0__inst_mult_6_80_sumout ;
wire Xd_0__inst_mult_6_81 ;
wire Xd_0__inst_mult_1_674 ;
wire Xd_0__inst_mult_1_80_sumout ;
wire Xd_0__inst_mult_1_81 ;
wire Xd_0__inst_mult_0_674 ;
wire Xd_0__inst_mult_3_674 ;
wire Xd_0__inst_mult_2_719 ;
wire Xd_0__inst_mult_9_679 ;
wire Xd_0__inst_mult_9_680 ;
wire Xd_0__inst_mult_8_679 ;
wire Xd_0__inst_mult_8_680 ;
wire Xd_0__inst_mult_21_689 ;
wire Xd_0__inst_mult_21_690 ;
wire Xd_0__inst_mult_11_679 ;
wire Xd_0__inst_mult_11_680 ;
wire Xd_0__inst_mult_10_679 ;
wire Xd_0__inst_mult_10_680 ;
wire Xd_0__inst_mult_20_689 ;
wire Xd_0__inst_mult_20_690 ;
wire Xd_0__inst_mult_25_704 ;
wire Xd_0__inst_mult_25_705 ;
wire Xd_0__inst_mult_3_679 ;
wire Xd_0__inst_mult_3_680 ;
wire Xd_0__inst_mult_0_679 ;
wire Xd_0__inst_mult_0_680 ;
wire Xd_0__inst_mult_23_689 ;
wire Xd_0__inst_mult_23_690 ;
wire Xd_0__inst_mult_6_679 ;
wire Xd_0__inst_mult_6_680 ;
wire Xd_0__inst_mult_1_679 ;
wire Xd_0__inst_mult_1_680 ;
wire Xd_0__inst_mult_22_689 ;
wire Xd_0__inst_mult_22_690 ;
wire Xd_0__inst_mult_24_774 ;
wire Xd_0__inst_mult_24_775 ;
wire Xd_0__inst_mult_26_774 ;
wire Xd_0__inst_mult_26_775 ;
wire Xd_0__inst_mult_7_679 ;
wire Xd_0__inst_mult_7_680 ;
wire Xd_0__inst_mult_4_679 ;
wire Xd_0__inst_mult_4_680 ;
wire Xd_0__inst_mult_19_689 ;
wire Xd_0__inst_mult_19_690 ;
wire Xd_0__inst_mult_30_679 ;
wire Xd_0__inst_mult_30_680 ;
wire Xd_0__inst_mult_5_679 ;
wire Xd_0__inst_mult_5_680 ;
wire Xd_0__inst_mult_17_689 ;
wire Xd_0__inst_mult_17_690 ;
wire Xd_0__inst_mult_27_704 ;
wire Xd_0__inst_mult_27_705 ;
wire Xd_0__inst_mult_13_679 ;
wire Xd_0__inst_mult_13_680 ;
wire Xd_0__inst_mult_2_724 ;
wire Xd_0__inst_mult_2_725 ;
wire Xd_0__inst_mult_16_689 ;
wire Xd_0__inst_mult_16_690 ;
wire Xd_0__inst_mult_28_679 ;
wire Xd_0__inst_mult_28_680 ;
wire Xd_0__inst_mult_31_679 ;
wire Xd_0__inst_mult_31_680 ;
wire Xd_0__inst_mult_29_689 ;
wire Xd_0__inst_mult_29_690 ;
wire Xd_0__inst_mult_26_779 ;
wire Xd_0__inst_mult_26_780 ;
wire Xd_0__inst_mult_24_779 ;
wire Xd_0__inst_mult_24_780 ;
wire Xd_0__inst_mult_29_694 ;
wire Xd_0__inst_mult_29_695 ;
wire Xd_0__inst_mult_29_700 ;
wire Xd_0__inst_mult_28_684 ;
wire Xd_0__inst_mult_28_685 ;
wire Xd_0__inst_mult_28_690 ;
wire Xd_0__inst_mult_31_684 ;
wire Xd_0__inst_mult_31_685 ;
wire Xd_0__inst_mult_31_690 ;
wire Xd_0__inst_mult_30_684 ;
wire Xd_0__inst_mult_30_685 ;
wire Xd_0__inst_mult_30_690 ;
wire Xd_0__inst_mult_25_709 ;
wire Xd_0__inst_mult_25_710 ;
wire Xd_0__inst_mult_25_715 ;
wire Xd_0__inst_mult_24_784 ;
wire Xd_0__inst_mult_24_785 ;
wire Xd_0__inst_mult_24_790 ;
wire Xd_0__inst_mult_27_709 ;
wire Xd_0__inst_mult_27_710 ;
wire Xd_0__inst_mult_27_715 ;
wire Xd_0__inst_mult_26_784 ;
wire Xd_0__inst_mult_26_785 ;
wire Xd_0__inst_mult_26_790 ;
wire Xd_0__inst_mult_21_694 ;
wire Xd_0__inst_mult_21_695 ;
wire Xd_0__inst_mult_21_700 ;
wire Xd_0__inst_mult_20_694 ;
wire Xd_0__inst_mult_20_695 ;
wire Xd_0__inst_mult_20_700 ;
wire Xd_0__inst_mult_23_694 ;
wire Xd_0__inst_mult_23_695 ;
wire Xd_0__inst_mult_23_700 ;
wire Xd_0__inst_mult_22_694 ;
wire Xd_0__inst_mult_22_695 ;
wire Xd_0__inst_mult_22_700 ;
wire Xd_0__inst_mult_17_694 ;
wire Xd_0__inst_mult_17_695 ;
wire Xd_0__inst_mult_17_700 ;
wire Xd_0__inst_mult_16_694 ;
wire Xd_0__inst_mult_16_695 ;
wire Xd_0__inst_mult_16_700 ;
wire Xd_0__inst_mult_19_694 ;
wire Xd_0__inst_mult_19_695 ;
wire Xd_0__inst_mult_19_700 ;
wire Xd_0__inst_mult_18_674 ;
wire Xd_0__inst_mult_18_675 ;
wire Xd_0__inst_mult_18_680 ;
wire Xd_0__inst_mult_13_684 ;
wire Xd_0__inst_mult_13_685 ;
wire Xd_0__inst_mult_13_690 ;
wire Xd_0__inst_mult_12_674 ;
wire Xd_0__inst_mult_12_675 ;
wire Xd_0__inst_mult_12_680 ;
wire Xd_0__inst_mult_15_674 ;
wire Xd_0__inst_mult_15_675 ;
wire Xd_0__inst_mult_15_680 ;
wire Xd_0__inst_mult_14_674 ;
wire Xd_0__inst_mult_14_675 ;
wire Xd_0__inst_mult_14_680 ;
wire Xd_0__inst_mult_9_684 ;
wire Xd_0__inst_mult_9_685 ;
wire Xd_0__inst_mult_9_690 ;
wire Xd_0__inst_mult_8_684 ;
wire Xd_0__inst_mult_8_685 ;
wire Xd_0__inst_mult_8_690 ;
wire Xd_0__inst_mult_11_684 ;
wire Xd_0__inst_mult_11_685 ;
wire Xd_0__inst_mult_11_690 ;
wire Xd_0__inst_mult_10_684 ;
wire Xd_0__inst_mult_10_685 ;
wire Xd_0__inst_mult_10_690 ;
wire Xd_0__inst_mult_5_684 ;
wire Xd_0__inst_mult_5_685 ;
wire Xd_0__inst_mult_5_690 ;
wire Xd_0__inst_mult_4_684 ;
wire Xd_0__inst_mult_4_685 ;
wire Xd_0__inst_mult_4_690 ;
wire Xd_0__inst_mult_7_684 ;
wire Xd_0__inst_mult_7_685 ;
wire Xd_0__inst_mult_7_690 ;
wire Xd_0__inst_mult_6_684 ;
wire Xd_0__inst_mult_6_685 ;
wire Xd_0__inst_mult_6_690 ;
wire Xd_0__inst_mult_1_684 ;
wire Xd_0__inst_mult_1_685 ;
wire Xd_0__inst_mult_1_690 ;
wire Xd_0__inst_mult_0_684 ;
wire Xd_0__inst_mult_0_685 ;
wire Xd_0__inst_mult_0_690 ;
wire Xd_0__inst_mult_3_684 ;
wire Xd_0__inst_mult_3_685 ;
wire Xd_0__inst_mult_3_690 ;
wire Xd_0__inst_mult_2_729 ;
wire Xd_0__inst_mult_2_730 ;
wire Xd_0__inst_mult_2_735 ;
wire Xd_0__inst_mult_29_704 ;
wire Xd_0__inst_mult_29_705 ;
wire Xd_0__inst_mult_28_694 ;
wire Xd_0__inst_mult_28_695 ;
wire Xd_0__inst_mult_31_694 ;
wire Xd_0__inst_mult_31_695 ;
wire Xd_0__inst_mult_30_694 ;
wire Xd_0__inst_mult_30_695 ;
wire Xd_0__inst_mult_25_719 ;
wire Xd_0__inst_mult_25_720 ;
wire Xd_0__inst_mult_24_794 ;
wire Xd_0__inst_mult_24_795 ;
wire Xd_0__inst_mult_27_719 ;
wire Xd_0__inst_mult_27_720 ;
wire Xd_0__inst_mult_26_794 ;
wire Xd_0__inst_mult_26_795 ;
wire Xd_0__inst_mult_21_704 ;
wire Xd_0__inst_mult_21_705 ;
wire Xd_0__inst_mult_20_704 ;
wire Xd_0__inst_mult_20_705 ;
wire Xd_0__inst_mult_23_704 ;
wire Xd_0__inst_mult_23_705 ;
wire Xd_0__inst_mult_22_704 ;
wire Xd_0__inst_mult_22_705 ;
wire Xd_0__inst_mult_17_704 ;
wire Xd_0__inst_mult_17_705 ;
wire Xd_0__inst_mult_16_704 ;
wire Xd_0__inst_mult_16_705 ;
wire Xd_0__inst_mult_19_704 ;
wire Xd_0__inst_mult_19_705 ;
wire Xd_0__inst_mult_18_684 ;
wire Xd_0__inst_mult_18_685 ;
wire Xd_0__inst_mult_13_694 ;
wire Xd_0__inst_mult_13_695 ;
wire Xd_0__inst_mult_12_684 ;
wire Xd_0__inst_mult_12_685 ;
wire Xd_0__inst_mult_15_684 ;
wire Xd_0__inst_mult_15_685 ;
wire Xd_0__inst_mult_14_684 ;
wire Xd_0__inst_mult_14_685 ;
wire Xd_0__inst_mult_9_694 ;
wire Xd_0__inst_mult_9_695 ;
wire Xd_0__inst_mult_8_694 ;
wire Xd_0__inst_mult_8_695 ;
wire Xd_0__inst_mult_11_694 ;
wire Xd_0__inst_mult_11_695 ;
wire Xd_0__inst_mult_10_694 ;
wire Xd_0__inst_mult_10_695 ;
wire Xd_0__inst_mult_5_694 ;
wire Xd_0__inst_mult_5_695 ;
wire Xd_0__inst_mult_4_694 ;
wire Xd_0__inst_mult_4_695 ;
wire Xd_0__inst_mult_7_694 ;
wire Xd_0__inst_mult_7_695 ;
wire Xd_0__inst_mult_6_694 ;
wire Xd_0__inst_mult_6_695 ;
wire Xd_0__inst_mult_1_694 ;
wire Xd_0__inst_mult_1_695 ;
wire Xd_0__inst_mult_0_694 ;
wire Xd_0__inst_mult_0_695 ;
wire Xd_0__inst_mult_3_694 ;
wire Xd_0__inst_mult_3_695 ;
wire Xd_0__inst_mult_2_739 ;
wire Xd_0__inst_mult_2_740 ;
wire Xd_0__inst_mult_29_709 ;
wire Xd_0__inst_mult_29_710 ;
wire Xd_0__inst_mult_28_699 ;
wire Xd_0__inst_mult_28_700 ;
wire Xd_0__inst_mult_31_699 ;
wire Xd_0__inst_mult_31_700 ;
wire Xd_0__inst_mult_30_699 ;
wire Xd_0__inst_mult_30_700 ;
wire Xd_0__inst_mult_21_709 ;
wire Xd_0__inst_mult_21_710 ;
wire Xd_0__inst_mult_20_709 ;
wire Xd_0__inst_mult_20_710 ;
wire Xd_0__inst_mult_23_709 ;
wire Xd_0__inst_mult_23_710 ;
wire Xd_0__inst_mult_22_709 ;
wire Xd_0__inst_mult_22_710 ;
wire Xd_0__inst_mult_17_709 ;
wire Xd_0__inst_mult_17_710 ;
wire Xd_0__inst_mult_16_709 ;
wire Xd_0__inst_mult_16_710 ;
wire Xd_0__inst_mult_19_709 ;
wire Xd_0__inst_mult_19_710 ;
wire Xd_0__inst_mult_18_689 ;
wire Xd_0__inst_mult_18_690 ;
wire Xd_0__inst_mult_13_699 ;
wire Xd_0__inst_mult_13_700 ;
wire Xd_0__inst_mult_12_689 ;
wire Xd_0__inst_mult_12_690 ;
wire Xd_0__inst_mult_15_689 ;
wire Xd_0__inst_mult_15_690 ;
wire Xd_0__inst_mult_14_689 ;
wire Xd_0__inst_mult_14_690 ;
wire Xd_0__inst_mult_9_699 ;
wire Xd_0__inst_mult_9_700 ;
wire Xd_0__inst_mult_8_699 ;
wire Xd_0__inst_mult_8_700 ;
wire Xd_0__inst_mult_11_699 ;
wire Xd_0__inst_mult_11_700 ;
wire Xd_0__inst_mult_10_699 ;
wire Xd_0__inst_mult_10_700 ;
wire Xd_0__inst_mult_5_699 ;
wire Xd_0__inst_mult_5_700 ;
wire Xd_0__inst_mult_4_699 ;
wire Xd_0__inst_mult_4_700 ;
wire Xd_0__inst_mult_7_699 ;
wire Xd_0__inst_mult_7_700 ;
wire Xd_0__inst_mult_6_699 ;
wire Xd_0__inst_mult_6_700 ;
wire Xd_0__inst_mult_1_699 ;
wire Xd_0__inst_mult_1_700 ;
wire Xd_0__inst_mult_0_699 ;
wire Xd_0__inst_mult_0_700 ;
wire Xd_0__inst_mult_3_699 ;
wire Xd_0__inst_mult_3_700 ;
wire Xd_0__inst_mult_2_744 ;
wire Xd_0__inst_mult_2_745 ;
wire Xd_0__inst_mult_29_714 ;
wire Xd_0__inst_mult_29_715 ;
wire Xd_0__inst_mult_29_719 ;
wire Xd_0__inst_mult_29_720 ;
wire Xd_0__inst_mult_29_725 ;
wire Xd_0__inst_mult_28_704 ;
wire Xd_0__inst_mult_28_705 ;
wire Xd_0__inst_mult_28_709 ;
wire Xd_0__inst_mult_28_710 ;
wire Xd_0__inst_mult_28_715 ;
wire Xd_0__inst_mult_31_704 ;
wire Xd_0__inst_mult_31_705 ;
wire Xd_0__inst_mult_31_709 ;
wire Xd_0__inst_mult_31_710 ;
wire Xd_0__inst_mult_31_715 ;
wire Xd_0__inst_mult_30_704 ;
wire Xd_0__inst_mult_30_705 ;
wire Xd_0__inst_mult_30_709 ;
wire Xd_0__inst_mult_30_710 ;
wire Xd_0__inst_mult_30_715 ;
wire Xd_0__inst_mult_25_724 ;
wire Xd_0__inst_mult_25_725 ;
wire Xd_0__inst_mult_25_730 ;
wire Xd_0__inst_mult_24_799 ;
wire Xd_0__inst_mult_24_800 ;
wire Xd_0__inst_mult_24_805 ;
wire Xd_0__inst_mult_27_724 ;
wire Xd_0__inst_mult_27_725 ;
wire Xd_0__inst_mult_27_730 ;
wire Xd_0__inst_mult_26_799 ;
wire Xd_0__inst_mult_26_800 ;
wire Xd_0__inst_mult_26_805 ;
wire Xd_0__inst_mult_21_714 ;
wire Xd_0__inst_mult_21_715 ;
wire Xd_0__inst_mult_21_719 ;
wire Xd_0__inst_mult_21_720 ;
wire Xd_0__inst_mult_21_725 ;
wire Xd_0__inst_mult_20_714 ;
wire Xd_0__inst_mult_20_715 ;
wire Xd_0__inst_mult_20_719 ;
wire Xd_0__inst_mult_20_720 ;
wire Xd_0__inst_mult_20_725 ;
wire Xd_0__inst_mult_23_714 ;
wire Xd_0__inst_mult_23_715 ;
wire Xd_0__inst_mult_23_719 ;
wire Xd_0__inst_mult_23_720 ;
wire Xd_0__inst_mult_23_725 ;
wire Xd_0__inst_mult_22_714 ;
wire Xd_0__inst_mult_22_715 ;
wire Xd_0__inst_mult_22_719 ;
wire Xd_0__inst_mult_22_720 ;
wire Xd_0__inst_mult_22_725 ;
wire Xd_0__inst_mult_17_714 ;
wire Xd_0__inst_mult_17_715 ;
wire Xd_0__inst_mult_17_719 ;
wire Xd_0__inst_mult_17_720 ;
wire Xd_0__inst_mult_17_725 ;
wire Xd_0__inst_mult_16_714 ;
wire Xd_0__inst_mult_16_715 ;
wire Xd_0__inst_mult_16_719 ;
wire Xd_0__inst_mult_16_720 ;
wire Xd_0__inst_mult_16_725 ;
wire Xd_0__inst_mult_19_714 ;
wire Xd_0__inst_mult_19_715 ;
wire Xd_0__inst_mult_19_719 ;
wire Xd_0__inst_mult_19_720 ;
wire Xd_0__inst_mult_19_725 ;
wire Xd_0__inst_mult_18_694 ;
wire Xd_0__inst_mult_18_695 ;
wire Xd_0__inst_mult_18_699 ;
wire Xd_0__inst_mult_18_700 ;
wire Xd_0__inst_mult_18_705 ;
wire Xd_0__inst_mult_13_704 ;
wire Xd_0__inst_mult_13_705 ;
wire Xd_0__inst_mult_13_709 ;
wire Xd_0__inst_mult_13_710 ;
wire Xd_0__inst_mult_13_715 ;
wire Xd_0__inst_mult_12_694 ;
wire Xd_0__inst_mult_12_695 ;
wire Xd_0__inst_mult_12_699 ;
wire Xd_0__inst_mult_12_700 ;
wire Xd_0__inst_mult_12_705 ;
wire Xd_0__inst_mult_15_694 ;
wire Xd_0__inst_mult_15_695 ;
wire Xd_0__inst_mult_15_699 ;
wire Xd_0__inst_mult_15_700 ;
wire Xd_0__inst_mult_15_705 ;
wire Xd_0__inst_mult_14_694 ;
wire Xd_0__inst_mult_14_695 ;
wire Xd_0__inst_mult_14_699 ;
wire Xd_0__inst_mult_14_700 ;
wire Xd_0__inst_mult_14_705 ;
wire Xd_0__inst_mult_9_704 ;
wire Xd_0__inst_mult_9_705 ;
wire Xd_0__inst_mult_9_709 ;
wire Xd_0__inst_mult_9_710 ;
wire Xd_0__inst_mult_9_715 ;
wire Xd_0__inst_mult_8_704 ;
wire Xd_0__inst_mult_8_705 ;
wire Xd_0__inst_mult_8_709 ;
wire Xd_0__inst_mult_8_710 ;
wire Xd_0__inst_mult_8_715 ;
wire Xd_0__inst_mult_11_704 ;
wire Xd_0__inst_mult_11_705 ;
wire Xd_0__inst_mult_11_709 ;
wire Xd_0__inst_mult_11_710 ;
wire Xd_0__inst_mult_11_715 ;
wire Xd_0__inst_mult_10_704 ;
wire Xd_0__inst_mult_10_705 ;
wire Xd_0__inst_mult_10_709 ;
wire Xd_0__inst_mult_10_710 ;
wire Xd_0__inst_mult_10_715 ;
wire Xd_0__inst_mult_5_704 ;
wire Xd_0__inst_mult_5_705 ;
wire Xd_0__inst_mult_5_709 ;
wire Xd_0__inst_mult_5_710 ;
wire Xd_0__inst_mult_5_715 ;
wire Xd_0__inst_mult_4_704 ;
wire Xd_0__inst_mult_4_705 ;
wire Xd_0__inst_mult_4_709 ;
wire Xd_0__inst_mult_4_710 ;
wire Xd_0__inst_mult_4_715 ;
wire Xd_0__inst_mult_7_704 ;
wire Xd_0__inst_mult_7_705 ;
wire Xd_0__inst_mult_7_709 ;
wire Xd_0__inst_mult_7_710 ;
wire Xd_0__inst_mult_7_715 ;
wire Xd_0__inst_mult_6_704 ;
wire Xd_0__inst_mult_6_705 ;
wire Xd_0__inst_mult_6_709 ;
wire Xd_0__inst_mult_6_710 ;
wire Xd_0__inst_mult_6_715 ;
wire Xd_0__inst_mult_1_704 ;
wire Xd_0__inst_mult_1_705 ;
wire Xd_0__inst_mult_1_709 ;
wire Xd_0__inst_mult_1_710 ;
wire Xd_0__inst_mult_1_715 ;
wire Xd_0__inst_mult_0_704 ;
wire Xd_0__inst_mult_0_705 ;
wire Xd_0__inst_mult_0_709 ;
wire Xd_0__inst_mult_0_710 ;
wire Xd_0__inst_mult_0_715 ;
wire Xd_0__inst_mult_3_704 ;
wire Xd_0__inst_mult_3_705 ;
wire Xd_0__inst_mult_3_709 ;
wire Xd_0__inst_mult_3_710 ;
wire Xd_0__inst_mult_3_715 ;
wire Xd_0__inst_mult_2_749 ;
wire Xd_0__inst_mult_2_750 ;
wire Xd_0__inst_mult_2_755 ;
wire Xd_0__inst_mult_29_729 ;
wire Xd_0__inst_mult_29_730 ;
wire Xd_0__inst_mult_29_734 ;
wire Xd_0__inst_mult_29_735 ;
wire Xd_0__inst_mult_28_719 ;
wire Xd_0__inst_mult_28_720 ;
wire Xd_0__inst_mult_28_724 ;
wire Xd_0__inst_mult_28_725 ;
wire Xd_0__inst_mult_31_719 ;
wire Xd_0__inst_mult_31_720 ;
wire Xd_0__inst_mult_31_724 ;
wire Xd_0__inst_mult_31_725 ;
wire Xd_0__inst_mult_30_719 ;
wire Xd_0__inst_mult_30_720 ;
wire Xd_0__inst_mult_30_724 ;
wire Xd_0__inst_mult_30_725 ;
wire Xd_0__inst_mult_25_734 ;
wire Xd_0__inst_mult_25_735 ;
wire Xd_0__inst_mult_24_809 ;
wire Xd_0__inst_mult_24_810 ;
wire Xd_0__inst_mult_27_734 ;
wire Xd_0__inst_mult_27_735 ;
wire Xd_0__inst_mult_26_809 ;
wire Xd_0__inst_mult_26_810 ;
wire Xd_0__inst_mult_21_729 ;
wire Xd_0__inst_mult_21_730 ;
wire Xd_0__inst_mult_21_734 ;
wire Xd_0__inst_mult_21_735 ;
wire Xd_0__inst_mult_20_729 ;
wire Xd_0__inst_mult_20_730 ;
wire Xd_0__inst_mult_20_734 ;
wire Xd_0__inst_mult_20_735 ;
wire Xd_0__inst_mult_23_729 ;
wire Xd_0__inst_mult_23_730 ;
wire Xd_0__inst_mult_23_734 ;
wire Xd_0__inst_mult_23_735 ;
wire Xd_0__inst_mult_22_729 ;
wire Xd_0__inst_mult_22_730 ;
wire Xd_0__inst_mult_22_734 ;
wire Xd_0__inst_mult_22_735 ;
wire Xd_0__inst_mult_17_729 ;
wire Xd_0__inst_mult_17_730 ;
wire Xd_0__inst_mult_17_734 ;
wire Xd_0__inst_mult_17_735 ;
wire Xd_0__inst_mult_16_729 ;
wire Xd_0__inst_mult_16_730 ;
wire Xd_0__inst_mult_16_734 ;
wire Xd_0__inst_mult_16_735 ;
wire Xd_0__inst_mult_19_729 ;
wire Xd_0__inst_mult_19_730 ;
wire Xd_0__inst_mult_19_734 ;
wire Xd_0__inst_mult_19_735 ;
wire Xd_0__inst_mult_18_709 ;
wire Xd_0__inst_mult_18_710 ;
wire Xd_0__inst_mult_18_714 ;
wire Xd_0__inst_mult_18_715 ;
wire Xd_0__inst_mult_13_719 ;
wire Xd_0__inst_mult_13_720 ;
wire Xd_0__inst_mult_13_724 ;
wire Xd_0__inst_mult_13_725 ;
wire Xd_0__inst_mult_12_709 ;
wire Xd_0__inst_mult_12_710 ;
wire Xd_0__inst_mult_12_714 ;
wire Xd_0__inst_mult_12_715 ;
wire Xd_0__inst_mult_15_709 ;
wire Xd_0__inst_mult_15_710 ;
wire Xd_0__inst_mult_15_714 ;
wire Xd_0__inst_mult_15_715 ;
wire Xd_0__inst_mult_14_709 ;
wire Xd_0__inst_mult_14_710 ;
wire Xd_0__inst_mult_14_714 ;
wire Xd_0__inst_mult_14_715 ;
wire Xd_0__inst_mult_9_719 ;
wire Xd_0__inst_mult_9_720 ;
wire Xd_0__inst_mult_9_724 ;
wire Xd_0__inst_mult_9_725 ;
wire Xd_0__inst_mult_8_719 ;
wire Xd_0__inst_mult_8_720 ;
wire Xd_0__inst_mult_8_724 ;
wire Xd_0__inst_mult_8_725 ;
wire Xd_0__inst_mult_11_719 ;
wire Xd_0__inst_mult_11_720 ;
wire Xd_0__inst_mult_11_724 ;
wire Xd_0__inst_mult_11_725 ;
wire Xd_0__inst_mult_10_719 ;
wire Xd_0__inst_mult_10_720 ;
wire Xd_0__inst_mult_10_724 ;
wire Xd_0__inst_mult_10_725 ;
wire Xd_0__inst_mult_5_719 ;
wire Xd_0__inst_mult_5_720 ;
wire Xd_0__inst_mult_5_724 ;
wire Xd_0__inst_mult_5_725 ;
wire Xd_0__inst_mult_4_719 ;
wire Xd_0__inst_mult_4_720 ;
wire Xd_0__inst_mult_4_724 ;
wire Xd_0__inst_mult_4_725 ;
wire Xd_0__inst_mult_7_719 ;
wire Xd_0__inst_mult_7_720 ;
wire Xd_0__inst_mult_7_724 ;
wire Xd_0__inst_mult_7_725 ;
wire Xd_0__inst_mult_6_719 ;
wire Xd_0__inst_mult_6_720 ;
wire Xd_0__inst_mult_6_724 ;
wire Xd_0__inst_mult_6_725 ;
wire Xd_0__inst_mult_1_719 ;
wire Xd_0__inst_mult_1_720 ;
wire Xd_0__inst_mult_1_724 ;
wire Xd_0__inst_mult_1_725 ;
wire Xd_0__inst_mult_0_719 ;
wire Xd_0__inst_mult_0_720 ;
wire Xd_0__inst_mult_0_724 ;
wire Xd_0__inst_mult_0_725 ;
wire Xd_0__inst_mult_3_719 ;
wire Xd_0__inst_mult_3_720 ;
wire Xd_0__inst_mult_3_724 ;
wire Xd_0__inst_mult_3_725 ;
wire Xd_0__inst_mult_2_759 ;
wire Xd_0__inst_mult_2_760 ;
wire Xd_0__inst_mult_29_739 ;
wire Xd_0__inst_mult_29_740 ;
wire Xd_0__inst_mult_28_729 ;
wire Xd_0__inst_mult_28_730 ;
wire Xd_0__inst_mult_28_734 ;
wire Xd_0__inst_mult_28_735 ;
wire Xd_0__inst_mult_31_729 ;
wire Xd_0__inst_mult_31_730 ;
wire Xd_0__inst_mult_31_734 ;
wire Xd_0__inst_mult_31_735 ;
wire Xd_0__inst_mult_30_729 ;
wire Xd_0__inst_mult_30_730 ;
wire Xd_0__inst_mult_30_734 ;
wire Xd_0__inst_mult_30_735 ;
wire Xd_0__inst_mult_25_739 ;
wire Xd_0__inst_mult_25_740 ;
wire Xd_0__inst_mult_27_739 ;
wire Xd_0__inst_mult_27_740 ;
wire Xd_0__inst_mult_21_739 ;
wire Xd_0__inst_mult_21_740 ;
wire Xd_0__inst_mult_20_739 ;
wire Xd_0__inst_mult_20_740 ;
wire Xd_0__inst_mult_23_739 ;
wire Xd_0__inst_mult_23_740 ;
wire Xd_0__inst_mult_22_739 ;
wire Xd_0__inst_mult_22_740 ;
wire Xd_0__inst_mult_17_739 ;
wire Xd_0__inst_mult_17_740 ;
wire Xd_0__inst_mult_16_739 ;
wire Xd_0__inst_mult_16_740 ;
wire Xd_0__inst_mult_19_739 ;
wire Xd_0__inst_mult_19_740 ;
wire Xd_0__inst_mult_18_719 ;
wire Xd_0__inst_mult_18_720 ;
wire Xd_0__inst_mult_18_724 ;
wire Xd_0__inst_mult_18_725 ;
wire Xd_0__inst_mult_13_729 ;
wire Xd_0__inst_mult_13_730 ;
wire Xd_0__inst_mult_13_734 ;
wire Xd_0__inst_mult_13_735 ;
wire Xd_0__inst_mult_12_719 ;
wire Xd_0__inst_mult_12_720 ;
wire Xd_0__inst_mult_12_724 ;
wire Xd_0__inst_mult_12_725 ;
wire Xd_0__inst_mult_15_719 ;
wire Xd_0__inst_mult_15_720 ;
wire Xd_0__inst_mult_15_724 ;
wire Xd_0__inst_mult_15_725 ;
wire Xd_0__inst_mult_14_719 ;
wire Xd_0__inst_mult_14_720 ;
wire Xd_0__inst_mult_14_724 ;
wire Xd_0__inst_mult_14_725 ;
wire Xd_0__inst_mult_9_729 ;
wire Xd_0__inst_mult_9_730 ;
wire Xd_0__inst_mult_9_734 ;
wire Xd_0__inst_mult_9_735 ;
wire Xd_0__inst_mult_8_729 ;
wire Xd_0__inst_mult_8_730 ;
wire Xd_0__inst_mult_8_734 ;
wire Xd_0__inst_mult_8_735 ;
wire Xd_0__inst_mult_11_729 ;
wire Xd_0__inst_mult_11_730 ;
wire Xd_0__inst_mult_11_734 ;
wire Xd_0__inst_mult_11_735 ;
wire Xd_0__inst_mult_10_729 ;
wire Xd_0__inst_mult_10_730 ;
wire Xd_0__inst_mult_10_734 ;
wire Xd_0__inst_mult_10_735 ;
wire Xd_0__inst_mult_5_729 ;
wire Xd_0__inst_mult_5_730 ;
wire Xd_0__inst_mult_5_734 ;
wire Xd_0__inst_mult_5_735 ;
wire Xd_0__inst_mult_4_729 ;
wire Xd_0__inst_mult_4_730 ;
wire Xd_0__inst_mult_4_734 ;
wire Xd_0__inst_mult_4_735 ;
wire Xd_0__inst_mult_7_729 ;
wire Xd_0__inst_mult_7_730 ;
wire Xd_0__inst_mult_7_734 ;
wire Xd_0__inst_mult_7_735 ;
wire Xd_0__inst_mult_6_729 ;
wire Xd_0__inst_mult_6_730 ;
wire Xd_0__inst_mult_6_734 ;
wire Xd_0__inst_mult_6_735 ;
wire Xd_0__inst_mult_1_729 ;
wire Xd_0__inst_mult_1_730 ;
wire Xd_0__inst_mult_1_734 ;
wire Xd_0__inst_mult_1_735 ;
wire Xd_0__inst_mult_0_729 ;
wire Xd_0__inst_mult_0_730 ;
wire Xd_0__inst_mult_0_734 ;
wire Xd_0__inst_mult_0_735 ;
wire Xd_0__inst_mult_3_729 ;
wire Xd_0__inst_mult_3_730 ;
wire Xd_0__inst_mult_3_734 ;
wire Xd_0__inst_mult_3_735 ;
wire Xd_0__inst_mult_2_764 ;
wire Xd_0__inst_mult_2_765 ;
wire Xd_0__inst_mult_29_744 ;
wire Xd_0__inst_mult_29_745 ;
wire Xd_0__inst_mult_29_749 ;
wire Xd_0__inst_mult_29_750 ;
wire Xd_0__inst_mult_29_754 ;
wire Xd_0__inst_mult_29_755 ;
wire Xd_0__inst_mult_28_739 ;
wire Xd_0__inst_mult_28_740 ;
wire Xd_0__inst_mult_28_744 ;
wire Xd_0__inst_mult_28_745 ;
wire Xd_0__inst_mult_28_749 ;
wire Xd_0__inst_mult_28_750 ;
wire Xd_0__inst_mult_28_754 ;
wire Xd_0__inst_mult_28_755 ;
wire Xd_0__inst_mult_31_739 ;
wire Xd_0__inst_mult_31_740 ;
wire Xd_0__inst_mult_31_744 ;
wire Xd_0__inst_mult_31_745 ;
wire Xd_0__inst_mult_31_749 ;
wire Xd_0__inst_mult_31_750 ;
wire Xd_0__inst_mult_31_754 ;
wire Xd_0__inst_mult_31_755 ;
wire Xd_0__inst_mult_30_739 ;
wire Xd_0__inst_mult_30_740 ;
wire Xd_0__inst_mult_30_744 ;
wire Xd_0__inst_mult_30_745 ;
wire Xd_0__inst_mult_30_749 ;
wire Xd_0__inst_mult_30_750 ;
wire Xd_0__inst_mult_30_754 ;
wire Xd_0__inst_mult_30_755 ;
wire Xd_0__inst_mult_25_744 ;
wire Xd_0__inst_mult_25_745 ;
wire Xd_0__inst_mult_25_749 ;
wire Xd_0__inst_mult_25_750 ;
wire Xd_0__inst_mult_25_754 ;
wire Xd_0__inst_mult_25_755 ;
wire Xd_0__inst_mult_27_744 ;
wire Xd_0__inst_mult_27_745 ;
wire Xd_0__inst_mult_27_749 ;
wire Xd_0__inst_mult_27_750 ;
wire Xd_0__inst_mult_27_754 ;
wire Xd_0__inst_mult_27_755 ;
wire Xd_0__inst_mult_21_744 ;
wire Xd_0__inst_mult_21_745 ;
wire Xd_0__inst_mult_21_749 ;
wire Xd_0__inst_mult_21_750 ;
wire Xd_0__inst_mult_21_754 ;
wire Xd_0__inst_mult_21_755 ;
wire Xd_0__inst_mult_20_744 ;
wire Xd_0__inst_mult_20_745 ;
wire Xd_0__inst_mult_20_749 ;
wire Xd_0__inst_mult_20_750 ;
wire Xd_0__inst_mult_20_754 ;
wire Xd_0__inst_mult_20_755 ;
wire Xd_0__inst_mult_23_744 ;
wire Xd_0__inst_mult_23_745 ;
wire Xd_0__inst_mult_23_749 ;
wire Xd_0__inst_mult_23_750 ;
wire Xd_0__inst_mult_23_754 ;
wire Xd_0__inst_mult_23_755 ;
wire Xd_0__inst_mult_22_744 ;
wire Xd_0__inst_mult_22_745 ;
wire Xd_0__inst_mult_22_749 ;
wire Xd_0__inst_mult_22_750 ;
wire Xd_0__inst_mult_22_754 ;
wire Xd_0__inst_mult_22_755 ;
wire Xd_0__inst_mult_17_744 ;
wire Xd_0__inst_mult_17_745 ;
wire Xd_0__inst_mult_17_749 ;
wire Xd_0__inst_mult_17_750 ;
wire Xd_0__inst_mult_17_754 ;
wire Xd_0__inst_mult_17_755 ;
wire Xd_0__inst_mult_16_744 ;
wire Xd_0__inst_mult_16_745 ;
wire Xd_0__inst_mult_16_749 ;
wire Xd_0__inst_mult_16_750 ;
wire Xd_0__inst_mult_16_754 ;
wire Xd_0__inst_mult_16_755 ;
wire Xd_0__inst_mult_19_744 ;
wire Xd_0__inst_mult_19_745 ;
wire Xd_0__inst_mult_19_749 ;
wire Xd_0__inst_mult_19_750 ;
wire Xd_0__inst_mult_19_754 ;
wire Xd_0__inst_mult_19_755 ;
wire Xd_0__inst_mult_18_729 ;
wire Xd_0__inst_mult_18_730 ;
wire Xd_0__inst_mult_18_734 ;
wire Xd_0__inst_mult_18_735 ;
wire Xd_0__inst_mult_18_739 ;
wire Xd_0__inst_mult_18_740 ;
wire Xd_0__inst_mult_18_744 ;
wire Xd_0__inst_mult_18_745 ;
wire Xd_0__inst_mult_13_739 ;
wire Xd_0__inst_mult_13_740 ;
wire Xd_0__inst_mult_13_744 ;
wire Xd_0__inst_mult_13_745 ;
wire Xd_0__inst_mult_13_749 ;
wire Xd_0__inst_mult_13_750 ;
wire Xd_0__inst_mult_13_754 ;
wire Xd_0__inst_mult_13_755 ;
wire Xd_0__inst_mult_12_729 ;
wire Xd_0__inst_mult_12_730 ;
wire Xd_0__inst_mult_12_734 ;
wire Xd_0__inst_mult_12_735 ;
wire Xd_0__inst_mult_12_739 ;
wire Xd_0__inst_mult_12_740 ;
wire Xd_0__inst_mult_12_744 ;
wire Xd_0__inst_mult_12_745 ;
wire Xd_0__inst_mult_15_729 ;
wire Xd_0__inst_mult_15_730 ;
wire Xd_0__inst_mult_15_734 ;
wire Xd_0__inst_mult_15_735 ;
wire Xd_0__inst_mult_15_739 ;
wire Xd_0__inst_mult_15_740 ;
wire Xd_0__inst_mult_15_744 ;
wire Xd_0__inst_mult_15_745 ;
wire Xd_0__inst_mult_14_729 ;
wire Xd_0__inst_mult_14_730 ;
wire Xd_0__inst_mult_14_734 ;
wire Xd_0__inst_mult_14_735 ;
wire Xd_0__inst_mult_14_739 ;
wire Xd_0__inst_mult_14_740 ;
wire Xd_0__inst_mult_14_744 ;
wire Xd_0__inst_mult_14_745 ;
wire Xd_0__inst_mult_9_739 ;
wire Xd_0__inst_mult_9_740 ;
wire Xd_0__inst_mult_9_744 ;
wire Xd_0__inst_mult_9_745 ;
wire Xd_0__inst_mult_9_749 ;
wire Xd_0__inst_mult_9_750 ;
wire Xd_0__inst_mult_9_754 ;
wire Xd_0__inst_mult_9_755 ;
wire Xd_0__inst_mult_8_739 ;
wire Xd_0__inst_mult_8_740 ;
wire Xd_0__inst_mult_8_744 ;
wire Xd_0__inst_mult_8_745 ;
wire Xd_0__inst_mult_8_749 ;
wire Xd_0__inst_mult_8_750 ;
wire Xd_0__inst_mult_8_754 ;
wire Xd_0__inst_mult_8_755 ;
wire Xd_0__inst_mult_11_739 ;
wire Xd_0__inst_mult_11_740 ;
wire Xd_0__inst_mult_11_744 ;
wire Xd_0__inst_mult_11_745 ;
wire Xd_0__inst_mult_11_749 ;
wire Xd_0__inst_mult_11_750 ;
wire Xd_0__inst_mult_11_754 ;
wire Xd_0__inst_mult_11_755 ;
wire Xd_0__inst_mult_10_739 ;
wire Xd_0__inst_mult_10_740 ;
wire Xd_0__inst_mult_10_744 ;
wire Xd_0__inst_mult_10_745 ;
wire Xd_0__inst_mult_10_749 ;
wire Xd_0__inst_mult_10_750 ;
wire Xd_0__inst_mult_10_754 ;
wire Xd_0__inst_mult_10_755 ;
wire Xd_0__inst_mult_5_739 ;
wire Xd_0__inst_mult_5_740 ;
wire Xd_0__inst_mult_5_744 ;
wire Xd_0__inst_mult_5_745 ;
wire Xd_0__inst_mult_5_749 ;
wire Xd_0__inst_mult_5_750 ;
wire Xd_0__inst_mult_5_754 ;
wire Xd_0__inst_mult_5_755 ;
wire Xd_0__inst_mult_4_739 ;
wire Xd_0__inst_mult_4_740 ;
wire Xd_0__inst_mult_4_744 ;
wire Xd_0__inst_mult_4_745 ;
wire Xd_0__inst_mult_4_749 ;
wire Xd_0__inst_mult_4_750 ;
wire Xd_0__inst_mult_4_754 ;
wire Xd_0__inst_mult_4_755 ;
wire Xd_0__inst_mult_7_739 ;
wire Xd_0__inst_mult_7_740 ;
wire Xd_0__inst_mult_7_744 ;
wire Xd_0__inst_mult_7_745 ;
wire Xd_0__inst_mult_7_749 ;
wire Xd_0__inst_mult_7_750 ;
wire Xd_0__inst_mult_7_754 ;
wire Xd_0__inst_mult_7_755 ;
wire Xd_0__inst_mult_6_739 ;
wire Xd_0__inst_mult_6_740 ;
wire Xd_0__inst_mult_6_744 ;
wire Xd_0__inst_mult_6_745 ;
wire Xd_0__inst_mult_6_749 ;
wire Xd_0__inst_mult_6_750 ;
wire Xd_0__inst_mult_6_754 ;
wire Xd_0__inst_mult_6_755 ;
wire Xd_0__inst_mult_1_739 ;
wire Xd_0__inst_mult_1_740 ;
wire Xd_0__inst_mult_1_744 ;
wire Xd_0__inst_mult_1_745 ;
wire Xd_0__inst_mult_1_749 ;
wire Xd_0__inst_mult_1_750 ;
wire Xd_0__inst_mult_1_754 ;
wire Xd_0__inst_mult_1_755 ;
wire Xd_0__inst_mult_0_739 ;
wire Xd_0__inst_mult_0_740 ;
wire Xd_0__inst_mult_0_744 ;
wire Xd_0__inst_mult_0_745 ;
wire Xd_0__inst_mult_0_749 ;
wire Xd_0__inst_mult_0_750 ;
wire Xd_0__inst_mult_0_754 ;
wire Xd_0__inst_mult_0_755 ;
wire Xd_0__inst_mult_3_739 ;
wire Xd_0__inst_mult_3_740 ;
wire Xd_0__inst_mult_3_744 ;
wire Xd_0__inst_mult_3_745 ;
wire Xd_0__inst_mult_3_749 ;
wire Xd_0__inst_mult_3_750 ;
wire Xd_0__inst_mult_3_754 ;
wire Xd_0__inst_mult_3_755 ;
wire Xd_0__inst_mult_2_769 ;
wire Xd_0__inst_mult_2_770 ;
wire Xd_0__inst_mult_2_774 ;
wire Xd_0__inst_mult_2_775 ;
wire Xd_0__inst_mult_2_779 ;
wire Xd_0__inst_mult_2_780 ;
wire Xd_0__inst_mult_29_759 ;
wire Xd_0__inst_mult_29_760 ;
wire Xd_0__inst_mult_29_764 ;
wire Xd_0__inst_mult_29_765 ;
wire Xd_0__inst_mult_28_759 ;
wire Xd_0__inst_mult_28_760 ;
wire Xd_0__inst_mult_28_764 ;
wire Xd_0__inst_mult_28_765 ;
wire Xd_0__inst_mult_31_759 ;
wire Xd_0__inst_mult_31_760 ;
wire Xd_0__inst_mult_31_764 ;
wire Xd_0__inst_mult_31_765 ;
wire Xd_0__inst_mult_30_759 ;
wire Xd_0__inst_mult_30_760 ;
wire Xd_0__inst_mult_30_764 ;
wire Xd_0__inst_mult_30_765 ;
wire Xd_0__inst_mult_25_759 ;
wire Xd_0__inst_mult_25_760 ;
wire Xd_0__inst_mult_25_764 ;
wire Xd_0__inst_mult_25_765 ;
wire Xd_0__inst_mult_27_759 ;
wire Xd_0__inst_mult_27_760 ;
wire Xd_0__inst_mult_27_764 ;
wire Xd_0__inst_mult_27_765 ;
wire Xd_0__inst_mult_21_759 ;
wire Xd_0__inst_mult_21_760 ;
wire Xd_0__inst_mult_21_764 ;
wire Xd_0__inst_mult_21_765 ;
wire Xd_0__inst_mult_20_759 ;
wire Xd_0__inst_mult_20_760 ;
wire Xd_0__inst_mult_20_764 ;
wire Xd_0__inst_mult_20_765 ;
wire Xd_0__inst_mult_23_759 ;
wire Xd_0__inst_mult_23_760 ;
wire Xd_0__inst_mult_23_764 ;
wire Xd_0__inst_mult_23_765 ;
wire Xd_0__inst_mult_22_759 ;
wire Xd_0__inst_mult_22_760 ;
wire Xd_0__inst_mult_22_764 ;
wire Xd_0__inst_mult_22_765 ;
wire Xd_0__inst_mult_17_759 ;
wire Xd_0__inst_mult_17_760 ;
wire Xd_0__inst_mult_17_764 ;
wire Xd_0__inst_mult_17_765 ;
wire Xd_0__inst_mult_16_759 ;
wire Xd_0__inst_mult_16_760 ;
wire Xd_0__inst_mult_16_764 ;
wire Xd_0__inst_mult_16_765 ;
wire Xd_0__inst_mult_19_759 ;
wire Xd_0__inst_mult_19_760 ;
wire Xd_0__inst_mult_19_764 ;
wire Xd_0__inst_mult_19_765 ;
wire Xd_0__inst_mult_18_749 ;
wire Xd_0__inst_mult_18_750 ;
wire Xd_0__inst_mult_18_754 ;
wire Xd_0__inst_mult_18_755 ;
wire Xd_0__inst_mult_18_759 ;
wire Xd_0__inst_mult_18_760 ;
wire Xd_0__inst_mult_13_759 ;
wire Xd_0__inst_mult_13_760 ;
wire Xd_0__inst_mult_13_764 ;
wire Xd_0__inst_mult_13_765 ;
wire Xd_0__inst_mult_12_749 ;
wire Xd_0__inst_mult_12_750 ;
wire Xd_0__inst_mult_12_754 ;
wire Xd_0__inst_mult_12_755 ;
wire Xd_0__inst_mult_12_759 ;
wire Xd_0__inst_mult_12_760 ;
wire Xd_0__inst_mult_15_749 ;
wire Xd_0__inst_mult_15_750 ;
wire Xd_0__inst_mult_15_754 ;
wire Xd_0__inst_mult_15_755 ;
wire Xd_0__inst_mult_15_759 ;
wire Xd_0__inst_mult_15_760 ;
wire Xd_0__inst_mult_14_749 ;
wire Xd_0__inst_mult_14_750 ;
wire Xd_0__inst_mult_14_754 ;
wire Xd_0__inst_mult_14_755 ;
wire Xd_0__inst_mult_14_759 ;
wire Xd_0__inst_mult_14_760 ;
wire Xd_0__inst_mult_9_759 ;
wire Xd_0__inst_mult_9_760 ;
wire Xd_0__inst_mult_9_764 ;
wire Xd_0__inst_mult_9_765 ;
wire Xd_0__inst_mult_8_759 ;
wire Xd_0__inst_mult_8_760 ;
wire Xd_0__inst_mult_8_764 ;
wire Xd_0__inst_mult_8_765 ;
wire Xd_0__inst_mult_11_759 ;
wire Xd_0__inst_mult_11_760 ;
wire Xd_0__inst_mult_11_764 ;
wire Xd_0__inst_mult_11_765 ;
wire Xd_0__inst_mult_10_759 ;
wire Xd_0__inst_mult_10_760 ;
wire Xd_0__inst_mult_10_764 ;
wire Xd_0__inst_mult_10_765 ;
wire Xd_0__inst_mult_5_759 ;
wire Xd_0__inst_mult_5_760 ;
wire Xd_0__inst_mult_5_764 ;
wire Xd_0__inst_mult_5_765 ;
wire Xd_0__inst_mult_4_759 ;
wire Xd_0__inst_mult_4_760 ;
wire Xd_0__inst_mult_4_764 ;
wire Xd_0__inst_mult_4_765 ;
wire Xd_0__inst_mult_7_759 ;
wire Xd_0__inst_mult_7_760 ;
wire Xd_0__inst_mult_7_764 ;
wire Xd_0__inst_mult_7_765 ;
wire Xd_0__inst_mult_6_759 ;
wire Xd_0__inst_mult_6_760 ;
wire Xd_0__inst_mult_6_764 ;
wire Xd_0__inst_mult_6_765 ;
wire Xd_0__inst_mult_1_759 ;
wire Xd_0__inst_mult_1_760 ;
wire Xd_0__inst_mult_1_764 ;
wire Xd_0__inst_mult_1_765 ;
wire Xd_0__inst_mult_0_759 ;
wire Xd_0__inst_mult_0_760 ;
wire Xd_0__inst_mult_0_764 ;
wire Xd_0__inst_mult_0_765 ;
wire Xd_0__inst_mult_3_759 ;
wire Xd_0__inst_mult_3_760 ;
wire Xd_0__inst_mult_3_764 ;
wire Xd_0__inst_mult_3_765 ;
wire Xd_0__inst_mult_2_784 ;
wire Xd_0__inst_mult_2_785 ;
wire Xd_0__inst_mult_29_769 ;
wire Xd_0__inst_mult_29_770 ;
wire Xd_0__inst_mult_29_774 ;
wire Xd_0__inst_mult_29_775 ;
wire Xd_0__inst_mult_28_769 ;
wire Xd_0__inst_mult_28_770 ;
wire Xd_0__inst_mult_28_774 ;
wire Xd_0__inst_mult_28_775 ;
wire Xd_0__inst_mult_31_769 ;
wire Xd_0__inst_mult_31_770 ;
wire Xd_0__inst_mult_31_774 ;
wire Xd_0__inst_mult_31_775 ;
wire Xd_0__inst_mult_30_769 ;
wire Xd_0__inst_mult_30_770 ;
wire Xd_0__inst_mult_30_774 ;
wire Xd_0__inst_mult_30_775 ;
wire Xd_0__inst_mult_25_769 ;
wire Xd_0__inst_mult_25_770 ;
wire Xd_0__inst_mult_25_774 ;
wire Xd_0__inst_mult_25_775 ;
wire Xd_0__inst_mult_27_769 ;
wire Xd_0__inst_mult_27_770 ;
wire Xd_0__inst_mult_27_774 ;
wire Xd_0__inst_mult_27_775 ;
wire Xd_0__inst_mult_21_769 ;
wire Xd_0__inst_mult_21_770 ;
wire Xd_0__inst_mult_21_774 ;
wire Xd_0__inst_mult_21_775 ;
wire Xd_0__inst_mult_20_769 ;
wire Xd_0__inst_mult_20_770 ;
wire Xd_0__inst_mult_20_774 ;
wire Xd_0__inst_mult_20_775 ;
wire Xd_0__inst_mult_23_769 ;
wire Xd_0__inst_mult_23_770 ;
wire Xd_0__inst_mult_23_774 ;
wire Xd_0__inst_mult_23_775 ;
wire Xd_0__inst_mult_22_769 ;
wire Xd_0__inst_mult_22_770 ;
wire Xd_0__inst_mult_22_774 ;
wire Xd_0__inst_mult_22_775 ;
wire Xd_0__inst_mult_17_769 ;
wire Xd_0__inst_mult_17_770 ;
wire Xd_0__inst_mult_17_774 ;
wire Xd_0__inst_mult_17_775 ;
wire Xd_0__inst_mult_16_769 ;
wire Xd_0__inst_mult_16_770 ;
wire Xd_0__inst_mult_16_774 ;
wire Xd_0__inst_mult_16_775 ;
wire Xd_0__inst_mult_19_769 ;
wire Xd_0__inst_mult_19_770 ;
wire Xd_0__inst_mult_19_774 ;
wire Xd_0__inst_mult_19_775 ;
wire Xd_0__inst_mult_18_764 ;
wire Xd_0__inst_mult_18_769 ;
wire Xd_0__inst_mult_18_770 ;
wire Xd_0__inst_mult_18_774 ;
wire Xd_0__inst_mult_18_775 ;
wire Xd_0__inst_mult_13_769 ;
wire Xd_0__inst_mult_13_770 ;
wire Xd_0__inst_mult_13_774 ;
wire Xd_0__inst_mult_13_775 ;
wire Xd_0__inst_mult_12_764 ;
wire Xd_0__inst_mult_12_769 ;
wire Xd_0__inst_mult_12_770 ;
wire Xd_0__inst_mult_12_774 ;
wire Xd_0__inst_mult_12_775 ;
wire Xd_0__inst_mult_15_764 ;
wire Xd_0__inst_mult_15_769 ;
wire Xd_0__inst_mult_15_770 ;
wire Xd_0__inst_mult_15_774 ;
wire Xd_0__inst_mult_15_775 ;
wire Xd_0__inst_mult_14_764 ;
wire Xd_0__inst_mult_14_769 ;
wire Xd_0__inst_mult_14_770 ;
wire Xd_0__inst_mult_14_774 ;
wire Xd_0__inst_mult_14_775 ;
wire Xd_0__inst_mult_9_769 ;
wire Xd_0__inst_mult_9_770 ;
wire Xd_0__inst_mult_9_774 ;
wire Xd_0__inst_mult_9_775 ;
wire Xd_0__inst_mult_8_769 ;
wire Xd_0__inst_mult_8_770 ;
wire Xd_0__inst_mult_8_774 ;
wire Xd_0__inst_mult_8_775 ;
wire Xd_0__inst_mult_11_769 ;
wire Xd_0__inst_mult_11_770 ;
wire Xd_0__inst_mult_11_774 ;
wire Xd_0__inst_mult_11_775 ;
wire Xd_0__inst_mult_10_769 ;
wire Xd_0__inst_mult_10_770 ;
wire Xd_0__inst_mult_10_774 ;
wire Xd_0__inst_mult_10_775 ;
wire Xd_0__inst_mult_5_769 ;
wire Xd_0__inst_mult_5_770 ;
wire Xd_0__inst_mult_5_774 ;
wire Xd_0__inst_mult_5_775 ;
wire Xd_0__inst_mult_4_769 ;
wire Xd_0__inst_mult_4_770 ;
wire Xd_0__inst_mult_4_774 ;
wire Xd_0__inst_mult_4_775 ;
wire Xd_0__inst_mult_7_769 ;
wire Xd_0__inst_mult_7_770 ;
wire Xd_0__inst_mult_7_774 ;
wire Xd_0__inst_mult_7_775 ;
wire Xd_0__inst_mult_6_769 ;
wire Xd_0__inst_mult_6_770 ;
wire Xd_0__inst_mult_6_774 ;
wire Xd_0__inst_mult_6_775 ;
wire Xd_0__inst_mult_1_769 ;
wire Xd_0__inst_mult_1_770 ;
wire Xd_0__inst_mult_1_774 ;
wire Xd_0__inst_mult_1_775 ;
wire Xd_0__inst_mult_0_769 ;
wire Xd_0__inst_mult_0_770 ;
wire Xd_0__inst_mult_0_774 ;
wire Xd_0__inst_mult_0_775 ;
wire Xd_0__inst_mult_3_769 ;
wire Xd_0__inst_mult_3_770 ;
wire Xd_0__inst_mult_3_774 ;
wire Xd_0__inst_mult_3_775 ;
wire Xd_0__inst_mult_2_789 ;
wire Xd_0__inst_mult_2_790 ;
wire Xd_0__inst_mult_29_779 ;
wire Xd_0__inst_mult_29_780 ;
wire Xd_0__inst_mult_29_784 ;
wire Xd_0__inst_mult_29_785 ;
wire Xd_0__inst_mult_28_779 ;
wire Xd_0__inst_mult_28_780 ;
wire Xd_0__inst_mult_28_784 ;
wire Xd_0__inst_mult_28_785 ;
wire Xd_0__inst_mult_31_779 ;
wire Xd_0__inst_mult_31_780 ;
wire Xd_0__inst_mult_31_784 ;
wire Xd_0__inst_mult_31_785 ;
wire Xd_0__inst_mult_30_779 ;
wire Xd_0__inst_mult_30_780 ;
wire Xd_0__inst_mult_30_784 ;
wire Xd_0__inst_mult_30_785 ;
wire Xd_0__inst_mult_25_779 ;
wire Xd_0__inst_mult_25_780 ;
wire Xd_0__inst_mult_25_784 ;
wire Xd_0__inst_mult_25_785 ;
wire Xd_0__inst_mult_27_779 ;
wire Xd_0__inst_mult_27_780 ;
wire Xd_0__inst_mult_27_784 ;
wire Xd_0__inst_mult_27_785 ;
wire Xd_0__inst_mult_21_779 ;
wire Xd_0__inst_mult_21_780 ;
wire Xd_0__inst_mult_21_784 ;
wire Xd_0__inst_mult_21_785 ;
wire Xd_0__inst_mult_20_779 ;
wire Xd_0__inst_mult_20_780 ;
wire Xd_0__inst_mult_20_784 ;
wire Xd_0__inst_mult_20_785 ;
wire Xd_0__inst_mult_23_779 ;
wire Xd_0__inst_mult_23_780 ;
wire Xd_0__inst_mult_23_784 ;
wire Xd_0__inst_mult_23_785 ;
wire Xd_0__inst_mult_22_779 ;
wire Xd_0__inst_mult_22_780 ;
wire Xd_0__inst_mult_22_784 ;
wire Xd_0__inst_mult_22_785 ;
wire Xd_0__inst_mult_17_779 ;
wire Xd_0__inst_mult_17_780 ;
wire Xd_0__inst_mult_17_784 ;
wire Xd_0__inst_mult_17_785 ;
wire Xd_0__inst_mult_16_779 ;
wire Xd_0__inst_mult_16_780 ;
wire Xd_0__inst_mult_16_784 ;
wire Xd_0__inst_mult_16_785 ;
wire Xd_0__inst_mult_19_779 ;
wire Xd_0__inst_mult_19_780 ;
wire Xd_0__inst_mult_19_784 ;
wire Xd_0__inst_mult_19_785 ;
wire Xd_0__inst_mult_18_779 ;
wire Xd_0__inst_mult_18_780 ;
wire Xd_0__inst_mult_18_784 ;
wire Xd_0__inst_mult_18_785 ;
wire Xd_0__inst_mult_13_779 ;
wire Xd_0__inst_mult_13_780 ;
wire Xd_0__inst_mult_13_784 ;
wire Xd_0__inst_mult_13_785 ;
wire Xd_0__inst_mult_12_779 ;
wire Xd_0__inst_mult_12_780 ;
wire Xd_0__inst_mult_12_784 ;
wire Xd_0__inst_mult_12_785 ;
wire Xd_0__inst_mult_15_779 ;
wire Xd_0__inst_mult_15_780 ;
wire Xd_0__inst_mult_15_784 ;
wire Xd_0__inst_mult_15_785 ;
wire Xd_0__inst_mult_14_779 ;
wire Xd_0__inst_mult_14_780 ;
wire Xd_0__inst_mult_14_784 ;
wire Xd_0__inst_mult_14_785 ;
wire Xd_0__inst_mult_9_779 ;
wire Xd_0__inst_mult_9_780 ;
wire Xd_0__inst_mult_9_784 ;
wire Xd_0__inst_mult_9_785 ;
wire Xd_0__inst_mult_8_779 ;
wire Xd_0__inst_mult_8_780 ;
wire Xd_0__inst_mult_8_784 ;
wire Xd_0__inst_mult_8_785 ;
wire Xd_0__inst_mult_11_779 ;
wire Xd_0__inst_mult_11_780 ;
wire Xd_0__inst_mult_11_784 ;
wire Xd_0__inst_mult_11_785 ;
wire Xd_0__inst_mult_10_779 ;
wire Xd_0__inst_mult_10_780 ;
wire Xd_0__inst_mult_10_784 ;
wire Xd_0__inst_mult_10_785 ;
wire Xd_0__inst_mult_5_779 ;
wire Xd_0__inst_mult_5_780 ;
wire Xd_0__inst_mult_5_784 ;
wire Xd_0__inst_mult_5_785 ;
wire Xd_0__inst_mult_4_779 ;
wire Xd_0__inst_mult_4_780 ;
wire Xd_0__inst_mult_4_784 ;
wire Xd_0__inst_mult_4_785 ;
wire Xd_0__inst_mult_7_779 ;
wire Xd_0__inst_mult_7_780 ;
wire Xd_0__inst_mult_7_784 ;
wire Xd_0__inst_mult_7_785 ;
wire Xd_0__inst_mult_6_779 ;
wire Xd_0__inst_mult_6_780 ;
wire Xd_0__inst_mult_6_784 ;
wire Xd_0__inst_mult_6_785 ;
wire Xd_0__inst_mult_1_779 ;
wire Xd_0__inst_mult_1_780 ;
wire Xd_0__inst_mult_1_784 ;
wire Xd_0__inst_mult_1_785 ;
wire Xd_0__inst_mult_0_779 ;
wire Xd_0__inst_mult_0_780 ;
wire Xd_0__inst_mult_0_784 ;
wire Xd_0__inst_mult_0_785 ;
wire Xd_0__inst_mult_3_779 ;
wire Xd_0__inst_mult_3_780 ;
wire Xd_0__inst_mult_3_784 ;
wire Xd_0__inst_mult_3_785 ;
wire Xd_0__inst_mult_2_794 ;
wire Xd_0__inst_mult_2_795 ;
wire Xd_0__inst_mult_29_789 ;
wire Xd_0__inst_mult_29_790 ;
wire Xd_0__inst_mult_29_794 ;
wire Xd_0__inst_mult_29_795 ;
wire Xd_0__inst_mult_28_789 ;
wire Xd_0__inst_mult_28_790 ;
wire Xd_0__inst_mult_28_794 ;
wire Xd_0__inst_mult_28_795 ;
wire Xd_0__inst_mult_31_789 ;
wire Xd_0__inst_mult_31_790 ;
wire Xd_0__inst_mult_31_794 ;
wire Xd_0__inst_mult_31_795 ;
wire Xd_0__inst_mult_30_789 ;
wire Xd_0__inst_mult_30_790 ;
wire Xd_0__inst_mult_30_794 ;
wire Xd_0__inst_mult_30_795 ;
wire Xd_0__inst_mult_25_789 ;
wire Xd_0__inst_mult_25_790 ;
wire Xd_0__inst_mult_25_794 ;
wire Xd_0__inst_mult_25_795 ;
wire Xd_0__inst_mult_27_789 ;
wire Xd_0__inst_mult_27_790 ;
wire Xd_0__inst_mult_27_794 ;
wire Xd_0__inst_mult_27_795 ;
wire Xd_0__inst_mult_21_789 ;
wire Xd_0__inst_mult_21_790 ;
wire Xd_0__inst_mult_21_794 ;
wire Xd_0__inst_mult_21_795 ;
wire Xd_0__inst_mult_20_789 ;
wire Xd_0__inst_mult_20_790 ;
wire Xd_0__inst_mult_20_794 ;
wire Xd_0__inst_mult_20_795 ;
wire Xd_0__inst_mult_23_789 ;
wire Xd_0__inst_mult_23_790 ;
wire Xd_0__inst_mult_23_794 ;
wire Xd_0__inst_mult_23_795 ;
wire Xd_0__inst_mult_22_789 ;
wire Xd_0__inst_mult_22_790 ;
wire Xd_0__inst_mult_22_794 ;
wire Xd_0__inst_mult_22_795 ;
wire Xd_0__inst_mult_17_789 ;
wire Xd_0__inst_mult_17_790 ;
wire Xd_0__inst_mult_17_794 ;
wire Xd_0__inst_mult_17_795 ;
wire Xd_0__inst_mult_16_789 ;
wire Xd_0__inst_mult_16_790 ;
wire Xd_0__inst_mult_16_794 ;
wire Xd_0__inst_mult_16_795 ;
wire Xd_0__inst_mult_19_789 ;
wire Xd_0__inst_mult_19_790 ;
wire Xd_0__inst_mult_19_794 ;
wire Xd_0__inst_mult_19_795 ;
wire Xd_0__inst_mult_18_789 ;
wire Xd_0__inst_mult_18_790 ;
wire Xd_0__inst_mult_18_794 ;
wire Xd_0__inst_mult_18_795 ;
wire Xd_0__inst_mult_13_789 ;
wire Xd_0__inst_mult_13_790 ;
wire Xd_0__inst_mult_13_794 ;
wire Xd_0__inst_mult_13_795 ;
wire Xd_0__inst_mult_12_789 ;
wire Xd_0__inst_mult_12_790 ;
wire Xd_0__inst_mult_12_794 ;
wire Xd_0__inst_mult_12_795 ;
wire Xd_0__inst_mult_15_789 ;
wire Xd_0__inst_mult_15_790 ;
wire Xd_0__inst_mult_15_794 ;
wire Xd_0__inst_mult_15_795 ;
wire Xd_0__inst_mult_14_789 ;
wire Xd_0__inst_mult_14_790 ;
wire Xd_0__inst_mult_14_794 ;
wire Xd_0__inst_mult_14_795 ;
wire Xd_0__inst_mult_9_789 ;
wire Xd_0__inst_mult_9_790 ;
wire Xd_0__inst_mult_9_794 ;
wire Xd_0__inst_mult_9_795 ;
wire Xd_0__inst_mult_8_789 ;
wire Xd_0__inst_mult_8_790 ;
wire Xd_0__inst_mult_8_794 ;
wire Xd_0__inst_mult_8_795 ;
wire Xd_0__inst_mult_11_789 ;
wire Xd_0__inst_mult_11_790 ;
wire Xd_0__inst_mult_11_794 ;
wire Xd_0__inst_mult_11_795 ;
wire Xd_0__inst_mult_10_789 ;
wire Xd_0__inst_mult_10_790 ;
wire Xd_0__inst_mult_10_794 ;
wire Xd_0__inst_mult_10_795 ;
wire Xd_0__inst_mult_5_789 ;
wire Xd_0__inst_mult_5_790 ;
wire Xd_0__inst_mult_5_794 ;
wire Xd_0__inst_mult_5_795 ;
wire Xd_0__inst_mult_4_789 ;
wire Xd_0__inst_mult_4_790 ;
wire Xd_0__inst_mult_4_794 ;
wire Xd_0__inst_mult_4_795 ;
wire Xd_0__inst_mult_7_789 ;
wire Xd_0__inst_mult_7_790 ;
wire Xd_0__inst_mult_7_794 ;
wire Xd_0__inst_mult_7_795 ;
wire Xd_0__inst_mult_6_789 ;
wire Xd_0__inst_mult_6_790 ;
wire Xd_0__inst_mult_6_794 ;
wire Xd_0__inst_mult_6_795 ;
wire Xd_0__inst_mult_1_789 ;
wire Xd_0__inst_mult_1_790 ;
wire Xd_0__inst_mult_1_794 ;
wire Xd_0__inst_mult_1_795 ;
wire Xd_0__inst_mult_0_789 ;
wire Xd_0__inst_mult_0_790 ;
wire Xd_0__inst_mult_0_794 ;
wire Xd_0__inst_mult_0_795 ;
wire Xd_0__inst_mult_3_789 ;
wire Xd_0__inst_mult_3_790 ;
wire Xd_0__inst_mult_3_794 ;
wire Xd_0__inst_mult_3_795 ;
wire Xd_0__inst_mult_2_799 ;
wire Xd_0__inst_mult_2_800 ;
wire Xd_0__inst_mult_29_799 ;
wire Xd_0__inst_mult_29_804 ;
wire Xd_0__inst_mult_29_805 ;
wire Xd_0__inst_mult_28_799 ;
wire Xd_0__inst_mult_28_804 ;
wire Xd_0__inst_mult_28_805 ;
wire Xd_0__inst_mult_31_799 ;
wire Xd_0__inst_mult_31_804 ;
wire Xd_0__inst_mult_31_805 ;
wire Xd_0__inst_mult_30_799 ;
wire Xd_0__inst_mult_30_804 ;
wire Xd_0__inst_mult_30_805 ;
wire Xd_0__inst_mult_25_799 ;
wire Xd_0__inst_mult_25_804 ;
wire Xd_0__inst_mult_25_805 ;
wire Xd_0__inst_mult_27_799 ;
wire Xd_0__inst_mult_27_804 ;
wire Xd_0__inst_mult_27_805 ;
wire Xd_0__inst_mult_21_799 ;
wire Xd_0__inst_mult_21_804 ;
wire Xd_0__inst_mult_21_805 ;
wire Xd_0__inst_mult_20_799 ;
wire Xd_0__inst_mult_20_804 ;
wire Xd_0__inst_mult_20_805 ;
wire Xd_0__inst_mult_23_799 ;
wire Xd_0__inst_mult_23_804 ;
wire Xd_0__inst_mult_23_805 ;
wire Xd_0__inst_mult_22_799 ;
wire Xd_0__inst_mult_22_804 ;
wire Xd_0__inst_mult_22_805 ;
wire Xd_0__inst_mult_17_799 ;
wire Xd_0__inst_mult_17_804 ;
wire Xd_0__inst_mult_17_805 ;
wire Xd_0__inst_mult_16_799 ;
wire Xd_0__inst_mult_16_804 ;
wire Xd_0__inst_mult_16_805 ;
wire Xd_0__inst_mult_19_799 ;
wire Xd_0__inst_mult_19_804 ;
wire Xd_0__inst_mult_19_805 ;
wire Xd_0__inst_mult_18_799 ;
wire Xd_0__inst_mult_18_804 ;
wire Xd_0__inst_mult_18_805 ;
wire Xd_0__inst_mult_13_799 ;
wire Xd_0__inst_mult_13_804 ;
wire Xd_0__inst_mult_13_805 ;
wire Xd_0__inst_mult_12_799 ;
wire Xd_0__inst_mult_12_804 ;
wire Xd_0__inst_mult_12_805 ;
wire Xd_0__inst_mult_15_799 ;
wire Xd_0__inst_mult_15_804 ;
wire Xd_0__inst_mult_15_805 ;
wire Xd_0__inst_mult_14_799 ;
wire Xd_0__inst_mult_14_804 ;
wire Xd_0__inst_mult_14_805 ;
wire Xd_0__inst_mult_9_799 ;
wire Xd_0__inst_mult_9_804 ;
wire Xd_0__inst_mult_9_805 ;
wire Xd_0__inst_mult_8_799 ;
wire Xd_0__inst_mult_8_804 ;
wire Xd_0__inst_mult_8_805 ;
wire Xd_0__inst_mult_11_799 ;
wire Xd_0__inst_mult_11_804 ;
wire Xd_0__inst_mult_11_805 ;
wire Xd_0__inst_mult_10_799 ;
wire Xd_0__inst_mult_10_804 ;
wire Xd_0__inst_mult_10_805 ;
wire Xd_0__inst_mult_5_799 ;
wire Xd_0__inst_mult_5_804 ;
wire Xd_0__inst_mult_5_805 ;
wire Xd_0__inst_mult_4_799 ;
wire Xd_0__inst_mult_4_804 ;
wire Xd_0__inst_mult_4_805 ;
wire Xd_0__inst_mult_7_799 ;
wire Xd_0__inst_mult_7_804 ;
wire Xd_0__inst_mult_7_805 ;
wire Xd_0__inst_mult_6_799 ;
wire Xd_0__inst_mult_6_804 ;
wire Xd_0__inst_mult_6_805 ;
wire Xd_0__inst_mult_1_799 ;
wire Xd_0__inst_mult_1_804 ;
wire Xd_0__inst_mult_1_805 ;
wire Xd_0__inst_mult_0_799 ;
wire Xd_0__inst_mult_0_804 ;
wire Xd_0__inst_mult_0_805 ;
wire Xd_0__inst_mult_3_799 ;
wire Xd_0__inst_mult_3_804 ;
wire Xd_0__inst_mult_3_805 ;
wire Xd_0__inst_mult_2_804 ;
wire Xd_0__inst_mult_2_805 ;
wire Xd_0__inst_mult_29_809 ;
wire Xd_0__inst_mult_29_810 ;
wire Xd_0__inst_mult_28_809 ;
wire Xd_0__inst_mult_28_810 ;
wire Xd_0__inst_mult_31_809 ;
wire Xd_0__inst_mult_31_810 ;
wire Xd_0__inst_mult_30_809 ;
wire Xd_0__inst_mult_30_810 ;
wire Xd_0__inst_mult_25_809 ;
wire Xd_0__inst_mult_25_810 ;
wire Xd_0__inst_mult_27_809 ;
wire Xd_0__inst_mult_27_810 ;
wire Xd_0__inst_mult_21_809 ;
wire Xd_0__inst_mult_21_810 ;
wire Xd_0__inst_mult_20_809 ;
wire Xd_0__inst_mult_20_810 ;
wire Xd_0__inst_mult_23_809 ;
wire Xd_0__inst_mult_23_810 ;
wire Xd_0__inst_mult_22_809 ;
wire Xd_0__inst_mult_22_810 ;
wire Xd_0__inst_mult_17_809 ;
wire Xd_0__inst_mult_17_810 ;
wire Xd_0__inst_mult_16_809 ;
wire Xd_0__inst_mult_16_810 ;
wire Xd_0__inst_mult_19_809 ;
wire Xd_0__inst_mult_19_810 ;
wire Xd_0__inst_mult_18_809 ;
wire Xd_0__inst_mult_18_810 ;
wire Xd_0__inst_mult_13_809 ;
wire Xd_0__inst_mult_13_810 ;
wire Xd_0__inst_mult_12_809 ;
wire Xd_0__inst_mult_12_810 ;
wire Xd_0__inst_mult_15_809 ;
wire Xd_0__inst_mult_15_810 ;
wire Xd_0__inst_mult_14_809 ;
wire Xd_0__inst_mult_14_810 ;
wire Xd_0__inst_mult_9_809 ;
wire Xd_0__inst_mult_9_810 ;
wire Xd_0__inst_mult_8_809 ;
wire Xd_0__inst_mult_8_810 ;
wire Xd_0__inst_mult_11_809 ;
wire Xd_0__inst_mult_11_810 ;
wire Xd_0__inst_mult_10_809 ;
wire Xd_0__inst_mult_10_810 ;
wire Xd_0__inst_mult_5_809 ;
wire Xd_0__inst_mult_5_810 ;
wire Xd_0__inst_mult_4_809 ;
wire Xd_0__inst_mult_4_810 ;
wire Xd_0__inst_mult_7_809 ;
wire Xd_0__inst_mult_7_810 ;
wire Xd_0__inst_mult_6_809 ;
wire Xd_0__inst_mult_6_810 ;
wire Xd_0__inst_mult_1_809 ;
wire Xd_0__inst_mult_1_810 ;
wire Xd_0__inst_mult_0_809 ;
wire Xd_0__inst_mult_0_810 ;
wire Xd_0__inst_mult_3_809 ;
wire Xd_0__inst_mult_3_810 ;
wire Xd_0__inst_mult_2_809 ;
wire Xd_0__inst_mult_2_810 ;
wire Xd_0__inst_inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_inst_first_level_1__18__q ;
wire Xd_0__inst_inst_inst_first_level_0__18__q ;
wire Xd_0__inst_inst_inst_first_level_1__19__q ;
wire Xd_0__inst_inst_inst_first_level_0__19__q ;
wire Xd_0__inst_inst_inst_first_level_1__20__q ;
wire Xd_0__inst_inst_inst_first_level_0__20__q ;
wire Xd_0__inst_inst_inst_first_level_1__21__q ;
wire Xd_0__inst_inst_inst_first_level_0__21__q ;
wire Xd_0__inst_inst_inst_first_level_1__22__q ;
wire Xd_0__inst_inst_inst_first_level_0__22__q ;
wire Xd_0__inst_inst_inst_first_level_1__23__q ;
wire Xd_0__inst_inst_inst_first_level_0__23__q ;
wire Xd_0__inst_inst_inst_first_level_1__24__q ;
wire Xd_0__inst_inst_inst_first_level_0__24__q ;
wire Xd_0__inst_inst_inst_first_level_1__25__q ;
wire Xd_0__inst_inst_inst_first_level_0__25__q ;
wire Xd_0__inst_inst_inst_first_level_1__26__q ;
wire Xd_0__inst_inst_inst_first_level_0__26__q ;
wire Xd_0__inst_inst_first_level_3__0__q ;
wire Xd_0__inst_inst_first_level_2__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_3__1__q ;
wire Xd_0__inst_inst_first_level_2__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_3__2__q ;
wire Xd_0__inst_inst_first_level_2__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_3__3__q ;
wire Xd_0__inst_inst_first_level_2__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_3__4__q ;
wire Xd_0__inst_inst_first_level_2__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_3__5__q ;
wire Xd_0__inst_inst_first_level_2__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_3__6__q ;
wire Xd_0__inst_inst_first_level_2__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_3__7__q ;
wire Xd_0__inst_inst_first_level_2__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_3__8__q ;
wire Xd_0__inst_inst_first_level_2__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_3__9__q ;
wire Xd_0__inst_inst_first_level_2__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_3__10__q ;
wire Xd_0__inst_inst_first_level_2__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_3__11__q ;
wire Xd_0__inst_inst_first_level_2__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_3__12__q ;
wire Xd_0__inst_inst_first_level_2__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_3__13__q ;
wire Xd_0__inst_inst_first_level_2__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_3__14__q ;
wire Xd_0__inst_inst_first_level_2__14__q ;
wire Xd_0__inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_first_level_3__15__q ;
wire Xd_0__inst_inst_first_level_2__15__q ;
wire Xd_0__inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_first_level_3__16__q ;
wire Xd_0__inst_inst_first_level_2__16__q ;
wire Xd_0__inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_first_level_3__17__q ;
wire Xd_0__inst_inst_first_level_2__17__q ;
wire Xd_0__inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_first_level_3__18__q ;
wire Xd_0__inst_inst_first_level_2__18__q ;
wire Xd_0__inst_inst_first_level_1__18__q ;
wire Xd_0__inst_inst_first_level_0__18__q ;
wire Xd_0__inst_inst_first_level_3__19__q ;
wire Xd_0__inst_inst_first_level_2__19__q ;
wire Xd_0__inst_inst_first_level_1__19__q ;
wire Xd_0__inst_inst_first_level_0__19__q ;
wire Xd_0__inst_inst_first_level_3__20__q ;
wire Xd_0__inst_inst_first_level_2__20__q ;
wire Xd_0__inst_inst_first_level_1__20__q ;
wire Xd_0__inst_inst_first_level_0__20__q ;
wire Xd_0__inst_inst_first_level_3__21__q ;
wire Xd_0__inst_inst_first_level_2__21__q ;
wire Xd_0__inst_inst_first_level_1__21__q ;
wire Xd_0__inst_inst_first_level_0__21__q ;
wire Xd_0__inst_inst_first_level_3__22__q ;
wire Xd_0__inst_inst_first_level_2__22__q ;
wire Xd_0__inst_inst_first_level_1__22__q ;
wire Xd_0__inst_inst_first_level_0__22__q ;
wire Xd_0__inst_inst_first_level_3__23__q ;
wire Xd_0__inst_inst_first_level_2__23__q ;
wire Xd_0__inst_inst_first_level_1__23__q ;
wire Xd_0__inst_inst_first_level_0__23__q ;
wire Xd_0__inst_inst_first_level_3__24__q ;
wire Xd_0__inst_inst_first_level_2__24__q ;
wire Xd_0__inst_inst_first_level_1__24__q ;
wire Xd_0__inst_inst_first_level_0__24__q ;
wire Xd_0__inst_inst_first_level_3__25__q ;
wire Xd_0__inst_inst_first_level_2__25__q ;
wire Xd_0__inst_inst_first_level_1__25__q ;
wire Xd_0__inst_inst_first_level_0__25__q ;
wire Xd_0__inst_r_sum2_7__0__q ;
wire Xd_0__inst_r_sum2_6__0__q ;
wire Xd_0__inst_r_sum2_5__0__q ;
wire Xd_0__inst_r_sum2_4__0__q ;
wire Xd_0__inst_r_sum2_3__0__q ;
wire Xd_0__inst_r_sum2_2__0__q ;
wire Xd_0__inst_r_sum2_1__0__q ;
wire Xd_0__inst_r_sum2_0__0__q ;
wire Xd_0__inst_r_sum2_7__1__q ;
wire Xd_0__inst_r_sum2_6__1__q ;
wire Xd_0__inst_r_sum2_5__1__q ;
wire Xd_0__inst_r_sum2_4__1__q ;
wire Xd_0__inst_r_sum2_3__1__q ;
wire Xd_0__inst_r_sum2_2__1__q ;
wire Xd_0__inst_r_sum2_1__1__q ;
wire Xd_0__inst_r_sum2_0__1__q ;
wire Xd_0__inst_r_sum2_7__2__q ;
wire Xd_0__inst_r_sum2_6__2__q ;
wire Xd_0__inst_r_sum2_5__2__q ;
wire Xd_0__inst_r_sum2_4__2__q ;
wire Xd_0__inst_r_sum2_3__2__q ;
wire Xd_0__inst_r_sum2_2__2__q ;
wire Xd_0__inst_r_sum2_1__2__q ;
wire Xd_0__inst_r_sum2_0__2__q ;
wire Xd_0__inst_r_sum2_7__3__q ;
wire Xd_0__inst_r_sum2_6__3__q ;
wire Xd_0__inst_r_sum2_5__3__q ;
wire Xd_0__inst_r_sum2_4__3__q ;
wire Xd_0__inst_r_sum2_3__3__q ;
wire Xd_0__inst_r_sum2_2__3__q ;
wire Xd_0__inst_r_sum2_1__3__q ;
wire Xd_0__inst_r_sum2_0__3__q ;
wire Xd_0__inst_r_sum2_7__4__q ;
wire Xd_0__inst_r_sum2_6__4__q ;
wire Xd_0__inst_r_sum2_5__4__q ;
wire Xd_0__inst_r_sum2_4__4__q ;
wire Xd_0__inst_r_sum2_3__4__q ;
wire Xd_0__inst_r_sum2_2__4__q ;
wire Xd_0__inst_r_sum2_1__4__q ;
wire Xd_0__inst_r_sum2_0__4__q ;
wire Xd_0__inst_r_sum2_7__5__q ;
wire Xd_0__inst_r_sum2_6__5__q ;
wire Xd_0__inst_r_sum2_5__5__q ;
wire Xd_0__inst_r_sum2_4__5__q ;
wire Xd_0__inst_r_sum2_3__5__q ;
wire Xd_0__inst_r_sum2_2__5__q ;
wire Xd_0__inst_r_sum2_1__5__q ;
wire Xd_0__inst_r_sum2_0__5__q ;
wire Xd_0__inst_r_sum2_7__6__q ;
wire Xd_0__inst_r_sum2_6__6__q ;
wire Xd_0__inst_r_sum2_5__6__q ;
wire Xd_0__inst_r_sum2_4__6__q ;
wire Xd_0__inst_r_sum2_3__6__q ;
wire Xd_0__inst_r_sum2_2__6__q ;
wire Xd_0__inst_r_sum2_1__6__q ;
wire Xd_0__inst_r_sum2_0__6__q ;
wire Xd_0__inst_r_sum2_7__7__q ;
wire Xd_0__inst_r_sum2_6__7__q ;
wire Xd_0__inst_r_sum2_5__7__q ;
wire Xd_0__inst_r_sum2_4__7__q ;
wire Xd_0__inst_r_sum2_3__7__q ;
wire Xd_0__inst_r_sum2_2__7__q ;
wire Xd_0__inst_r_sum2_1__7__q ;
wire Xd_0__inst_r_sum2_0__7__q ;
wire Xd_0__inst_r_sum2_7__8__q ;
wire Xd_0__inst_r_sum2_6__8__q ;
wire Xd_0__inst_r_sum2_5__8__q ;
wire Xd_0__inst_r_sum2_4__8__q ;
wire Xd_0__inst_r_sum2_3__8__q ;
wire Xd_0__inst_r_sum2_2__8__q ;
wire Xd_0__inst_r_sum2_1__8__q ;
wire Xd_0__inst_r_sum2_0__8__q ;
wire Xd_0__inst_r_sum2_7__9__q ;
wire Xd_0__inst_r_sum2_6__9__q ;
wire Xd_0__inst_r_sum2_5__9__q ;
wire Xd_0__inst_r_sum2_4__9__q ;
wire Xd_0__inst_r_sum2_3__9__q ;
wire Xd_0__inst_r_sum2_2__9__q ;
wire Xd_0__inst_r_sum2_1__9__q ;
wire Xd_0__inst_r_sum2_0__9__q ;
wire Xd_0__inst_r_sum2_7__10__q ;
wire Xd_0__inst_r_sum2_6__10__q ;
wire Xd_0__inst_r_sum2_5__10__q ;
wire Xd_0__inst_r_sum2_4__10__q ;
wire Xd_0__inst_r_sum2_3__10__q ;
wire Xd_0__inst_r_sum2_2__10__q ;
wire Xd_0__inst_r_sum2_1__10__q ;
wire Xd_0__inst_r_sum2_0__10__q ;
wire Xd_0__inst_r_sum2_7__11__q ;
wire Xd_0__inst_r_sum2_6__11__q ;
wire Xd_0__inst_r_sum2_5__11__q ;
wire Xd_0__inst_r_sum2_4__11__q ;
wire Xd_0__inst_r_sum2_3__11__q ;
wire Xd_0__inst_r_sum2_2__11__q ;
wire Xd_0__inst_r_sum2_1__11__q ;
wire Xd_0__inst_r_sum2_0__11__q ;
wire Xd_0__inst_r_sum2_7__12__q ;
wire Xd_0__inst_r_sum2_6__12__q ;
wire Xd_0__inst_r_sum2_5__12__q ;
wire Xd_0__inst_r_sum2_4__12__q ;
wire Xd_0__inst_r_sum2_3__12__q ;
wire Xd_0__inst_r_sum2_2__12__q ;
wire Xd_0__inst_r_sum2_1__12__q ;
wire Xd_0__inst_r_sum2_0__12__q ;
wire Xd_0__inst_r_sum2_7__13__q ;
wire Xd_0__inst_r_sum2_6__13__q ;
wire Xd_0__inst_r_sum2_5__13__q ;
wire Xd_0__inst_r_sum2_4__13__q ;
wire Xd_0__inst_r_sum2_3__13__q ;
wire Xd_0__inst_r_sum2_2__13__q ;
wire Xd_0__inst_r_sum2_1__13__q ;
wire Xd_0__inst_r_sum2_0__13__q ;
wire Xd_0__inst_r_sum2_7__14__q ;
wire Xd_0__inst_r_sum2_6__14__q ;
wire Xd_0__inst_r_sum2_5__14__q ;
wire Xd_0__inst_r_sum2_4__14__q ;
wire Xd_0__inst_r_sum2_3__14__q ;
wire Xd_0__inst_r_sum2_2__14__q ;
wire Xd_0__inst_r_sum2_1__14__q ;
wire Xd_0__inst_r_sum2_0__14__q ;
wire Xd_0__inst_r_sum2_7__15__q ;
wire Xd_0__inst_r_sum2_6__15__q ;
wire Xd_0__inst_r_sum2_5__15__q ;
wire Xd_0__inst_r_sum2_4__15__q ;
wire Xd_0__inst_r_sum2_3__15__q ;
wire Xd_0__inst_r_sum2_2__15__q ;
wire Xd_0__inst_r_sum2_1__15__q ;
wire Xd_0__inst_r_sum2_0__15__q ;
wire Xd_0__inst_r_sum2_7__16__q ;
wire Xd_0__inst_r_sum2_6__16__q ;
wire Xd_0__inst_r_sum2_5__16__q ;
wire Xd_0__inst_r_sum2_4__16__q ;
wire Xd_0__inst_r_sum2_3__16__q ;
wire Xd_0__inst_r_sum2_2__16__q ;
wire Xd_0__inst_r_sum2_1__16__q ;
wire Xd_0__inst_r_sum2_0__16__q ;
wire Xd_0__inst_r_sum2_7__17__q ;
wire Xd_0__inst_r_sum2_6__17__q ;
wire Xd_0__inst_r_sum2_5__17__q ;
wire Xd_0__inst_r_sum2_4__17__q ;
wire Xd_0__inst_r_sum2_3__17__q ;
wire Xd_0__inst_r_sum2_2__17__q ;
wire Xd_0__inst_r_sum2_1__17__q ;
wire Xd_0__inst_r_sum2_0__17__q ;
wire Xd_0__inst_r_sum2_7__18__q ;
wire Xd_0__inst_r_sum2_6__18__q ;
wire Xd_0__inst_r_sum2_5__18__q ;
wire Xd_0__inst_r_sum2_4__18__q ;
wire Xd_0__inst_r_sum2_3__18__q ;
wire Xd_0__inst_r_sum2_2__18__q ;
wire Xd_0__inst_r_sum2_1__18__q ;
wire Xd_0__inst_r_sum2_0__18__q ;
wire Xd_0__inst_r_sum2_7__19__q ;
wire Xd_0__inst_r_sum2_6__19__q ;
wire Xd_0__inst_r_sum2_5__19__q ;
wire Xd_0__inst_r_sum2_4__19__q ;
wire Xd_0__inst_r_sum2_3__19__q ;
wire Xd_0__inst_r_sum2_2__19__q ;
wire Xd_0__inst_r_sum2_1__19__q ;
wire Xd_0__inst_r_sum2_0__19__q ;
wire Xd_0__inst_r_sum2_7__20__q ;
wire Xd_0__inst_r_sum2_6__20__q ;
wire Xd_0__inst_r_sum2_5__20__q ;
wire Xd_0__inst_r_sum2_4__20__q ;
wire Xd_0__inst_r_sum2_3__20__q ;
wire Xd_0__inst_r_sum2_2__20__q ;
wire Xd_0__inst_r_sum2_1__20__q ;
wire Xd_0__inst_r_sum2_0__20__q ;
wire Xd_0__inst_r_sum2_7__21__q ;
wire Xd_0__inst_r_sum2_6__21__q ;
wire Xd_0__inst_r_sum2_5__21__q ;
wire Xd_0__inst_r_sum2_4__21__q ;
wire Xd_0__inst_r_sum2_3__21__q ;
wire Xd_0__inst_r_sum2_2__21__q ;
wire Xd_0__inst_r_sum2_1__21__q ;
wire Xd_0__inst_r_sum2_0__21__q ;
wire Xd_0__inst_r_sum2_7__22__q ;
wire Xd_0__inst_r_sum2_6__22__q ;
wire Xd_0__inst_r_sum2_5__22__q ;
wire Xd_0__inst_r_sum2_4__22__q ;
wire Xd_0__inst_r_sum2_3__22__q ;
wire Xd_0__inst_r_sum2_2__22__q ;
wire Xd_0__inst_r_sum2_1__22__q ;
wire Xd_0__inst_r_sum2_0__22__q ;
wire Xd_0__inst_r_sum2_7__23__q ;
wire Xd_0__inst_r_sum2_6__23__q ;
wire Xd_0__inst_r_sum2_5__23__q ;
wire Xd_0__inst_r_sum2_4__23__q ;
wire Xd_0__inst_r_sum2_3__23__q ;
wire Xd_0__inst_r_sum2_2__23__q ;
wire Xd_0__inst_r_sum2_1__23__q ;
wire Xd_0__inst_r_sum2_0__23__q ;
wire Xd_0__inst_r_sum2_7__24__q ;
wire Xd_0__inst_r_sum2_6__24__q ;
wire Xd_0__inst_r_sum2_5__24__q ;
wire Xd_0__inst_r_sum2_4__24__q ;
wire Xd_0__inst_r_sum2_3__24__q ;
wire Xd_0__inst_r_sum2_2__24__q ;
wire Xd_0__inst_r_sum2_1__24__q ;
wire Xd_0__inst_r_sum2_0__24__q ;
wire Xd_0__inst_r_sum1_15__0__q ;
wire Xd_0__inst_r_sum1_14__0__q ;
wire Xd_0__inst_r_sum1_13__0__q ;
wire Xd_0__inst_r_sum1_12__0__q ;
wire Xd_0__inst_r_sum1_11__0__q ;
wire Xd_0__inst_r_sum1_10__0__q ;
wire Xd_0__inst_r_sum1_9__0__q ;
wire Xd_0__inst_r_sum1_8__0__q ;
wire Xd_0__inst_r_sum1_7__0__q ;
wire Xd_0__inst_r_sum1_6__0__q ;
wire Xd_0__inst_r_sum1_5__0__q ;
wire Xd_0__inst_r_sum1_4__0__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_14__1__q ;
wire Xd_0__inst_r_sum1_15__1__q ;
wire Xd_0__inst_r_sum1_12__1__q ;
wire Xd_0__inst_r_sum1_13__1__q ;
wire Xd_0__inst_r_sum1_10__1__q ;
wire Xd_0__inst_r_sum1_11__1__q ;
wire Xd_0__inst_r_sum1_8__1__q ;
wire Xd_0__inst_r_sum1_9__1__q ;
wire Xd_0__inst_r_sum1_6__1__q ;
wire Xd_0__inst_r_sum1_7__1__q ;
wire Xd_0__inst_r_sum1_4__1__q ;
wire Xd_0__inst_r_sum1_5__1__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_14__2__q ;
wire Xd_0__inst_r_sum1_15__2__q ;
wire Xd_0__inst_r_sum1_12__2__q ;
wire Xd_0__inst_r_sum1_13__2__q ;
wire Xd_0__inst_r_sum1_10__2__q ;
wire Xd_0__inst_r_sum1_11__2__q ;
wire Xd_0__inst_r_sum1_8__2__q ;
wire Xd_0__inst_r_sum1_9__2__q ;
wire Xd_0__inst_r_sum1_6__2__q ;
wire Xd_0__inst_r_sum1_7__2__q ;
wire Xd_0__inst_r_sum1_4__2__q ;
wire Xd_0__inst_r_sum1_5__2__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_14__3__q ;
wire Xd_0__inst_r_sum1_15__3__q ;
wire Xd_0__inst_r_sum1_12__3__q ;
wire Xd_0__inst_r_sum1_13__3__q ;
wire Xd_0__inst_r_sum1_10__3__q ;
wire Xd_0__inst_r_sum1_11__3__q ;
wire Xd_0__inst_r_sum1_8__3__q ;
wire Xd_0__inst_r_sum1_9__3__q ;
wire Xd_0__inst_r_sum1_6__3__q ;
wire Xd_0__inst_r_sum1_7__3__q ;
wire Xd_0__inst_r_sum1_4__3__q ;
wire Xd_0__inst_r_sum1_5__3__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_14__4__q ;
wire Xd_0__inst_r_sum1_15__4__q ;
wire Xd_0__inst_r_sum1_12__4__q ;
wire Xd_0__inst_r_sum1_13__4__q ;
wire Xd_0__inst_r_sum1_10__4__q ;
wire Xd_0__inst_r_sum1_11__4__q ;
wire Xd_0__inst_r_sum1_8__4__q ;
wire Xd_0__inst_r_sum1_9__4__q ;
wire Xd_0__inst_r_sum1_6__4__q ;
wire Xd_0__inst_r_sum1_7__4__q ;
wire Xd_0__inst_r_sum1_4__4__q ;
wire Xd_0__inst_r_sum1_5__4__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_14__5__q ;
wire Xd_0__inst_r_sum1_15__5__q ;
wire Xd_0__inst_r_sum1_12__5__q ;
wire Xd_0__inst_r_sum1_13__5__q ;
wire Xd_0__inst_r_sum1_10__5__q ;
wire Xd_0__inst_r_sum1_11__5__q ;
wire Xd_0__inst_r_sum1_8__5__q ;
wire Xd_0__inst_r_sum1_9__5__q ;
wire Xd_0__inst_r_sum1_6__5__q ;
wire Xd_0__inst_r_sum1_7__5__q ;
wire Xd_0__inst_r_sum1_4__5__q ;
wire Xd_0__inst_r_sum1_5__5__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_14__6__q ;
wire Xd_0__inst_r_sum1_15__6__q ;
wire Xd_0__inst_r_sum1_12__6__q ;
wire Xd_0__inst_r_sum1_13__6__q ;
wire Xd_0__inst_r_sum1_10__6__q ;
wire Xd_0__inst_r_sum1_11__6__q ;
wire Xd_0__inst_r_sum1_8__6__q ;
wire Xd_0__inst_r_sum1_9__6__q ;
wire Xd_0__inst_r_sum1_6__6__q ;
wire Xd_0__inst_r_sum1_7__6__q ;
wire Xd_0__inst_r_sum1_4__6__q ;
wire Xd_0__inst_r_sum1_5__6__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_14__7__q ;
wire Xd_0__inst_r_sum1_15__7__q ;
wire Xd_0__inst_r_sum1_12__7__q ;
wire Xd_0__inst_r_sum1_13__7__q ;
wire Xd_0__inst_r_sum1_10__7__q ;
wire Xd_0__inst_r_sum1_11__7__q ;
wire Xd_0__inst_r_sum1_8__7__q ;
wire Xd_0__inst_r_sum1_9__7__q ;
wire Xd_0__inst_r_sum1_6__7__q ;
wire Xd_0__inst_r_sum1_7__7__q ;
wire Xd_0__inst_r_sum1_4__7__q ;
wire Xd_0__inst_r_sum1_5__7__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_14__8__q ;
wire Xd_0__inst_r_sum1_15__8__q ;
wire Xd_0__inst_r_sum1_12__8__q ;
wire Xd_0__inst_r_sum1_13__8__q ;
wire Xd_0__inst_r_sum1_10__8__q ;
wire Xd_0__inst_r_sum1_11__8__q ;
wire Xd_0__inst_r_sum1_8__8__q ;
wire Xd_0__inst_r_sum1_9__8__q ;
wire Xd_0__inst_r_sum1_6__8__q ;
wire Xd_0__inst_r_sum1_7__8__q ;
wire Xd_0__inst_r_sum1_4__8__q ;
wire Xd_0__inst_r_sum1_5__8__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_14__9__q ;
wire Xd_0__inst_r_sum1_15__9__q ;
wire Xd_0__inst_r_sum1_12__9__q ;
wire Xd_0__inst_r_sum1_13__9__q ;
wire Xd_0__inst_r_sum1_10__9__q ;
wire Xd_0__inst_r_sum1_11__9__q ;
wire Xd_0__inst_r_sum1_8__9__q ;
wire Xd_0__inst_r_sum1_9__9__q ;
wire Xd_0__inst_r_sum1_6__9__q ;
wire Xd_0__inst_r_sum1_7__9__q ;
wire Xd_0__inst_r_sum1_4__9__q ;
wire Xd_0__inst_r_sum1_5__9__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_14__10__q ;
wire Xd_0__inst_r_sum1_15__10__q ;
wire Xd_0__inst_r_sum1_12__10__q ;
wire Xd_0__inst_r_sum1_13__10__q ;
wire Xd_0__inst_r_sum1_10__10__q ;
wire Xd_0__inst_r_sum1_11__10__q ;
wire Xd_0__inst_r_sum1_8__10__q ;
wire Xd_0__inst_r_sum1_9__10__q ;
wire Xd_0__inst_r_sum1_6__10__q ;
wire Xd_0__inst_r_sum1_7__10__q ;
wire Xd_0__inst_r_sum1_4__10__q ;
wire Xd_0__inst_r_sum1_5__10__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_14__11__q ;
wire Xd_0__inst_r_sum1_15__11__q ;
wire Xd_0__inst_r_sum1_12__11__q ;
wire Xd_0__inst_r_sum1_13__11__q ;
wire Xd_0__inst_r_sum1_10__11__q ;
wire Xd_0__inst_r_sum1_11__11__q ;
wire Xd_0__inst_r_sum1_8__11__q ;
wire Xd_0__inst_r_sum1_9__11__q ;
wire Xd_0__inst_r_sum1_6__11__q ;
wire Xd_0__inst_r_sum1_7__11__q ;
wire Xd_0__inst_r_sum1_4__11__q ;
wire Xd_0__inst_r_sum1_5__11__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_14__12__q ;
wire Xd_0__inst_r_sum1_15__12__q ;
wire Xd_0__inst_r_sum1_12__12__q ;
wire Xd_0__inst_r_sum1_13__12__q ;
wire Xd_0__inst_r_sum1_10__12__q ;
wire Xd_0__inst_r_sum1_11__12__q ;
wire Xd_0__inst_r_sum1_8__12__q ;
wire Xd_0__inst_r_sum1_9__12__q ;
wire Xd_0__inst_r_sum1_6__12__q ;
wire Xd_0__inst_r_sum1_7__12__q ;
wire Xd_0__inst_r_sum1_4__12__q ;
wire Xd_0__inst_r_sum1_5__12__q ;
wire Xd_0__inst_r_sum1_2__12__q ;
wire Xd_0__inst_r_sum1_3__12__q ;
wire Xd_0__inst_r_sum1_0__12__q ;
wire Xd_0__inst_r_sum1_1__12__q ;
wire Xd_0__inst_r_sum1_14__13__q ;
wire Xd_0__inst_r_sum1_15__13__q ;
wire Xd_0__inst_r_sum1_12__13__q ;
wire Xd_0__inst_r_sum1_13__13__q ;
wire Xd_0__inst_r_sum1_10__13__q ;
wire Xd_0__inst_r_sum1_11__13__q ;
wire Xd_0__inst_r_sum1_8__13__q ;
wire Xd_0__inst_r_sum1_9__13__q ;
wire Xd_0__inst_r_sum1_6__13__q ;
wire Xd_0__inst_r_sum1_7__13__q ;
wire Xd_0__inst_r_sum1_4__13__q ;
wire Xd_0__inst_r_sum1_5__13__q ;
wire Xd_0__inst_r_sum1_2__13__q ;
wire Xd_0__inst_r_sum1_3__13__q ;
wire Xd_0__inst_r_sum1_0__13__q ;
wire Xd_0__inst_r_sum1_1__13__q ;
wire Xd_0__inst_r_sum1_14__14__q ;
wire Xd_0__inst_r_sum1_15__14__q ;
wire Xd_0__inst_r_sum1_12__14__q ;
wire Xd_0__inst_r_sum1_13__14__q ;
wire Xd_0__inst_r_sum1_10__14__q ;
wire Xd_0__inst_r_sum1_11__14__q ;
wire Xd_0__inst_r_sum1_8__14__q ;
wire Xd_0__inst_r_sum1_9__14__q ;
wire Xd_0__inst_r_sum1_6__14__q ;
wire Xd_0__inst_r_sum1_7__14__q ;
wire Xd_0__inst_r_sum1_4__14__q ;
wire Xd_0__inst_r_sum1_5__14__q ;
wire Xd_0__inst_r_sum1_2__14__q ;
wire Xd_0__inst_r_sum1_3__14__q ;
wire Xd_0__inst_r_sum1_0__14__q ;
wire Xd_0__inst_r_sum1_1__14__q ;
wire Xd_0__inst_r_sum1_14__15__q ;
wire Xd_0__inst_r_sum1_15__15__q ;
wire Xd_0__inst_r_sum1_12__15__q ;
wire Xd_0__inst_r_sum1_13__15__q ;
wire Xd_0__inst_r_sum1_10__15__q ;
wire Xd_0__inst_r_sum1_11__15__q ;
wire Xd_0__inst_r_sum1_8__15__q ;
wire Xd_0__inst_r_sum1_9__15__q ;
wire Xd_0__inst_r_sum1_6__15__q ;
wire Xd_0__inst_r_sum1_7__15__q ;
wire Xd_0__inst_r_sum1_4__15__q ;
wire Xd_0__inst_r_sum1_5__15__q ;
wire Xd_0__inst_r_sum1_2__15__q ;
wire Xd_0__inst_r_sum1_3__15__q ;
wire Xd_0__inst_r_sum1_0__15__q ;
wire Xd_0__inst_r_sum1_1__15__q ;
wire Xd_0__inst_r_sum1_14__16__q ;
wire Xd_0__inst_r_sum1_15__16__q ;
wire Xd_0__inst_r_sum1_12__16__q ;
wire Xd_0__inst_r_sum1_13__16__q ;
wire Xd_0__inst_r_sum1_10__16__q ;
wire Xd_0__inst_r_sum1_11__16__q ;
wire Xd_0__inst_r_sum1_8__16__q ;
wire Xd_0__inst_r_sum1_9__16__q ;
wire Xd_0__inst_r_sum1_6__16__q ;
wire Xd_0__inst_r_sum1_7__16__q ;
wire Xd_0__inst_r_sum1_4__16__q ;
wire Xd_0__inst_r_sum1_5__16__q ;
wire Xd_0__inst_r_sum1_2__16__q ;
wire Xd_0__inst_r_sum1_3__16__q ;
wire Xd_0__inst_r_sum1_0__16__q ;
wire Xd_0__inst_r_sum1_1__16__q ;
wire Xd_0__inst_r_sum1_14__17__q ;
wire Xd_0__inst_r_sum1_15__17__q ;
wire Xd_0__inst_r_sum1_12__17__q ;
wire Xd_0__inst_r_sum1_13__17__q ;
wire Xd_0__inst_r_sum1_10__17__q ;
wire Xd_0__inst_r_sum1_11__17__q ;
wire Xd_0__inst_r_sum1_8__17__q ;
wire Xd_0__inst_r_sum1_9__17__q ;
wire Xd_0__inst_r_sum1_6__17__q ;
wire Xd_0__inst_r_sum1_7__17__q ;
wire Xd_0__inst_r_sum1_4__17__q ;
wire Xd_0__inst_r_sum1_5__17__q ;
wire Xd_0__inst_r_sum1_2__17__q ;
wire Xd_0__inst_r_sum1_3__17__q ;
wire Xd_0__inst_r_sum1_0__17__q ;
wire Xd_0__inst_r_sum1_1__17__q ;
wire Xd_0__inst_r_sum1_14__18__q ;
wire Xd_0__inst_r_sum1_15__18__q ;
wire Xd_0__inst_r_sum1_12__18__q ;
wire Xd_0__inst_r_sum1_13__18__q ;
wire Xd_0__inst_r_sum1_10__18__q ;
wire Xd_0__inst_r_sum1_11__18__q ;
wire Xd_0__inst_r_sum1_8__18__q ;
wire Xd_0__inst_r_sum1_9__18__q ;
wire Xd_0__inst_r_sum1_6__18__q ;
wire Xd_0__inst_r_sum1_7__18__q ;
wire Xd_0__inst_r_sum1_4__18__q ;
wire Xd_0__inst_r_sum1_5__18__q ;
wire Xd_0__inst_r_sum1_2__18__q ;
wire Xd_0__inst_r_sum1_3__18__q ;
wire Xd_0__inst_r_sum1_0__18__q ;
wire Xd_0__inst_r_sum1_1__18__q ;
wire Xd_0__inst_r_sum1_14__19__q ;
wire Xd_0__inst_r_sum1_15__19__q ;
wire Xd_0__inst_r_sum1_12__19__q ;
wire Xd_0__inst_r_sum1_13__19__q ;
wire Xd_0__inst_r_sum1_10__19__q ;
wire Xd_0__inst_r_sum1_11__19__q ;
wire Xd_0__inst_r_sum1_8__19__q ;
wire Xd_0__inst_r_sum1_9__19__q ;
wire Xd_0__inst_r_sum1_6__19__q ;
wire Xd_0__inst_r_sum1_7__19__q ;
wire Xd_0__inst_r_sum1_4__19__q ;
wire Xd_0__inst_r_sum1_5__19__q ;
wire Xd_0__inst_r_sum1_2__19__q ;
wire Xd_0__inst_r_sum1_3__19__q ;
wire Xd_0__inst_r_sum1_0__19__q ;
wire Xd_0__inst_r_sum1_1__19__q ;
wire Xd_0__inst_r_sum1_14__20__q ;
wire Xd_0__inst_r_sum1_15__20__q ;
wire Xd_0__inst_r_sum1_12__20__q ;
wire Xd_0__inst_r_sum1_13__20__q ;
wire Xd_0__inst_r_sum1_10__20__q ;
wire Xd_0__inst_r_sum1_11__20__q ;
wire Xd_0__inst_r_sum1_8__20__q ;
wire Xd_0__inst_r_sum1_9__20__q ;
wire Xd_0__inst_r_sum1_6__20__q ;
wire Xd_0__inst_r_sum1_7__20__q ;
wire Xd_0__inst_r_sum1_4__20__q ;
wire Xd_0__inst_r_sum1_5__20__q ;
wire Xd_0__inst_r_sum1_2__20__q ;
wire Xd_0__inst_r_sum1_3__20__q ;
wire Xd_0__inst_r_sum1_0__20__q ;
wire Xd_0__inst_r_sum1_1__20__q ;
wire Xd_0__inst_r_sum1_14__21__q ;
wire Xd_0__inst_r_sum1_15__21__q ;
wire Xd_0__inst_r_sum1_12__21__q ;
wire Xd_0__inst_r_sum1_13__21__q ;
wire Xd_0__inst_r_sum1_10__21__q ;
wire Xd_0__inst_r_sum1_11__21__q ;
wire Xd_0__inst_r_sum1_8__21__q ;
wire Xd_0__inst_r_sum1_9__21__q ;
wire Xd_0__inst_r_sum1_6__21__q ;
wire Xd_0__inst_r_sum1_7__21__q ;
wire Xd_0__inst_r_sum1_4__21__q ;
wire Xd_0__inst_r_sum1_5__21__q ;
wire Xd_0__inst_r_sum1_2__21__q ;
wire Xd_0__inst_r_sum1_3__21__q ;
wire Xd_0__inst_r_sum1_0__21__q ;
wire Xd_0__inst_r_sum1_1__21__q ;
wire Xd_0__inst_r_sum1_14__22__q ;
wire Xd_0__inst_r_sum1_15__22__q ;
wire Xd_0__inst_r_sum1_12__22__q ;
wire Xd_0__inst_r_sum1_13__22__q ;
wire Xd_0__inst_r_sum1_10__22__q ;
wire Xd_0__inst_r_sum1_11__22__q ;
wire Xd_0__inst_r_sum1_8__22__q ;
wire Xd_0__inst_r_sum1_9__22__q ;
wire Xd_0__inst_r_sum1_6__22__q ;
wire Xd_0__inst_r_sum1_7__22__q ;
wire Xd_0__inst_r_sum1_4__22__q ;
wire Xd_0__inst_r_sum1_5__22__q ;
wire Xd_0__inst_r_sum1_2__22__q ;
wire Xd_0__inst_r_sum1_3__22__q ;
wire Xd_0__inst_r_sum1_0__22__q ;
wire Xd_0__inst_r_sum1_1__22__q ;
wire Xd_0__inst_r_sum1_14__23__q ;
wire Xd_0__inst_r_sum1_15__23__q ;
wire Xd_0__inst_r_sum1_12__23__q ;
wire Xd_0__inst_r_sum1_13__23__q ;
wire Xd_0__inst_r_sum1_10__23__q ;
wire Xd_0__inst_r_sum1_11__23__q ;
wire Xd_0__inst_r_sum1_8__23__q ;
wire Xd_0__inst_r_sum1_9__23__q ;
wire Xd_0__inst_r_sum1_6__23__q ;
wire Xd_0__inst_r_sum1_7__23__q ;
wire Xd_0__inst_r_sum1_4__23__q ;
wire Xd_0__inst_r_sum1_5__23__q ;
wire Xd_0__inst_r_sum1_2__23__q ;
wire Xd_0__inst_r_sum1_3__23__q ;
wire Xd_0__inst_r_sum1_0__23__q ;
wire Xd_0__inst_r_sum1_1__23__q ;
wire Xd_0__inst_product_31__0__q ;
wire Xd_0__inst_product_30__0__q ;
wire Xd_0__inst_product_29__0__q ;
wire Xd_0__inst_product_28__0__q ;
wire Xd_0__inst_product_27__0__q ;
wire Xd_0__inst_product_26__0__q ;
wire Xd_0__inst_product_25__0__q ;
wire Xd_0__inst_product_24__0__q ;
wire Xd_0__inst_product_23__0__q ;
wire Xd_0__inst_product_22__0__q ;
wire Xd_0__inst_product_21__0__q ;
wire Xd_0__inst_product_20__0__q ;
wire Xd_0__inst_product_19__0__q ;
wire Xd_0__inst_product_18__0__q ;
wire Xd_0__inst_product_17__0__q ;
wire Xd_0__inst_product_16__0__q ;
wire Xd_0__inst_product_15__0__q ;
wire Xd_0__inst_product_14__0__q ;
wire Xd_0__inst_product_13__0__q ;
wire Xd_0__inst_product_12__0__q ;
wire Xd_0__inst_product_11__0__q ;
wire Xd_0__inst_product_10__0__q ;
wire Xd_0__inst_product_9__0__q ;
wire Xd_0__inst_product_8__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_29__1__q ;
wire Xd_0__inst_product_28__1__q ;
wire Xd_0__inst_product_31__1__q ;
wire Xd_0__inst_product_30__1__q ;
wire Xd_0__inst_product_25__1__q ;
wire Xd_0__inst_product_24__1__q ;
wire Xd_0__inst_product_27__1__q ;
wire Xd_0__inst_product_26__1__q ;
wire Xd_0__inst_product_21__1__q ;
wire Xd_0__inst_product_20__1__q ;
wire Xd_0__inst_product_23__1__q ;
wire Xd_0__inst_product_22__1__q ;
wire Xd_0__inst_product_17__1__q ;
wire Xd_0__inst_product_16__1__q ;
wire Xd_0__inst_product_19__1__q ;
wire Xd_0__inst_product_18__1__q ;
wire Xd_0__inst_product_13__1__q ;
wire Xd_0__inst_product_12__1__q ;
wire Xd_0__inst_product_15__1__q ;
wire Xd_0__inst_product_14__1__q ;
wire Xd_0__inst_product_9__1__q ;
wire Xd_0__inst_product_8__1__q ;
wire Xd_0__inst_product_11__1__q ;
wire Xd_0__inst_product_10__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_29__2__q ;
wire Xd_0__inst_product_28__2__q ;
wire Xd_0__inst_product_31__2__q ;
wire Xd_0__inst_product_30__2__q ;
wire Xd_0__inst_product_25__2__q ;
wire Xd_0__inst_product_24__2__q ;
wire Xd_0__inst_product_27__2__q ;
wire Xd_0__inst_product_26__2__q ;
wire Xd_0__inst_product_21__2__q ;
wire Xd_0__inst_product_20__2__q ;
wire Xd_0__inst_product_23__2__q ;
wire Xd_0__inst_product_22__2__q ;
wire Xd_0__inst_product_17__2__q ;
wire Xd_0__inst_product_16__2__q ;
wire Xd_0__inst_product_19__2__q ;
wire Xd_0__inst_product_18__2__q ;
wire Xd_0__inst_product_13__2__q ;
wire Xd_0__inst_product_12__2__q ;
wire Xd_0__inst_product_15__2__q ;
wire Xd_0__inst_product_14__2__q ;
wire Xd_0__inst_product_9__2__q ;
wire Xd_0__inst_product_8__2__q ;
wire Xd_0__inst_product_11__2__q ;
wire Xd_0__inst_product_10__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_29__3__q ;
wire Xd_0__inst_product_28__3__q ;
wire Xd_0__inst_product_31__3__q ;
wire Xd_0__inst_product_30__3__q ;
wire Xd_0__inst_product_25__3__q ;
wire Xd_0__inst_product_24__3__q ;
wire Xd_0__inst_product_27__3__q ;
wire Xd_0__inst_product_26__3__q ;
wire Xd_0__inst_product_21__3__q ;
wire Xd_0__inst_product_20__3__q ;
wire Xd_0__inst_product_23__3__q ;
wire Xd_0__inst_product_22__3__q ;
wire Xd_0__inst_product_17__3__q ;
wire Xd_0__inst_product_16__3__q ;
wire Xd_0__inst_product_19__3__q ;
wire Xd_0__inst_product_18__3__q ;
wire Xd_0__inst_product_13__3__q ;
wire Xd_0__inst_product_12__3__q ;
wire Xd_0__inst_product_15__3__q ;
wire Xd_0__inst_product_14__3__q ;
wire Xd_0__inst_product_9__3__q ;
wire Xd_0__inst_product_8__3__q ;
wire Xd_0__inst_product_11__3__q ;
wire Xd_0__inst_product_10__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_29__4__q ;
wire Xd_0__inst_product_28__4__q ;
wire Xd_0__inst_product_31__4__q ;
wire Xd_0__inst_product_30__4__q ;
wire Xd_0__inst_product_25__4__q ;
wire Xd_0__inst_product_24__4__q ;
wire Xd_0__inst_product_27__4__q ;
wire Xd_0__inst_product_26__4__q ;
wire Xd_0__inst_product_21__4__q ;
wire Xd_0__inst_product_20__4__q ;
wire Xd_0__inst_product_23__4__q ;
wire Xd_0__inst_product_22__4__q ;
wire Xd_0__inst_product_17__4__q ;
wire Xd_0__inst_product_16__4__q ;
wire Xd_0__inst_product_19__4__q ;
wire Xd_0__inst_product_18__4__q ;
wire Xd_0__inst_product_13__4__q ;
wire Xd_0__inst_product_12__4__q ;
wire Xd_0__inst_product_15__4__q ;
wire Xd_0__inst_product_14__4__q ;
wire Xd_0__inst_product_9__4__q ;
wire Xd_0__inst_product_8__4__q ;
wire Xd_0__inst_product_11__4__q ;
wire Xd_0__inst_product_10__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_29__5__q ;
wire Xd_0__inst_product_28__5__q ;
wire Xd_0__inst_product_31__5__q ;
wire Xd_0__inst_product_30__5__q ;
wire Xd_0__inst_product_25__5__q ;
wire Xd_0__inst_product_24__5__q ;
wire Xd_0__inst_product_27__5__q ;
wire Xd_0__inst_product_26__5__q ;
wire Xd_0__inst_product_21__5__q ;
wire Xd_0__inst_product_20__5__q ;
wire Xd_0__inst_product_23__5__q ;
wire Xd_0__inst_product_22__5__q ;
wire Xd_0__inst_product_17__5__q ;
wire Xd_0__inst_product_16__5__q ;
wire Xd_0__inst_product_19__5__q ;
wire Xd_0__inst_product_18__5__q ;
wire Xd_0__inst_product_13__5__q ;
wire Xd_0__inst_product_12__5__q ;
wire Xd_0__inst_product_15__5__q ;
wire Xd_0__inst_product_14__5__q ;
wire Xd_0__inst_product_9__5__q ;
wire Xd_0__inst_product_8__5__q ;
wire Xd_0__inst_product_11__5__q ;
wire Xd_0__inst_product_10__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_29__6__q ;
wire Xd_0__inst_product_28__6__q ;
wire Xd_0__inst_product_31__6__q ;
wire Xd_0__inst_product_30__6__q ;
wire Xd_0__inst_product_25__6__q ;
wire Xd_0__inst_product_24__6__q ;
wire Xd_0__inst_product_27__6__q ;
wire Xd_0__inst_product_26__6__q ;
wire Xd_0__inst_product_21__6__q ;
wire Xd_0__inst_product_20__6__q ;
wire Xd_0__inst_product_23__6__q ;
wire Xd_0__inst_product_22__6__q ;
wire Xd_0__inst_product_17__6__q ;
wire Xd_0__inst_product_16__6__q ;
wire Xd_0__inst_product_19__6__q ;
wire Xd_0__inst_product_18__6__q ;
wire Xd_0__inst_product_13__6__q ;
wire Xd_0__inst_product_12__6__q ;
wire Xd_0__inst_product_15__6__q ;
wire Xd_0__inst_product_14__6__q ;
wire Xd_0__inst_product_9__6__q ;
wire Xd_0__inst_product_8__6__q ;
wire Xd_0__inst_product_11__6__q ;
wire Xd_0__inst_product_10__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_29__7__q ;
wire Xd_0__inst_product_28__7__q ;
wire Xd_0__inst_product_31__7__q ;
wire Xd_0__inst_product_30__7__q ;
wire Xd_0__inst_product_25__7__q ;
wire Xd_0__inst_product_24__7__q ;
wire Xd_0__inst_product_27__7__q ;
wire Xd_0__inst_product_26__7__q ;
wire Xd_0__inst_product_21__7__q ;
wire Xd_0__inst_product_20__7__q ;
wire Xd_0__inst_product_23__7__q ;
wire Xd_0__inst_product_22__7__q ;
wire Xd_0__inst_product_17__7__q ;
wire Xd_0__inst_product_16__7__q ;
wire Xd_0__inst_product_19__7__q ;
wire Xd_0__inst_product_18__7__q ;
wire Xd_0__inst_product_13__7__q ;
wire Xd_0__inst_product_12__7__q ;
wire Xd_0__inst_product_15__7__q ;
wire Xd_0__inst_product_14__7__q ;
wire Xd_0__inst_product_9__7__q ;
wire Xd_0__inst_product_8__7__q ;
wire Xd_0__inst_product_11__7__q ;
wire Xd_0__inst_product_10__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_29__8__q ;
wire Xd_0__inst_product_28__8__q ;
wire Xd_0__inst_product_31__8__q ;
wire Xd_0__inst_product_30__8__q ;
wire Xd_0__inst_product_25__8__q ;
wire Xd_0__inst_product_24__8__q ;
wire Xd_0__inst_product_27__8__q ;
wire Xd_0__inst_product_26__8__q ;
wire Xd_0__inst_product_21__8__q ;
wire Xd_0__inst_product_20__8__q ;
wire Xd_0__inst_product_23__8__q ;
wire Xd_0__inst_product_22__8__q ;
wire Xd_0__inst_product_17__8__q ;
wire Xd_0__inst_product_16__8__q ;
wire Xd_0__inst_product_19__8__q ;
wire Xd_0__inst_product_18__8__q ;
wire Xd_0__inst_product_13__8__q ;
wire Xd_0__inst_product_12__8__q ;
wire Xd_0__inst_product_15__8__q ;
wire Xd_0__inst_product_14__8__q ;
wire Xd_0__inst_product_9__8__q ;
wire Xd_0__inst_product_8__8__q ;
wire Xd_0__inst_product_11__8__q ;
wire Xd_0__inst_product_10__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_29__9__q ;
wire Xd_0__inst_product_28__9__q ;
wire Xd_0__inst_product_31__9__q ;
wire Xd_0__inst_product_30__9__q ;
wire Xd_0__inst_product_25__9__q ;
wire Xd_0__inst_product_24__9__q ;
wire Xd_0__inst_product_27__9__q ;
wire Xd_0__inst_product_26__9__q ;
wire Xd_0__inst_product_21__9__q ;
wire Xd_0__inst_product_20__9__q ;
wire Xd_0__inst_product_23__9__q ;
wire Xd_0__inst_product_22__9__q ;
wire Xd_0__inst_product_17__9__q ;
wire Xd_0__inst_product_16__9__q ;
wire Xd_0__inst_product_19__9__q ;
wire Xd_0__inst_product_18__9__q ;
wire Xd_0__inst_product_13__9__q ;
wire Xd_0__inst_product_12__9__q ;
wire Xd_0__inst_product_15__9__q ;
wire Xd_0__inst_product_14__9__q ;
wire Xd_0__inst_product_9__9__q ;
wire Xd_0__inst_product_8__9__q ;
wire Xd_0__inst_product_11__9__q ;
wire Xd_0__inst_product_10__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_29__10__q ;
wire Xd_0__inst_product_28__10__q ;
wire Xd_0__inst_product_31__10__q ;
wire Xd_0__inst_product_30__10__q ;
wire Xd_0__inst_product_25__10__q ;
wire Xd_0__inst_product_24__10__q ;
wire Xd_0__inst_product_27__10__q ;
wire Xd_0__inst_product_26__10__q ;
wire Xd_0__inst_product_21__10__q ;
wire Xd_0__inst_product_20__10__q ;
wire Xd_0__inst_product_23__10__q ;
wire Xd_0__inst_product_22__10__q ;
wire Xd_0__inst_product_17__10__q ;
wire Xd_0__inst_product_16__10__q ;
wire Xd_0__inst_product_19__10__q ;
wire Xd_0__inst_product_18__10__q ;
wire Xd_0__inst_product_13__10__q ;
wire Xd_0__inst_product_12__10__q ;
wire Xd_0__inst_product_15__10__q ;
wire Xd_0__inst_product_14__10__q ;
wire Xd_0__inst_product_9__10__q ;
wire Xd_0__inst_product_8__10__q ;
wire Xd_0__inst_product_11__10__q ;
wire Xd_0__inst_product_10__10__q ;
wire Xd_0__inst_product_5__10__q ;
wire Xd_0__inst_product_4__10__q ;
wire Xd_0__inst_product_7__10__q ;
wire Xd_0__inst_product_6__10__q ;
wire Xd_0__inst_product_1__10__q ;
wire Xd_0__inst_product_0__10__q ;
wire Xd_0__inst_product_3__10__q ;
wire Xd_0__inst_product_2__10__q ;
wire Xd_0__inst_product_29__11__q ;
wire Xd_0__inst_product_28__11__q ;
wire Xd_0__inst_product_31__11__q ;
wire Xd_0__inst_product_30__11__q ;
wire Xd_0__inst_product_25__11__q ;
wire Xd_0__inst_product_24__11__q ;
wire Xd_0__inst_product_27__11__q ;
wire Xd_0__inst_product_26__11__q ;
wire Xd_0__inst_product_21__11__q ;
wire Xd_0__inst_product_20__11__q ;
wire Xd_0__inst_product_23__11__q ;
wire Xd_0__inst_product_22__11__q ;
wire Xd_0__inst_product_17__11__q ;
wire Xd_0__inst_product_16__11__q ;
wire Xd_0__inst_product_19__11__q ;
wire Xd_0__inst_product_18__11__q ;
wire Xd_0__inst_product_13__11__q ;
wire Xd_0__inst_product_12__11__q ;
wire Xd_0__inst_product_15__11__q ;
wire Xd_0__inst_product_14__11__q ;
wire Xd_0__inst_product_9__11__q ;
wire Xd_0__inst_product_8__11__q ;
wire Xd_0__inst_product_11__11__q ;
wire Xd_0__inst_product_10__11__q ;
wire Xd_0__inst_product_5__11__q ;
wire Xd_0__inst_product_4__11__q ;
wire Xd_0__inst_product_7__11__q ;
wire Xd_0__inst_product_6__11__q ;
wire Xd_0__inst_product_1__11__q ;
wire Xd_0__inst_product_0__11__q ;
wire Xd_0__inst_product_3__11__q ;
wire Xd_0__inst_product_2__11__q ;
wire Xd_0__inst_product_29__12__q ;
wire Xd_0__inst_product_28__12__q ;
wire Xd_0__inst_product_31__12__q ;
wire Xd_0__inst_product_30__12__q ;
wire Xd_0__inst_product_25__12__q ;
wire Xd_0__inst_product_24__12__q ;
wire Xd_0__inst_product_27__12__q ;
wire Xd_0__inst_product_26__12__q ;
wire Xd_0__inst_product_21__12__q ;
wire Xd_0__inst_product_20__12__q ;
wire Xd_0__inst_product_23__12__q ;
wire Xd_0__inst_product_22__12__q ;
wire Xd_0__inst_product_17__12__q ;
wire Xd_0__inst_product_16__12__q ;
wire Xd_0__inst_product_19__12__q ;
wire Xd_0__inst_product_18__12__q ;
wire Xd_0__inst_product_13__12__q ;
wire Xd_0__inst_product_12__12__q ;
wire Xd_0__inst_product_15__12__q ;
wire Xd_0__inst_product_14__12__q ;
wire Xd_0__inst_product_9__12__q ;
wire Xd_0__inst_product_8__12__q ;
wire Xd_0__inst_product_11__12__q ;
wire Xd_0__inst_product_10__12__q ;
wire Xd_0__inst_product_5__12__q ;
wire Xd_0__inst_product_4__12__q ;
wire Xd_0__inst_product_7__12__q ;
wire Xd_0__inst_product_6__12__q ;
wire Xd_0__inst_product_1__12__q ;
wire Xd_0__inst_product_0__12__q ;
wire Xd_0__inst_product_3__12__q ;
wire Xd_0__inst_product_2__12__q ;
wire Xd_0__inst_product_29__13__q ;
wire Xd_0__inst_product_28__13__q ;
wire Xd_0__inst_product_31__13__q ;
wire Xd_0__inst_product_30__13__q ;
wire Xd_0__inst_product_25__13__q ;
wire Xd_0__inst_product_24__13__q ;
wire Xd_0__inst_product_27__13__q ;
wire Xd_0__inst_product_26__13__q ;
wire Xd_0__inst_product_21__13__q ;
wire Xd_0__inst_product_20__13__q ;
wire Xd_0__inst_product_23__13__q ;
wire Xd_0__inst_product_22__13__q ;
wire Xd_0__inst_product_17__13__q ;
wire Xd_0__inst_product_16__13__q ;
wire Xd_0__inst_product_19__13__q ;
wire Xd_0__inst_product_18__13__q ;
wire Xd_0__inst_product_13__13__q ;
wire Xd_0__inst_product_12__13__q ;
wire Xd_0__inst_product_15__13__q ;
wire Xd_0__inst_product_14__13__q ;
wire Xd_0__inst_product_9__13__q ;
wire Xd_0__inst_product_8__13__q ;
wire Xd_0__inst_product_11__13__q ;
wire Xd_0__inst_product_10__13__q ;
wire Xd_0__inst_product_5__13__q ;
wire Xd_0__inst_product_4__13__q ;
wire Xd_0__inst_product_7__13__q ;
wire Xd_0__inst_product_6__13__q ;
wire Xd_0__inst_product_1__13__q ;
wire Xd_0__inst_product_0__13__q ;
wire Xd_0__inst_product_3__13__q ;
wire Xd_0__inst_product_2__13__q ;
wire Xd_0__inst_product_29__14__q ;
wire Xd_0__inst_product_28__14__q ;
wire Xd_0__inst_product_31__14__q ;
wire Xd_0__inst_product_30__14__q ;
wire Xd_0__inst_product_25__14__q ;
wire Xd_0__inst_product_24__14__q ;
wire Xd_0__inst_product_27__14__q ;
wire Xd_0__inst_product_26__14__q ;
wire Xd_0__inst_product_21__14__q ;
wire Xd_0__inst_product_20__14__q ;
wire Xd_0__inst_product_23__14__q ;
wire Xd_0__inst_product_22__14__q ;
wire Xd_0__inst_product_17__14__q ;
wire Xd_0__inst_product_16__14__q ;
wire Xd_0__inst_product_19__14__q ;
wire Xd_0__inst_product_18__14__q ;
wire Xd_0__inst_product_13__14__q ;
wire Xd_0__inst_product_12__14__q ;
wire Xd_0__inst_product_15__14__q ;
wire Xd_0__inst_product_14__14__q ;
wire Xd_0__inst_product_9__14__q ;
wire Xd_0__inst_product_8__14__q ;
wire Xd_0__inst_product_11__14__q ;
wire Xd_0__inst_product_10__14__q ;
wire Xd_0__inst_product_5__14__q ;
wire Xd_0__inst_product_4__14__q ;
wire Xd_0__inst_product_7__14__q ;
wire Xd_0__inst_product_6__14__q ;
wire Xd_0__inst_product_1__14__q ;
wire Xd_0__inst_product_0__14__q ;
wire Xd_0__inst_product_3__14__q ;
wire Xd_0__inst_product_2__14__q ;
wire Xd_0__inst_product_29__15__q ;
wire Xd_0__inst_product_28__15__q ;
wire Xd_0__inst_product_31__15__q ;
wire Xd_0__inst_product_30__15__q ;
wire Xd_0__inst_product_25__15__q ;
wire Xd_0__inst_product_24__15__q ;
wire Xd_0__inst_product_27__15__q ;
wire Xd_0__inst_product_26__15__q ;
wire Xd_0__inst_product_21__15__q ;
wire Xd_0__inst_product_20__15__q ;
wire Xd_0__inst_product_23__15__q ;
wire Xd_0__inst_product_22__15__q ;
wire Xd_0__inst_product_17__15__q ;
wire Xd_0__inst_product_16__15__q ;
wire Xd_0__inst_product_19__15__q ;
wire Xd_0__inst_product_18__15__q ;
wire Xd_0__inst_product_13__15__q ;
wire Xd_0__inst_product_12__15__q ;
wire Xd_0__inst_product_15__15__q ;
wire Xd_0__inst_product_14__15__q ;
wire Xd_0__inst_product_9__15__q ;
wire Xd_0__inst_product_8__15__q ;
wire Xd_0__inst_product_11__15__q ;
wire Xd_0__inst_product_10__15__q ;
wire Xd_0__inst_product_5__15__q ;
wire Xd_0__inst_product_4__15__q ;
wire Xd_0__inst_product_7__15__q ;
wire Xd_0__inst_product_6__15__q ;
wire Xd_0__inst_product_1__15__q ;
wire Xd_0__inst_product_0__15__q ;
wire Xd_0__inst_product_3__15__q ;
wire Xd_0__inst_product_2__15__q ;
wire Xd_0__inst_product_29__16__q ;
wire Xd_0__inst_product_28__16__q ;
wire Xd_0__inst_product_31__16__q ;
wire Xd_0__inst_product_30__16__q ;
wire Xd_0__inst_product_25__16__q ;
wire Xd_0__inst_product_24__16__q ;
wire Xd_0__inst_product_27__16__q ;
wire Xd_0__inst_product_26__16__q ;
wire Xd_0__inst_product_21__16__q ;
wire Xd_0__inst_product_20__16__q ;
wire Xd_0__inst_product_23__16__q ;
wire Xd_0__inst_product_22__16__q ;
wire Xd_0__inst_product_17__16__q ;
wire Xd_0__inst_product_16__16__q ;
wire Xd_0__inst_product_19__16__q ;
wire Xd_0__inst_product_18__16__q ;
wire Xd_0__inst_product_13__16__q ;
wire Xd_0__inst_product_12__16__q ;
wire Xd_0__inst_product_15__16__q ;
wire Xd_0__inst_product_14__16__q ;
wire Xd_0__inst_product_9__16__q ;
wire Xd_0__inst_product_8__16__q ;
wire Xd_0__inst_product_11__16__q ;
wire Xd_0__inst_product_10__16__q ;
wire Xd_0__inst_product_5__16__q ;
wire Xd_0__inst_product_4__16__q ;
wire Xd_0__inst_product_7__16__q ;
wire Xd_0__inst_product_6__16__q ;
wire Xd_0__inst_product_1__16__q ;
wire Xd_0__inst_product_0__16__q ;
wire Xd_0__inst_product_3__16__q ;
wire Xd_0__inst_product_2__16__q ;
wire Xd_0__inst_product_29__17__q ;
wire Xd_0__inst_product_28__17__q ;
wire Xd_0__inst_product_31__17__q ;
wire Xd_0__inst_product_30__17__q ;
wire Xd_0__inst_product_25__17__q ;
wire Xd_0__inst_product_24__17__q ;
wire Xd_0__inst_product_27__17__q ;
wire Xd_0__inst_product_26__17__q ;
wire Xd_0__inst_product_21__17__q ;
wire Xd_0__inst_product_20__17__q ;
wire Xd_0__inst_product_23__17__q ;
wire Xd_0__inst_product_22__17__q ;
wire Xd_0__inst_product_17__17__q ;
wire Xd_0__inst_product_16__17__q ;
wire Xd_0__inst_product_19__17__q ;
wire Xd_0__inst_product_18__17__q ;
wire Xd_0__inst_product_13__17__q ;
wire Xd_0__inst_product_12__17__q ;
wire Xd_0__inst_product_15__17__q ;
wire Xd_0__inst_product_14__17__q ;
wire Xd_0__inst_product_9__17__q ;
wire Xd_0__inst_product_8__17__q ;
wire Xd_0__inst_product_11__17__q ;
wire Xd_0__inst_product_10__17__q ;
wire Xd_0__inst_product_5__17__q ;
wire Xd_0__inst_product_4__17__q ;
wire Xd_0__inst_product_7__17__q ;
wire Xd_0__inst_product_6__17__q ;
wire Xd_0__inst_product_1__17__q ;
wire Xd_0__inst_product_0__17__q ;
wire Xd_0__inst_product_3__17__q ;
wire Xd_0__inst_product_2__17__q ;
wire Xd_0__inst_product_29__18__q ;
wire Xd_0__inst_product_28__18__q ;
wire Xd_0__inst_product_31__18__q ;
wire Xd_0__inst_product_30__18__q ;
wire Xd_0__inst_product_25__18__q ;
wire Xd_0__inst_product_24__18__q ;
wire Xd_0__inst_product_27__18__q ;
wire Xd_0__inst_product_26__18__q ;
wire Xd_0__inst_product_21__18__q ;
wire Xd_0__inst_product_20__18__q ;
wire Xd_0__inst_product_23__18__q ;
wire Xd_0__inst_product_22__18__q ;
wire Xd_0__inst_product_17__18__q ;
wire Xd_0__inst_product_16__18__q ;
wire Xd_0__inst_product_19__18__q ;
wire Xd_0__inst_product_18__18__q ;
wire Xd_0__inst_product_13__18__q ;
wire Xd_0__inst_product_12__18__q ;
wire Xd_0__inst_product_15__18__q ;
wire Xd_0__inst_product_14__18__q ;
wire Xd_0__inst_product_9__18__q ;
wire Xd_0__inst_product_8__18__q ;
wire Xd_0__inst_product_11__18__q ;
wire Xd_0__inst_product_10__18__q ;
wire Xd_0__inst_product_5__18__q ;
wire Xd_0__inst_product_4__18__q ;
wire Xd_0__inst_product_7__18__q ;
wire Xd_0__inst_product_6__18__q ;
wire Xd_0__inst_product_1__18__q ;
wire Xd_0__inst_product_0__18__q ;
wire Xd_0__inst_product_3__18__q ;
wire Xd_0__inst_product_2__18__q ;
wire Xd_0__inst_product_29__19__q ;
wire Xd_0__inst_product_28__19__q ;
wire Xd_0__inst_product_31__19__q ;
wire Xd_0__inst_product_30__19__q ;
wire Xd_0__inst_product_25__19__q ;
wire Xd_0__inst_product_24__19__q ;
wire Xd_0__inst_product_27__19__q ;
wire Xd_0__inst_product_26__19__q ;
wire Xd_0__inst_product_21__19__q ;
wire Xd_0__inst_product_20__19__q ;
wire Xd_0__inst_product_23__19__q ;
wire Xd_0__inst_product_22__19__q ;
wire Xd_0__inst_product_17__19__q ;
wire Xd_0__inst_product_16__19__q ;
wire Xd_0__inst_product_19__19__q ;
wire Xd_0__inst_product_18__19__q ;
wire Xd_0__inst_product_13__19__q ;
wire Xd_0__inst_product_12__19__q ;
wire Xd_0__inst_product_15__19__q ;
wire Xd_0__inst_product_14__19__q ;
wire Xd_0__inst_product_9__19__q ;
wire Xd_0__inst_product_8__19__q ;
wire Xd_0__inst_product_11__19__q ;
wire Xd_0__inst_product_10__19__q ;
wire Xd_0__inst_product_5__19__q ;
wire Xd_0__inst_product_4__19__q ;
wire Xd_0__inst_product_7__19__q ;
wire Xd_0__inst_product_6__19__q ;
wire Xd_0__inst_product_1__19__q ;
wire Xd_0__inst_product_0__19__q ;
wire Xd_0__inst_product_3__19__q ;
wire Xd_0__inst_product_2__19__q ;
wire Xd_0__inst_product_29__20__q ;
wire Xd_0__inst_product_28__20__q ;
wire Xd_0__inst_product_31__20__q ;
wire Xd_0__inst_product_30__20__q ;
wire Xd_0__inst_product_25__20__q ;
wire Xd_0__inst_product_24__20__q ;
wire Xd_0__inst_product_27__20__q ;
wire Xd_0__inst_product_26__20__q ;
wire Xd_0__inst_product_21__20__q ;
wire Xd_0__inst_product_20__20__q ;
wire Xd_0__inst_product_23__20__q ;
wire Xd_0__inst_product_22__20__q ;
wire Xd_0__inst_product_17__20__q ;
wire Xd_0__inst_product_16__20__q ;
wire Xd_0__inst_product_19__20__q ;
wire Xd_0__inst_product_18__20__q ;
wire Xd_0__inst_product_13__20__q ;
wire Xd_0__inst_product_12__20__q ;
wire Xd_0__inst_product_15__20__q ;
wire Xd_0__inst_product_14__20__q ;
wire Xd_0__inst_product_9__20__q ;
wire Xd_0__inst_product_8__20__q ;
wire Xd_0__inst_product_11__20__q ;
wire Xd_0__inst_product_10__20__q ;
wire Xd_0__inst_product_5__20__q ;
wire Xd_0__inst_product_4__20__q ;
wire Xd_0__inst_product_7__20__q ;
wire Xd_0__inst_product_6__20__q ;
wire Xd_0__inst_product_1__20__q ;
wire Xd_0__inst_product_0__20__q ;
wire Xd_0__inst_product_3__20__q ;
wire Xd_0__inst_product_2__20__q ;
wire Xd_0__inst_product_29__21__q ;
wire Xd_0__inst_product_28__21__q ;
wire Xd_0__inst_product_31__21__q ;
wire Xd_0__inst_product_30__21__q ;
wire Xd_0__inst_product_25__21__q ;
wire Xd_0__inst_product_24__21__q ;
wire Xd_0__inst_product_27__21__q ;
wire Xd_0__inst_product_26__21__q ;
wire Xd_0__inst_product_21__21__q ;
wire Xd_0__inst_product_20__21__q ;
wire Xd_0__inst_product_23__21__q ;
wire Xd_0__inst_product_22__21__q ;
wire Xd_0__inst_product_17__21__q ;
wire Xd_0__inst_product_16__21__q ;
wire Xd_0__inst_product_19__21__q ;
wire Xd_0__inst_product_18__21__q ;
wire Xd_0__inst_product_13__21__q ;
wire Xd_0__inst_product_12__21__q ;
wire Xd_0__inst_product_15__21__q ;
wire Xd_0__inst_product_14__21__q ;
wire Xd_0__inst_product_9__21__q ;
wire Xd_0__inst_product_8__21__q ;
wire Xd_0__inst_product_11__21__q ;
wire Xd_0__inst_product_10__21__q ;
wire Xd_0__inst_product_5__21__q ;
wire Xd_0__inst_product_4__21__q ;
wire Xd_0__inst_product_7__21__q ;
wire Xd_0__inst_product_6__21__q ;
wire Xd_0__inst_product_1__21__q ;
wire Xd_0__inst_product_0__21__q ;
wire Xd_0__inst_product_3__21__q ;
wire Xd_0__inst_product_2__21__q ;
wire Xd_0__inst_product1_31__0__q ;
wire Xd_0__inst_product1_30__0__q ;
wire Xd_0__inst_product1_29__0__q ;
wire Xd_0__inst_product1_28__0__q ;
wire Xd_0__inst_product1_27__0__q ;
wire Xd_0__inst_product1_26__0__q ;
wire Xd_0__inst_product1_25__0__q ;
wire Xd_0__inst_product1_24__0__q ;
wire Xd_0__inst_product1_23__0__q ;
wire Xd_0__inst_product1_22__0__q ;
wire Xd_0__inst_product1_21__0__q ;
wire Xd_0__inst_product1_20__0__q ;
wire Xd_0__inst_product1_19__0__q ;
wire Xd_0__inst_product1_18__0__q ;
wire Xd_0__inst_product1_17__0__q ;
wire Xd_0__inst_product1_16__0__q ;
wire Xd_0__inst_product1_15__0__q ;
wire Xd_0__inst_product1_14__0__q ;
wire Xd_0__inst_product1_13__0__q ;
wire Xd_0__inst_product1_12__0__q ;
wire Xd_0__inst_product1_11__0__q ;
wire Xd_0__inst_product1_10__0__q ;
wire Xd_0__inst_product1_9__0__q ;
wire Xd_0__inst_product1_8__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_29__1__q ;
wire Xd_0__inst_product1_28__1__q ;
wire Xd_0__inst_product1_31__1__q ;
wire Xd_0__inst_product1_30__1__q ;
wire Xd_0__inst_product1_25__1__q ;
wire Xd_0__inst_product1_24__1__q ;
wire Xd_0__inst_product1_27__1__q ;
wire Xd_0__inst_product1_26__1__q ;
wire Xd_0__inst_product1_21__1__q ;
wire Xd_0__inst_product1_20__1__q ;
wire Xd_0__inst_product1_23__1__q ;
wire Xd_0__inst_product1_22__1__q ;
wire Xd_0__inst_product1_17__1__q ;
wire Xd_0__inst_product1_16__1__q ;
wire Xd_0__inst_product1_19__1__q ;
wire Xd_0__inst_product1_18__1__q ;
wire Xd_0__inst_product1_13__1__q ;
wire Xd_0__inst_product1_12__1__q ;
wire Xd_0__inst_product1_15__1__q ;
wire Xd_0__inst_product1_14__1__q ;
wire Xd_0__inst_product1_9__1__q ;
wire Xd_0__inst_product1_8__1__q ;
wire Xd_0__inst_product1_11__1__q ;
wire Xd_0__inst_product1_10__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_29__2__q ;
wire Xd_0__inst_product1_28__2__q ;
wire Xd_0__inst_product1_31__2__q ;
wire Xd_0__inst_product1_30__2__q ;
wire Xd_0__inst_product1_25__2__q ;
wire Xd_0__inst_product1_24__2__q ;
wire Xd_0__inst_product1_27__2__q ;
wire Xd_0__inst_product1_26__2__q ;
wire Xd_0__inst_product1_21__2__q ;
wire Xd_0__inst_product1_20__2__q ;
wire Xd_0__inst_product1_23__2__q ;
wire Xd_0__inst_product1_22__2__q ;
wire Xd_0__inst_product1_17__2__q ;
wire Xd_0__inst_product1_16__2__q ;
wire Xd_0__inst_product1_19__2__q ;
wire Xd_0__inst_product1_18__2__q ;
wire Xd_0__inst_product1_13__2__q ;
wire Xd_0__inst_product1_12__2__q ;
wire Xd_0__inst_product1_15__2__q ;
wire Xd_0__inst_product1_14__2__q ;
wire Xd_0__inst_product1_9__2__q ;
wire Xd_0__inst_product1_8__2__q ;
wire Xd_0__inst_product1_11__2__q ;
wire Xd_0__inst_product1_10__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_29__3__q ;
wire Xd_0__inst_product1_28__3__q ;
wire Xd_0__inst_product1_31__3__q ;
wire Xd_0__inst_product1_30__3__q ;
wire Xd_0__inst_product1_25__3__q ;
wire Xd_0__inst_product1_24__3__q ;
wire Xd_0__inst_product1_27__3__q ;
wire Xd_0__inst_product1_26__3__q ;
wire Xd_0__inst_product1_21__3__q ;
wire Xd_0__inst_product1_20__3__q ;
wire Xd_0__inst_product1_23__3__q ;
wire Xd_0__inst_product1_22__3__q ;
wire Xd_0__inst_product1_17__3__q ;
wire Xd_0__inst_product1_16__3__q ;
wire Xd_0__inst_product1_19__3__q ;
wire Xd_0__inst_product1_18__3__q ;
wire Xd_0__inst_product1_13__3__q ;
wire Xd_0__inst_product1_12__3__q ;
wire Xd_0__inst_product1_15__3__q ;
wire Xd_0__inst_product1_14__3__q ;
wire Xd_0__inst_product1_9__3__q ;
wire Xd_0__inst_product1_8__3__q ;
wire Xd_0__inst_product1_11__3__q ;
wire Xd_0__inst_product1_10__3__q ;
wire Xd_0__inst_product1_5__3__q ;
wire Xd_0__inst_product1_4__3__q ;
wire Xd_0__inst_product1_7__3__q ;
wire Xd_0__inst_product1_6__3__q ;
wire Xd_0__inst_product1_1__3__q ;
wire Xd_0__inst_product1_0__3__q ;
wire Xd_0__inst_product1_3__3__q ;
wire Xd_0__inst_product1_2__3__q ;
wire Xd_0__inst_product1_29__4__q ;
wire Xd_0__inst_product1_28__4__q ;
wire Xd_0__inst_product1_31__4__q ;
wire Xd_0__inst_product1_30__4__q ;
wire Xd_0__inst_product1_25__4__q ;
wire Xd_0__inst_product1_24__4__q ;
wire Xd_0__inst_product1_27__4__q ;
wire Xd_0__inst_product1_26__4__q ;
wire Xd_0__inst_product1_21__4__q ;
wire Xd_0__inst_product1_20__4__q ;
wire Xd_0__inst_product1_23__4__q ;
wire Xd_0__inst_product1_22__4__q ;
wire Xd_0__inst_product1_17__4__q ;
wire Xd_0__inst_product1_16__4__q ;
wire Xd_0__inst_product1_19__4__q ;
wire Xd_0__inst_product1_18__4__q ;
wire Xd_0__inst_product1_13__4__q ;
wire Xd_0__inst_product1_12__4__q ;
wire Xd_0__inst_product1_15__4__q ;
wire Xd_0__inst_product1_14__4__q ;
wire Xd_0__inst_product1_9__4__q ;
wire Xd_0__inst_product1_8__4__q ;
wire Xd_0__inst_product1_11__4__q ;
wire Xd_0__inst_product1_10__4__q ;
wire Xd_0__inst_product1_5__4__q ;
wire Xd_0__inst_product1_4__4__q ;
wire Xd_0__inst_product1_7__4__q ;
wire Xd_0__inst_product1_6__4__q ;
wire Xd_0__inst_product1_1__4__q ;
wire Xd_0__inst_product1_0__4__q ;
wire Xd_0__inst_product1_3__4__q ;
wire Xd_0__inst_product1_2__4__q ;
wire Xd_0__inst_mult_29_0_q ;
wire Xd_0__inst_mult_29_1_q ;
wire Xd_0__inst_mult_28_0_q ;
wire Xd_0__inst_mult_28_1_q ;
wire Xd_0__inst_mult_31_0_q ;
wire Xd_0__inst_mult_31_1_q ;
wire Xd_0__inst_mult_30_0_q ;
wire Xd_0__inst_mult_30_1_q ;
wire Xd_0__inst_mult_25_0_q ;
wire Xd_0__inst_mult_25_1_q ;
wire Xd_0__inst_mult_24_0_q ;
wire Xd_0__inst_mult_24_1_q ;
wire Xd_0__inst_mult_27_0_q ;
wire Xd_0__inst_mult_27_1_q ;
wire Xd_0__inst_mult_26_0_q ;
wire Xd_0__inst_mult_26_1_q ;
wire Xd_0__inst_mult_21_0_q ;
wire Xd_0__inst_mult_21_1_q ;
wire Xd_0__inst_mult_20_0_q ;
wire Xd_0__inst_mult_20_1_q ;
wire Xd_0__inst_mult_23_0_q ;
wire Xd_0__inst_mult_23_1_q ;
wire Xd_0__inst_mult_22_0_q ;
wire Xd_0__inst_mult_22_1_q ;
wire Xd_0__inst_mult_17_0_q ;
wire Xd_0__inst_mult_17_1_q ;
wire Xd_0__inst_mult_16_0_q ;
wire Xd_0__inst_mult_16_1_q ;
wire Xd_0__inst_mult_19_0_q ;
wire Xd_0__inst_mult_19_1_q ;
wire Xd_0__inst_mult_18_0_q ;
wire Xd_0__inst_mult_18_1_q ;
wire Xd_0__inst_mult_13_0_q ;
wire Xd_0__inst_mult_13_1_q ;
wire Xd_0__inst_mult_12_0_q ;
wire Xd_0__inst_mult_12_1_q ;
wire Xd_0__inst_mult_15_0_q ;
wire Xd_0__inst_mult_15_1_q ;
wire Xd_0__inst_mult_14_0_q ;
wire Xd_0__inst_mult_14_1_q ;
wire Xd_0__inst_mult_9_0_q ;
wire Xd_0__inst_mult_9_1_q ;
wire Xd_0__inst_mult_8_0_q ;
wire Xd_0__inst_mult_8_1_q ;
wire Xd_0__inst_mult_11_0_q ;
wire Xd_0__inst_mult_11_1_q ;
wire Xd_0__inst_mult_10_0_q ;
wire Xd_0__inst_mult_10_1_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_1_0_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_mult_29_2_q ;
wire Xd_0__inst_mult_29_3_q ;
wire Xd_0__inst_mult_28_2_q ;
wire Xd_0__inst_mult_28_3_q ;
wire Xd_0__inst_mult_31_2_q ;
wire Xd_0__inst_mult_31_3_q ;
wire Xd_0__inst_mult_30_2_q ;
wire Xd_0__inst_mult_30_3_q ;
wire Xd_0__inst_mult_25_2_q ;
wire Xd_0__inst_mult_25_3_q ;
wire Xd_0__inst_mult_24_2_q ;
wire Xd_0__inst_mult_24_3_q ;
wire Xd_0__inst_mult_27_2_q ;
wire Xd_0__inst_mult_27_3_q ;
wire Xd_0__inst_mult_26_2_q ;
wire Xd_0__inst_mult_26_3_q ;
wire Xd_0__inst_mult_21_2_q ;
wire Xd_0__inst_mult_21_3_q ;
wire Xd_0__inst_mult_20_2_q ;
wire Xd_0__inst_mult_20_3_q ;
wire Xd_0__inst_mult_23_2_q ;
wire Xd_0__inst_mult_23_3_q ;
wire Xd_0__inst_mult_22_2_q ;
wire Xd_0__inst_mult_22_3_q ;
wire Xd_0__inst_mult_17_2_q ;
wire Xd_0__inst_mult_17_3_q ;
wire Xd_0__inst_mult_16_2_q ;
wire Xd_0__inst_mult_16_3_q ;
wire Xd_0__inst_mult_19_2_q ;
wire Xd_0__inst_mult_19_3_q ;
wire Xd_0__inst_mult_18_2_q ;
wire Xd_0__inst_mult_18_3_q ;
wire Xd_0__inst_mult_13_2_q ;
wire Xd_0__inst_mult_13_3_q ;
wire Xd_0__inst_mult_12_2_q ;
wire Xd_0__inst_mult_12_3_q ;
wire Xd_0__inst_mult_15_2_q ;
wire Xd_0__inst_mult_15_3_q ;
wire Xd_0__inst_mult_14_2_q ;
wire Xd_0__inst_mult_14_3_q ;
wire Xd_0__inst_mult_9_2_q ;
wire Xd_0__inst_mult_9_3_q ;
wire Xd_0__inst_mult_8_2_q ;
wire Xd_0__inst_mult_8_3_q ;
wire Xd_0__inst_mult_11_2_q ;
wire Xd_0__inst_mult_11_3_q ;
wire Xd_0__inst_mult_10_2_q ;
wire Xd_0__inst_mult_10_3_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_29_4_q ;
wire Xd_0__inst_mult_29_5_q ;
wire Xd_0__inst_mult_28_4_q ;
wire Xd_0__inst_mult_28_5_q ;
wire Xd_0__inst_mult_31_4_q ;
wire Xd_0__inst_mult_31_5_q ;
wire Xd_0__inst_mult_30_4_q ;
wire Xd_0__inst_mult_30_5_q ;
wire Xd_0__inst_mult_25_4_q ;
wire Xd_0__inst_mult_25_5_q ;
wire Xd_0__inst_mult_24_4_q ;
wire Xd_0__inst_mult_24_5_q ;
wire Xd_0__inst_mult_27_4_q ;
wire Xd_0__inst_mult_27_5_q ;
wire Xd_0__inst_mult_26_4_q ;
wire Xd_0__inst_mult_26_5_q ;
wire Xd_0__inst_mult_21_4_q ;
wire Xd_0__inst_mult_21_5_q ;
wire Xd_0__inst_mult_20_4_q ;
wire Xd_0__inst_mult_20_5_q ;
wire Xd_0__inst_mult_23_4_q ;
wire Xd_0__inst_mult_23_5_q ;
wire Xd_0__inst_mult_22_4_q ;
wire Xd_0__inst_mult_22_5_q ;
wire Xd_0__inst_mult_17_4_q ;
wire Xd_0__inst_mult_17_5_q ;
wire Xd_0__inst_mult_16_4_q ;
wire Xd_0__inst_mult_16_5_q ;
wire Xd_0__inst_mult_19_4_q ;
wire Xd_0__inst_mult_19_5_q ;
wire Xd_0__inst_mult_18_4_q ;
wire Xd_0__inst_mult_18_5_q ;
wire Xd_0__inst_mult_13_4_q ;
wire Xd_0__inst_mult_13_5_q ;
wire Xd_0__inst_mult_12_4_q ;
wire Xd_0__inst_mult_12_5_q ;
wire Xd_0__inst_mult_15_4_q ;
wire Xd_0__inst_mult_15_5_q ;
wire Xd_0__inst_mult_14_4_q ;
wire Xd_0__inst_mult_14_5_q ;
wire Xd_0__inst_mult_9_4_q ;
wire Xd_0__inst_mult_9_5_q ;
wire Xd_0__inst_mult_8_4_q ;
wire Xd_0__inst_mult_8_5_q ;
wire Xd_0__inst_mult_11_4_q ;
wire Xd_0__inst_mult_11_5_q ;
wire Xd_0__inst_mult_10_4_q ;
wire Xd_0__inst_mult_10_5_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_29_6_q ;
wire Xd_0__inst_mult_29_7_q ;
wire Xd_0__inst_mult_28_6_q ;
wire Xd_0__inst_mult_28_7_q ;
wire Xd_0__inst_mult_31_6_q ;
wire Xd_0__inst_mult_31_7_q ;
wire Xd_0__inst_mult_30_6_q ;
wire Xd_0__inst_mult_30_7_q ;
wire Xd_0__inst_mult_25_6_q ;
wire Xd_0__inst_mult_25_7_q ;
wire Xd_0__inst_mult_24_6_q ;
wire Xd_0__inst_mult_24_7_q ;
wire Xd_0__inst_mult_27_6_q ;
wire Xd_0__inst_mult_27_7_q ;
wire Xd_0__inst_mult_26_6_q ;
wire Xd_0__inst_mult_26_7_q ;
wire Xd_0__inst_mult_21_6_q ;
wire Xd_0__inst_mult_21_7_q ;
wire Xd_0__inst_mult_20_6_q ;
wire Xd_0__inst_mult_20_7_q ;
wire Xd_0__inst_mult_23_6_q ;
wire Xd_0__inst_mult_23_7_q ;
wire Xd_0__inst_mult_22_6_q ;
wire Xd_0__inst_mult_22_7_q ;
wire Xd_0__inst_mult_17_6_q ;
wire Xd_0__inst_mult_17_7_q ;
wire Xd_0__inst_mult_16_6_q ;
wire Xd_0__inst_mult_16_7_q ;
wire Xd_0__inst_mult_19_6_q ;
wire Xd_0__inst_mult_19_7_q ;
wire Xd_0__inst_mult_18_6_q ;
wire Xd_0__inst_mult_18_7_q ;
wire Xd_0__inst_mult_13_6_q ;
wire Xd_0__inst_mult_13_7_q ;
wire Xd_0__inst_mult_12_6_q ;
wire Xd_0__inst_mult_12_7_q ;
wire Xd_0__inst_mult_15_6_q ;
wire Xd_0__inst_mult_15_7_q ;
wire Xd_0__inst_mult_14_6_q ;
wire Xd_0__inst_mult_14_7_q ;
wire Xd_0__inst_mult_9_6_q ;
wire Xd_0__inst_mult_9_7_q ;
wire Xd_0__inst_mult_8_6_q ;
wire Xd_0__inst_mult_8_7_q ;
wire Xd_0__inst_mult_11_6_q ;
wire Xd_0__inst_mult_11_7_q ;
wire Xd_0__inst_mult_10_6_q ;
wire Xd_0__inst_mult_10_7_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_29_8_q ;
wire Xd_0__inst_mult_29_9_q ;
wire Xd_0__inst_mult_28_8_q ;
wire Xd_0__inst_mult_28_9_q ;
wire Xd_0__inst_mult_31_8_q ;
wire Xd_0__inst_mult_31_9_q ;
wire Xd_0__inst_mult_30_8_q ;
wire Xd_0__inst_mult_30_9_q ;
wire Xd_0__inst_mult_25_8_q ;
wire Xd_0__inst_mult_25_9_q ;
wire Xd_0__inst_mult_24_8_q ;
wire Xd_0__inst_mult_24_9_q ;
wire Xd_0__inst_mult_27_8_q ;
wire Xd_0__inst_mult_27_9_q ;
wire Xd_0__inst_mult_26_8_q ;
wire Xd_0__inst_mult_26_9_q ;
wire Xd_0__inst_mult_21_8_q ;
wire Xd_0__inst_mult_21_9_q ;
wire Xd_0__inst_mult_20_8_q ;
wire Xd_0__inst_mult_20_9_q ;
wire Xd_0__inst_mult_23_8_q ;
wire Xd_0__inst_mult_23_9_q ;
wire Xd_0__inst_mult_22_8_q ;
wire Xd_0__inst_mult_22_9_q ;
wire Xd_0__inst_mult_17_8_q ;
wire Xd_0__inst_mult_17_9_q ;
wire Xd_0__inst_mult_16_8_q ;
wire Xd_0__inst_mult_16_9_q ;
wire Xd_0__inst_mult_19_8_q ;
wire Xd_0__inst_mult_19_9_q ;
wire Xd_0__inst_mult_18_8_q ;
wire Xd_0__inst_mult_18_9_q ;
wire Xd_0__inst_mult_13_8_q ;
wire Xd_0__inst_mult_13_9_q ;
wire Xd_0__inst_mult_12_8_q ;
wire Xd_0__inst_mult_12_9_q ;
wire Xd_0__inst_mult_15_8_q ;
wire Xd_0__inst_mult_15_9_q ;
wire Xd_0__inst_mult_14_8_q ;
wire Xd_0__inst_mult_14_9_q ;
wire Xd_0__inst_mult_9_8_q ;
wire Xd_0__inst_mult_9_9_q ;
wire Xd_0__inst_mult_8_8_q ;
wire Xd_0__inst_mult_8_9_q ;
wire Xd_0__inst_mult_11_8_q ;
wire Xd_0__inst_mult_11_9_q ;
wire Xd_0__inst_mult_10_8_q ;
wire Xd_0__inst_mult_10_9_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_29_10_q ;
wire Xd_0__inst_mult_29_11_q ;
wire Xd_0__inst_mult_28_10_q ;
wire Xd_0__inst_mult_28_11_q ;
wire Xd_0__inst_mult_31_10_q ;
wire Xd_0__inst_mult_31_11_q ;
wire Xd_0__inst_mult_30_10_q ;
wire Xd_0__inst_mult_30_11_q ;
wire Xd_0__inst_mult_25_10_q ;
wire Xd_0__inst_mult_25_11_q ;
wire Xd_0__inst_mult_24_10_q ;
wire Xd_0__inst_mult_24_11_q ;
wire Xd_0__inst_mult_27_10_q ;
wire Xd_0__inst_mult_27_11_q ;
wire Xd_0__inst_mult_26_10_q ;
wire Xd_0__inst_mult_26_11_q ;
wire Xd_0__inst_mult_21_10_q ;
wire Xd_0__inst_mult_21_11_q ;
wire Xd_0__inst_mult_20_10_q ;
wire Xd_0__inst_mult_20_11_q ;
wire Xd_0__inst_mult_23_10_q ;
wire Xd_0__inst_mult_23_11_q ;
wire Xd_0__inst_mult_22_10_q ;
wire Xd_0__inst_mult_22_11_q ;
wire Xd_0__inst_mult_17_10_q ;
wire Xd_0__inst_mult_17_11_q ;
wire Xd_0__inst_mult_16_10_q ;
wire Xd_0__inst_mult_16_11_q ;
wire Xd_0__inst_mult_19_10_q ;
wire Xd_0__inst_mult_19_11_q ;
wire Xd_0__inst_mult_18_10_q ;
wire Xd_0__inst_mult_18_11_q ;
wire Xd_0__inst_mult_13_10_q ;
wire Xd_0__inst_mult_13_11_q ;
wire Xd_0__inst_mult_12_10_q ;
wire Xd_0__inst_mult_12_11_q ;
wire Xd_0__inst_mult_15_10_q ;
wire Xd_0__inst_mult_15_11_q ;
wire Xd_0__inst_mult_14_10_q ;
wire Xd_0__inst_mult_14_11_q ;
wire Xd_0__inst_mult_9_10_q ;
wire Xd_0__inst_mult_9_11_q ;
wire Xd_0__inst_mult_8_10_q ;
wire Xd_0__inst_mult_8_11_q ;
wire Xd_0__inst_mult_11_10_q ;
wire Xd_0__inst_mult_11_11_q ;
wire Xd_0__inst_mult_10_10_q ;
wire Xd_0__inst_mult_10_11_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_29_12_q ;
wire Xd_0__inst_mult_29_13_q ;
wire Xd_0__inst_mult_28_12_q ;
wire Xd_0__inst_mult_28_13_q ;
wire Xd_0__inst_mult_31_12_q ;
wire Xd_0__inst_mult_31_13_q ;
wire Xd_0__inst_mult_30_12_q ;
wire Xd_0__inst_mult_30_13_q ;
wire Xd_0__inst_mult_25_12_q ;
wire Xd_0__inst_mult_25_13_q ;
wire Xd_0__inst_mult_24_12_q ;
wire Xd_0__inst_mult_24_13_q ;
wire Xd_0__inst_mult_27_12_q ;
wire Xd_0__inst_mult_27_13_q ;
wire Xd_0__inst_mult_26_12_q ;
wire Xd_0__inst_mult_26_13_q ;
wire Xd_0__inst_mult_21_12_q ;
wire Xd_0__inst_mult_21_13_q ;
wire Xd_0__inst_mult_20_12_q ;
wire Xd_0__inst_mult_20_13_q ;
wire Xd_0__inst_mult_23_12_q ;
wire Xd_0__inst_mult_23_13_q ;
wire Xd_0__inst_mult_22_12_q ;
wire Xd_0__inst_mult_22_13_q ;
wire Xd_0__inst_mult_17_12_q ;
wire Xd_0__inst_mult_17_13_q ;
wire Xd_0__inst_mult_16_12_q ;
wire Xd_0__inst_mult_16_13_q ;
wire Xd_0__inst_mult_19_12_q ;
wire Xd_0__inst_mult_19_13_q ;
wire Xd_0__inst_mult_18_12_q ;
wire Xd_0__inst_mult_18_13_q ;
wire Xd_0__inst_mult_13_12_q ;
wire Xd_0__inst_mult_13_13_q ;
wire Xd_0__inst_mult_12_12_q ;
wire Xd_0__inst_mult_12_13_q ;
wire Xd_0__inst_mult_15_12_q ;
wire Xd_0__inst_mult_15_13_q ;
wire Xd_0__inst_mult_14_12_q ;
wire Xd_0__inst_mult_14_13_q ;
wire Xd_0__inst_mult_9_12_q ;
wire Xd_0__inst_mult_9_13_q ;
wire Xd_0__inst_mult_8_12_q ;
wire Xd_0__inst_mult_8_13_q ;
wire Xd_0__inst_mult_11_12_q ;
wire Xd_0__inst_mult_11_13_q ;
wire Xd_0__inst_mult_10_12_q ;
wire Xd_0__inst_mult_10_13_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_29_14_q ;
wire Xd_0__inst_mult_29_15_q ;
wire Xd_0__inst_mult_28_14_q ;
wire Xd_0__inst_mult_28_15_q ;
wire Xd_0__inst_mult_31_14_q ;
wire Xd_0__inst_mult_31_15_q ;
wire Xd_0__inst_mult_30_14_q ;
wire Xd_0__inst_mult_30_15_q ;
wire Xd_0__inst_mult_25_14_q ;
wire Xd_0__inst_mult_25_15_q ;
wire Xd_0__inst_mult_24_14_q ;
wire Xd_0__inst_mult_24_15_q ;
wire Xd_0__inst_mult_27_14_q ;
wire Xd_0__inst_mult_27_15_q ;
wire Xd_0__inst_mult_26_14_q ;
wire Xd_0__inst_mult_26_15_q ;
wire Xd_0__inst_mult_21_14_q ;
wire Xd_0__inst_mult_21_15_q ;
wire Xd_0__inst_mult_20_14_q ;
wire Xd_0__inst_mult_20_15_q ;
wire Xd_0__inst_mult_23_14_q ;
wire Xd_0__inst_mult_23_15_q ;
wire Xd_0__inst_mult_22_14_q ;
wire Xd_0__inst_mult_22_15_q ;
wire Xd_0__inst_mult_17_14_q ;
wire Xd_0__inst_mult_17_15_q ;
wire Xd_0__inst_mult_16_14_q ;
wire Xd_0__inst_mult_16_15_q ;
wire Xd_0__inst_mult_19_14_q ;
wire Xd_0__inst_mult_19_15_q ;
wire Xd_0__inst_mult_18_14_q ;
wire Xd_0__inst_mult_18_15_q ;
wire Xd_0__inst_mult_13_14_q ;
wire Xd_0__inst_mult_13_15_q ;
wire Xd_0__inst_mult_12_14_q ;
wire Xd_0__inst_mult_12_15_q ;
wire Xd_0__inst_mult_15_14_q ;
wire Xd_0__inst_mult_15_15_q ;
wire Xd_0__inst_mult_14_14_q ;
wire Xd_0__inst_mult_14_15_q ;
wire Xd_0__inst_mult_9_14_q ;
wire Xd_0__inst_mult_9_15_q ;
wire Xd_0__inst_mult_8_14_q ;
wire Xd_0__inst_mult_8_15_q ;
wire Xd_0__inst_mult_11_14_q ;
wire Xd_0__inst_mult_11_15_q ;
wire Xd_0__inst_mult_10_14_q ;
wire Xd_0__inst_mult_10_15_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_29_16_q ;
wire Xd_0__inst_mult_29_17_q ;
wire Xd_0__inst_mult_28_16_q ;
wire Xd_0__inst_mult_28_17_q ;
wire Xd_0__inst_mult_31_16_q ;
wire Xd_0__inst_mult_31_17_q ;
wire Xd_0__inst_mult_30_16_q ;
wire Xd_0__inst_mult_30_17_q ;
wire Xd_0__inst_mult_25_16_q ;
wire Xd_0__inst_mult_25_17_q ;
wire Xd_0__inst_mult_24_16_q ;
wire Xd_0__inst_mult_24_17_q ;
wire Xd_0__inst_mult_27_16_q ;
wire Xd_0__inst_mult_27_17_q ;
wire Xd_0__inst_mult_26_16_q ;
wire Xd_0__inst_mult_26_17_q ;
wire Xd_0__inst_mult_21_16_q ;
wire Xd_0__inst_mult_21_17_q ;
wire Xd_0__inst_mult_20_16_q ;
wire Xd_0__inst_mult_20_17_q ;
wire Xd_0__inst_mult_23_16_q ;
wire Xd_0__inst_mult_23_17_q ;
wire Xd_0__inst_mult_22_16_q ;
wire Xd_0__inst_mult_22_17_q ;
wire Xd_0__inst_mult_17_16_q ;
wire Xd_0__inst_mult_17_17_q ;
wire Xd_0__inst_mult_16_16_q ;
wire Xd_0__inst_mult_16_17_q ;
wire Xd_0__inst_mult_19_16_q ;
wire Xd_0__inst_mult_19_17_q ;
wire Xd_0__inst_mult_18_16_q ;
wire Xd_0__inst_mult_18_17_q ;
wire Xd_0__inst_mult_13_16_q ;
wire Xd_0__inst_mult_13_17_q ;
wire Xd_0__inst_mult_12_16_q ;
wire Xd_0__inst_mult_12_17_q ;
wire Xd_0__inst_mult_15_16_q ;
wire Xd_0__inst_mult_15_17_q ;
wire Xd_0__inst_mult_14_16_q ;
wire Xd_0__inst_mult_14_17_q ;
wire Xd_0__inst_mult_9_16_q ;
wire Xd_0__inst_mult_9_17_q ;
wire Xd_0__inst_mult_8_16_q ;
wire Xd_0__inst_mult_8_17_q ;
wire Xd_0__inst_mult_11_16_q ;
wire Xd_0__inst_mult_11_17_q ;
wire Xd_0__inst_mult_10_16_q ;
wire Xd_0__inst_mult_10_17_q ;
wire Xd_0__inst_mult_5_16_q ;
wire Xd_0__inst_mult_5_17_q ;
wire Xd_0__inst_mult_4_16_q ;
wire Xd_0__inst_mult_4_17_q ;
wire Xd_0__inst_mult_7_16_q ;
wire Xd_0__inst_mult_7_17_q ;
wire Xd_0__inst_mult_6_16_q ;
wire Xd_0__inst_mult_6_17_q ;
wire Xd_0__inst_mult_1_16_q ;
wire Xd_0__inst_mult_1_17_q ;
wire Xd_0__inst_mult_0_16_q ;
wire Xd_0__inst_mult_0_17_q ;
wire Xd_0__inst_mult_3_16_q ;
wire Xd_0__inst_mult_3_17_q ;
wire Xd_0__inst_mult_2_16_q ;
wire Xd_0__inst_mult_2_17_q ;
wire Xd_0__inst_mult_29_18_q ;
wire Xd_0__inst_mult_29_19_q ;
wire Xd_0__inst_mult_28_18_q ;
wire Xd_0__inst_mult_28_19_q ;
wire Xd_0__inst_mult_31_18_q ;
wire Xd_0__inst_mult_31_19_q ;
wire Xd_0__inst_mult_30_18_q ;
wire Xd_0__inst_mult_30_19_q ;
wire Xd_0__inst_mult_25_18_q ;
wire Xd_0__inst_mult_25_19_q ;
wire Xd_0__inst_mult_24_18_q ;
wire Xd_0__inst_mult_24_19_q ;
wire Xd_0__inst_mult_27_18_q ;
wire Xd_0__inst_mult_27_19_q ;
wire Xd_0__inst_mult_26_18_q ;
wire Xd_0__inst_mult_26_19_q ;
wire Xd_0__inst_mult_21_18_q ;
wire Xd_0__inst_mult_21_19_q ;
wire Xd_0__inst_mult_20_18_q ;
wire Xd_0__inst_mult_20_19_q ;
wire Xd_0__inst_mult_23_18_q ;
wire Xd_0__inst_mult_23_19_q ;
wire Xd_0__inst_mult_22_18_q ;
wire Xd_0__inst_mult_22_19_q ;
wire Xd_0__inst_mult_17_18_q ;
wire Xd_0__inst_mult_17_19_q ;
wire Xd_0__inst_mult_16_18_q ;
wire Xd_0__inst_mult_16_19_q ;
wire Xd_0__inst_mult_19_18_q ;
wire Xd_0__inst_mult_19_19_q ;
wire Xd_0__inst_mult_18_18_q ;
wire Xd_0__inst_mult_18_19_q ;
wire Xd_0__inst_mult_13_18_q ;
wire Xd_0__inst_mult_13_19_q ;
wire Xd_0__inst_mult_12_18_q ;
wire Xd_0__inst_mult_12_19_q ;
wire Xd_0__inst_mult_15_18_q ;
wire Xd_0__inst_mult_15_19_q ;
wire Xd_0__inst_mult_14_18_q ;
wire Xd_0__inst_mult_14_19_q ;
wire Xd_0__inst_mult_9_18_q ;
wire Xd_0__inst_mult_9_19_q ;
wire Xd_0__inst_mult_8_18_q ;
wire Xd_0__inst_mult_8_19_q ;
wire Xd_0__inst_mult_11_18_q ;
wire Xd_0__inst_mult_11_19_q ;
wire Xd_0__inst_mult_10_18_q ;
wire Xd_0__inst_mult_10_19_q ;
wire Xd_0__inst_mult_5_18_q ;
wire Xd_0__inst_mult_5_19_q ;
wire Xd_0__inst_mult_4_18_q ;
wire Xd_0__inst_mult_4_19_q ;
wire Xd_0__inst_mult_7_18_q ;
wire Xd_0__inst_mult_7_19_q ;
wire Xd_0__inst_mult_6_18_q ;
wire Xd_0__inst_mult_6_19_q ;
wire Xd_0__inst_mult_1_18_q ;
wire Xd_0__inst_mult_1_19_q ;
wire Xd_0__inst_mult_0_18_q ;
wire Xd_0__inst_mult_0_19_q ;
wire Xd_0__inst_mult_3_18_q ;
wire Xd_0__inst_mult_3_19_q ;
wire Xd_0__inst_mult_2_18_q ;
wire Xd_0__inst_mult_2_19_q ;
wire Xd_0__inst_mult_29_20_q ;
wire Xd_0__inst_mult_29_21_q ;
wire Xd_0__inst_mult_29_22_q ;
wire Xd_0__inst_mult_29_23_q ;
wire Xd_0__inst_mult_28_20_q ;
wire Xd_0__inst_mult_28_21_q ;
wire Xd_0__inst_mult_28_22_q ;
wire Xd_0__inst_mult_28_23_q ;
wire Xd_0__inst_mult_31_20_q ;
wire Xd_0__inst_mult_31_21_q ;
wire Xd_0__inst_mult_31_22_q ;
wire Xd_0__inst_mult_31_23_q ;
wire Xd_0__inst_mult_30_20_q ;
wire Xd_0__inst_mult_30_21_q ;
wire Xd_0__inst_mult_30_22_q ;
wire Xd_0__inst_mult_30_23_q ;
wire Xd_0__inst_mult_25_20_q ;
wire Xd_0__inst_mult_25_21_q ;
wire Xd_0__inst_mult_25_22_q ;
wire Xd_0__inst_mult_25_23_q ;
wire Xd_0__inst_mult_24_20_q ;
wire Xd_0__inst_mult_24_21_q ;
wire Xd_0__inst_mult_24_22_q ;
wire Xd_0__inst_mult_24_23_q ;
wire Xd_0__inst_mult_27_20_q ;
wire Xd_0__inst_mult_27_21_q ;
wire Xd_0__inst_mult_27_22_q ;
wire Xd_0__inst_mult_27_23_q ;
wire Xd_0__inst_mult_26_20_q ;
wire Xd_0__inst_mult_26_21_q ;
wire Xd_0__inst_mult_26_22_q ;
wire Xd_0__inst_mult_26_23_q ;
wire Xd_0__inst_mult_21_20_q ;
wire Xd_0__inst_mult_21_21_q ;
wire Xd_0__inst_mult_21_22_q ;
wire Xd_0__inst_mult_21_23_q ;
wire Xd_0__inst_mult_20_20_q ;
wire Xd_0__inst_mult_20_21_q ;
wire Xd_0__inst_mult_20_22_q ;
wire Xd_0__inst_mult_20_23_q ;
wire Xd_0__inst_mult_23_20_q ;
wire Xd_0__inst_mult_23_21_q ;
wire Xd_0__inst_mult_23_22_q ;
wire Xd_0__inst_mult_23_23_q ;
wire Xd_0__inst_mult_22_20_q ;
wire Xd_0__inst_mult_22_21_q ;
wire Xd_0__inst_mult_22_22_q ;
wire Xd_0__inst_mult_22_23_q ;
wire Xd_0__inst_mult_17_20_q ;
wire Xd_0__inst_mult_17_21_q ;
wire Xd_0__inst_mult_17_22_q ;
wire Xd_0__inst_mult_17_23_q ;
wire Xd_0__inst_mult_16_20_q ;
wire Xd_0__inst_mult_16_21_q ;
wire Xd_0__inst_mult_16_22_q ;
wire Xd_0__inst_mult_16_23_q ;
wire Xd_0__inst_mult_19_20_q ;
wire Xd_0__inst_mult_19_21_q ;
wire Xd_0__inst_mult_19_22_q ;
wire Xd_0__inst_mult_19_23_q ;
wire Xd_0__inst_mult_18_20_q ;
wire Xd_0__inst_mult_18_21_q ;
wire Xd_0__inst_mult_18_22_q ;
wire Xd_0__inst_mult_18_23_q ;
wire Xd_0__inst_mult_13_20_q ;
wire Xd_0__inst_mult_13_21_q ;
wire Xd_0__inst_mult_13_22_q ;
wire Xd_0__inst_mult_13_23_q ;
wire Xd_0__inst_mult_12_20_q ;
wire Xd_0__inst_mult_12_21_q ;
wire Xd_0__inst_mult_12_22_q ;
wire Xd_0__inst_mult_12_23_q ;
wire Xd_0__inst_mult_15_20_q ;
wire Xd_0__inst_mult_15_21_q ;
wire Xd_0__inst_mult_15_22_q ;
wire Xd_0__inst_mult_15_23_q ;
wire Xd_0__inst_mult_14_20_q ;
wire Xd_0__inst_mult_14_21_q ;
wire Xd_0__inst_mult_14_22_q ;
wire Xd_0__inst_mult_14_23_q ;
wire Xd_0__inst_mult_9_20_q ;
wire Xd_0__inst_mult_9_21_q ;
wire Xd_0__inst_mult_9_22_q ;
wire Xd_0__inst_mult_9_23_q ;
wire Xd_0__inst_mult_8_20_q ;
wire Xd_0__inst_mult_8_21_q ;
wire Xd_0__inst_mult_8_22_q ;
wire Xd_0__inst_mult_8_23_q ;
wire Xd_0__inst_mult_11_20_q ;
wire Xd_0__inst_mult_11_21_q ;
wire Xd_0__inst_mult_11_22_q ;
wire Xd_0__inst_mult_11_23_q ;
wire Xd_0__inst_mult_10_20_q ;
wire Xd_0__inst_mult_10_21_q ;
wire Xd_0__inst_mult_10_22_q ;
wire Xd_0__inst_mult_10_23_q ;
wire Xd_0__inst_mult_5_20_q ;
wire Xd_0__inst_mult_5_21_q ;
wire Xd_0__inst_mult_5_22_q ;
wire Xd_0__inst_mult_5_23_q ;
wire Xd_0__inst_mult_4_20_q ;
wire Xd_0__inst_mult_4_21_q ;
wire Xd_0__inst_mult_4_22_q ;
wire Xd_0__inst_mult_4_23_q ;
wire Xd_0__inst_mult_7_20_q ;
wire Xd_0__inst_mult_7_21_q ;
wire Xd_0__inst_mult_7_22_q ;
wire Xd_0__inst_mult_7_23_q ;
wire Xd_0__inst_mult_6_20_q ;
wire Xd_0__inst_mult_6_21_q ;
wire Xd_0__inst_mult_6_22_q ;
wire Xd_0__inst_mult_6_23_q ;
wire Xd_0__inst_mult_1_20_q ;
wire Xd_0__inst_mult_1_21_q ;
wire Xd_0__inst_mult_1_22_q ;
wire Xd_0__inst_mult_1_23_q ;
wire Xd_0__inst_mult_0_20_q ;
wire Xd_0__inst_mult_0_21_q ;
wire Xd_0__inst_mult_0_22_q ;
wire Xd_0__inst_mult_0_23_q ;
wire Xd_0__inst_mult_3_20_q ;
wire Xd_0__inst_mult_3_21_q ;
wire Xd_0__inst_mult_3_22_q ;
wire Xd_0__inst_mult_3_23_q ;
wire Xd_0__inst_mult_2_20_q ;
wire Xd_0__inst_mult_2_21_q ;
wire Xd_0__inst_mult_2_22_q ;
wire Xd_0__inst_mult_2_23_q ;
wire Xd_0__inst_mult_29_24_q ;
wire Xd_0__inst_mult_29_25_q ;
wire Xd_0__inst_mult_28_24_q ;
wire Xd_0__inst_mult_28_25_q ;
wire Xd_0__inst_mult_31_24_q ;
wire Xd_0__inst_mult_31_25_q ;
wire Xd_0__inst_mult_30_24_q ;
wire Xd_0__inst_mult_30_25_q ;
wire Xd_0__inst_mult_25_24_q ;
wire Xd_0__inst_mult_25_25_q ;
wire Xd_0__inst_mult_24_24_q ;
wire Xd_0__inst_mult_24_25_q ;
wire Xd_0__inst_mult_27_24_q ;
wire Xd_0__inst_mult_27_25_q ;
wire Xd_0__inst_mult_26_24_q ;
wire Xd_0__inst_mult_26_25_q ;
wire Xd_0__inst_mult_21_24_q ;
wire Xd_0__inst_mult_21_25_q ;
wire Xd_0__inst_mult_20_24_q ;
wire Xd_0__inst_mult_20_25_q ;
wire Xd_0__inst_mult_23_24_q ;
wire Xd_0__inst_mult_23_25_q ;
wire Xd_0__inst_mult_22_24_q ;
wire Xd_0__inst_mult_22_25_q ;
wire Xd_0__inst_mult_17_24_q ;
wire Xd_0__inst_mult_17_25_q ;
wire Xd_0__inst_mult_16_24_q ;
wire Xd_0__inst_mult_16_25_q ;
wire Xd_0__inst_mult_19_24_q ;
wire Xd_0__inst_mult_19_25_q ;
wire Xd_0__inst_mult_18_24_q ;
wire Xd_0__inst_mult_18_25_q ;
wire Xd_0__inst_mult_13_24_q ;
wire Xd_0__inst_mult_13_25_q ;
wire Xd_0__inst_mult_12_24_q ;
wire Xd_0__inst_mult_12_25_q ;
wire Xd_0__inst_mult_15_24_q ;
wire Xd_0__inst_mult_15_25_q ;
wire Xd_0__inst_mult_14_24_q ;
wire Xd_0__inst_mult_14_25_q ;
wire Xd_0__inst_mult_9_24_q ;
wire Xd_0__inst_mult_9_25_q ;
wire Xd_0__inst_mult_8_24_q ;
wire Xd_0__inst_mult_8_25_q ;
wire Xd_0__inst_mult_11_24_q ;
wire Xd_0__inst_mult_11_25_q ;
wire Xd_0__inst_mult_10_24_q ;
wire Xd_0__inst_mult_10_25_q ;
wire Xd_0__inst_mult_5_24_q ;
wire Xd_0__inst_mult_5_25_q ;
wire Xd_0__inst_mult_4_24_q ;
wire Xd_0__inst_mult_4_25_q ;
wire Xd_0__inst_mult_7_24_q ;
wire Xd_0__inst_mult_7_25_q ;
wire Xd_0__inst_mult_6_24_q ;
wire Xd_0__inst_mult_6_25_q ;
wire Xd_0__inst_mult_1_24_q ;
wire Xd_0__inst_mult_1_25_q ;
wire Xd_0__inst_mult_0_24_q ;
wire Xd_0__inst_mult_0_25_q ;
wire Xd_0__inst_mult_3_24_q ;
wire Xd_0__inst_mult_3_25_q ;
wire Xd_0__inst_mult_2_24_q ;
wire Xd_0__inst_mult_2_25_q ;
wire Xd_0__inst_mult_29_26_q ;
wire Xd_0__inst_mult_29_27_q ;
wire Xd_0__inst_mult_28_26_q ;
wire Xd_0__inst_mult_28_27_q ;
wire Xd_0__inst_mult_31_26_q ;
wire Xd_0__inst_mult_31_27_q ;
wire Xd_0__inst_mult_30_26_q ;
wire Xd_0__inst_mult_30_27_q ;
wire Xd_0__inst_mult_25_26_q ;
wire Xd_0__inst_mult_25_27_q ;
wire Xd_0__inst_mult_24_26_q ;
wire Xd_0__inst_mult_24_27_q ;
wire Xd_0__inst_mult_27_26_q ;
wire Xd_0__inst_mult_27_27_q ;
wire Xd_0__inst_mult_26_26_q ;
wire Xd_0__inst_mult_26_27_q ;
wire Xd_0__inst_mult_21_26_q ;
wire Xd_0__inst_mult_21_27_q ;
wire Xd_0__inst_mult_20_26_q ;
wire Xd_0__inst_mult_20_27_q ;
wire Xd_0__inst_mult_23_26_q ;
wire Xd_0__inst_mult_23_27_q ;
wire Xd_0__inst_mult_22_26_q ;
wire Xd_0__inst_mult_22_27_q ;
wire Xd_0__inst_mult_17_26_q ;
wire Xd_0__inst_mult_17_27_q ;
wire Xd_0__inst_mult_16_26_q ;
wire Xd_0__inst_mult_16_27_q ;
wire Xd_0__inst_mult_19_26_q ;
wire Xd_0__inst_mult_19_27_q ;
wire Xd_0__inst_mult_18_26_q ;
wire Xd_0__inst_mult_18_27_q ;
wire Xd_0__inst_mult_13_26_q ;
wire Xd_0__inst_mult_13_27_q ;
wire Xd_0__inst_mult_12_26_q ;
wire Xd_0__inst_mult_12_27_q ;
wire Xd_0__inst_mult_15_26_q ;
wire Xd_0__inst_mult_15_27_q ;
wire Xd_0__inst_mult_14_26_q ;
wire Xd_0__inst_mult_14_27_q ;
wire Xd_0__inst_mult_9_26_q ;
wire Xd_0__inst_mult_9_27_q ;
wire Xd_0__inst_mult_8_26_q ;
wire Xd_0__inst_mult_8_27_q ;
wire Xd_0__inst_mult_11_26_q ;
wire Xd_0__inst_mult_11_27_q ;
wire Xd_0__inst_mult_10_26_q ;
wire Xd_0__inst_mult_10_27_q ;
wire Xd_0__inst_mult_5_26_q ;
wire Xd_0__inst_mult_5_27_q ;
wire Xd_0__inst_mult_4_26_q ;
wire Xd_0__inst_mult_4_27_q ;
wire Xd_0__inst_mult_7_26_q ;
wire Xd_0__inst_mult_7_27_q ;
wire Xd_0__inst_mult_6_26_q ;
wire Xd_0__inst_mult_6_27_q ;
wire Xd_0__inst_mult_1_26_q ;
wire Xd_0__inst_mult_1_27_q ;
wire Xd_0__inst_mult_0_26_q ;
wire Xd_0__inst_mult_0_27_q ;
wire Xd_0__inst_mult_3_26_q ;
wire Xd_0__inst_mult_3_27_q ;
wire Xd_0__inst_mult_2_26_q ;
wire Xd_0__inst_mult_2_27_q ;
wire Xd_0__inst_mult_29_28_q ;
wire Xd_0__inst_mult_29_29_q ;
wire Xd_0__inst_mult_28_28_q ;
wire Xd_0__inst_mult_28_29_q ;
wire Xd_0__inst_mult_31_28_q ;
wire Xd_0__inst_mult_31_29_q ;
wire Xd_0__inst_mult_30_28_q ;
wire Xd_0__inst_mult_30_29_q ;
wire Xd_0__inst_mult_25_28_q ;
wire Xd_0__inst_mult_25_29_q ;
wire Xd_0__inst_mult_24_28_q ;
wire Xd_0__inst_mult_24_29_q ;
wire Xd_0__inst_mult_27_28_q ;
wire Xd_0__inst_mult_27_29_q ;
wire Xd_0__inst_mult_26_28_q ;
wire Xd_0__inst_mult_26_29_q ;
wire Xd_0__inst_mult_21_28_q ;
wire Xd_0__inst_mult_21_29_q ;
wire Xd_0__inst_mult_20_28_q ;
wire Xd_0__inst_mult_20_29_q ;
wire Xd_0__inst_mult_23_28_q ;
wire Xd_0__inst_mult_23_29_q ;
wire Xd_0__inst_mult_22_28_q ;
wire Xd_0__inst_mult_22_29_q ;
wire Xd_0__inst_mult_17_28_q ;
wire Xd_0__inst_mult_17_29_q ;
wire Xd_0__inst_mult_16_28_q ;
wire Xd_0__inst_mult_16_29_q ;
wire Xd_0__inst_mult_19_28_q ;
wire Xd_0__inst_mult_19_29_q ;
wire Xd_0__inst_mult_18_28_q ;
wire Xd_0__inst_mult_18_29_q ;
wire Xd_0__inst_mult_13_28_q ;
wire Xd_0__inst_mult_13_29_q ;
wire Xd_0__inst_mult_12_28_q ;
wire Xd_0__inst_mult_12_29_q ;
wire Xd_0__inst_mult_15_28_q ;
wire Xd_0__inst_mult_15_29_q ;
wire Xd_0__inst_mult_14_28_q ;
wire Xd_0__inst_mult_14_29_q ;
wire Xd_0__inst_mult_9_28_q ;
wire Xd_0__inst_mult_9_29_q ;
wire Xd_0__inst_mult_8_28_q ;
wire Xd_0__inst_mult_8_29_q ;
wire Xd_0__inst_mult_11_28_q ;
wire Xd_0__inst_mult_11_29_q ;
wire Xd_0__inst_mult_10_28_q ;
wire Xd_0__inst_mult_10_29_q ;
wire Xd_0__inst_mult_5_28_q ;
wire Xd_0__inst_mult_5_29_q ;
wire Xd_0__inst_mult_4_28_q ;
wire Xd_0__inst_mult_4_29_q ;
wire Xd_0__inst_mult_7_28_q ;
wire Xd_0__inst_mult_7_29_q ;
wire Xd_0__inst_mult_6_28_q ;
wire Xd_0__inst_mult_6_29_q ;
wire Xd_0__inst_mult_1_28_q ;
wire Xd_0__inst_mult_1_29_q ;
wire Xd_0__inst_mult_0_28_q ;
wire Xd_0__inst_mult_0_29_q ;
wire Xd_0__inst_mult_3_28_q ;
wire Xd_0__inst_mult_3_29_q ;
wire Xd_0__inst_mult_2_28_q ;
wire Xd_0__inst_mult_2_29_q ;
wire Xd_0__inst_mult_29_30_q ;
wire Xd_0__inst_mult_29_31_q ;
wire Xd_0__inst_mult_28_30_q ;
wire Xd_0__inst_mult_28_31_q ;
wire Xd_0__inst_mult_31_30_q ;
wire Xd_0__inst_mult_31_31_q ;
wire Xd_0__inst_mult_30_30_q ;
wire Xd_0__inst_mult_30_31_q ;
wire Xd_0__inst_mult_25_30_q ;
wire Xd_0__inst_mult_25_31_q ;
wire Xd_0__inst_mult_24_30_q ;
wire Xd_0__inst_mult_24_31_q ;
wire Xd_0__inst_mult_27_30_q ;
wire Xd_0__inst_mult_27_31_q ;
wire Xd_0__inst_mult_26_30_q ;
wire Xd_0__inst_mult_26_31_q ;
wire Xd_0__inst_mult_21_30_q ;
wire Xd_0__inst_mult_21_31_q ;
wire Xd_0__inst_mult_20_30_q ;
wire Xd_0__inst_mult_20_31_q ;
wire Xd_0__inst_mult_23_30_q ;
wire Xd_0__inst_mult_23_31_q ;
wire Xd_0__inst_mult_22_30_q ;
wire Xd_0__inst_mult_22_31_q ;
wire Xd_0__inst_mult_17_30_q ;
wire Xd_0__inst_mult_17_31_q ;
wire Xd_0__inst_mult_16_30_q ;
wire Xd_0__inst_mult_16_31_q ;
wire Xd_0__inst_mult_19_30_q ;
wire Xd_0__inst_mult_19_31_q ;
wire Xd_0__inst_mult_18_30_q ;
wire Xd_0__inst_mult_18_31_q ;
wire Xd_0__inst_mult_13_30_q ;
wire Xd_0__inst_mult_13_31_q ;
wire Xd_0__inst_mult_12_30_q ;
wire Xd_0__inst_mult_12_31_q ;
wire Xd_0__inst_mult_15_30_q ;
wire Xd_0__inst_mult_15_31_q ;
wire Xd_0__inst_mult_14_30_q ;
wire Xd_0__inst_mult_14_31_q ;
wire Xd_0__inst_mult_9_30_q ;
wire Xd_0__inst_mult_9_31_q ;
wire Xd_0__inst_mult_8_30_q ;
wire Xd_0__inst_mult_8_31_q ;
wire Xd_0__inst_mult_11_30_q ;
wire Xd_0__inst_mult_11_31_q ;
wire Xd_0__inst_mult_10_30_q ;
wire Xd_0__inst_mult_10_31_q ;
wire Xd_0__inst_mult_5_30_q ;
wire Xd_0__inst_mult_5_31_q ;
wire Xd_0__inst_mult_4_30_q ;
wire Xd_0__inst_mult_4_31_q ;
wire Xd_0__inst_mult_7_30_q ;
wire Xd_0__inst_mult_7_31_q ;
wire Xd_0__inst_mult_6_30_q ;
wire Xd_0__inst_mult_6_31_q ;
wire Xd_0__inst_mult_1_30_q ;
wire Xd_0__inst_mult_1_31_q ;
wire Xd_0__inst_mult_0_30_q ;
wire Xd_0__inst_mult_0_31_q ;
wire Xd_0__inst_mult_3_30_q ;
wire Xd_0__inst_mult_3_31_q ;
wire Xd_0__inst_mult_2_30_q ;
wire Xd_0__inst_mult_2_31_q ;
wire Xd_0__inst_mult_29_32_q ;
wire Xd_0__inst_mult_29_33_q ;
wire Xd_0__inst_mult_28_32_q ;
wire Xd_0__inst_mult_28_33_q ;
wire Xd_0__inst_mult_31_32_q ;
wire Xd_0__inst_mult_31_33_q ;
wire Xd_0__inst_mult_30_32_q ;
wire Xd_0__inst_mult_30_33_q ;
wire Xd_0__inst_mult_25_32_q ;
wire Xd_0__inst_mult_25_33_q ;
wire Xd_0__inst_mult_24_32_q ;
wire Xd_0__inst_mult_24_33_q ;
wire Xd_0__inst_mult_27_32_q ;
wire Xd_0__inst_mult_27_33_q ;
wire Xd_0__inst_mult_26_32_q ;
wire Xd_0__inst_mult_26_33_q ;
wire Xd_0__inst_mult_21_32_q ;
wire Xd_0__inst_mult_21_33_q ;
wire Xd_0__inst_mult_20_32_q ;
wire Xd_0__inst_mult_20_33_q ;
wire Xd_0__inst_mult_23_32_q ;
wire Xd_0__inst_mult_23_33_q ;
wire Xd_0__inst_mult_22_32_q ;
wire Xd_0__inst_mult_22_33_q ;
wire Xd_0__inst_mult_17_32_q ;
wire Xd_0__inst_mult_17_33_q ;
wire Xd_0__inst_mult_16_32_q ;
wire Xd_0__inst_mult_16_33_q ;
wire Xd_0__inst_mult_19_32_q ;
wire Xd_0__inst_mult_19_33_q ;
wire Xd_0__inst_mult_18_32_q ;
wire Xd_0__inst_mult_18_33_q ;
wire Xd_0__inst_mult_13_32_q ;
wire Xd_0__inst_mult_13_33_q ;
wire Xd_0__inst_mult_12_32_q ;
wire Xd_0__inst_mult_12_33_q ;
wire Xd_0__inst_mult_15_32_q ;
wire Xd_0__inst_mult_15_33_q ;
wire Xd_0__inst_mult_14_32_q ;
wire Xd_0__inst_mult_14_33_q ;
wire Xd_0__inst_mult_9_32_q ;
wire Xd_0__inst_mult_9_33_q ;
wire Xd_0__inst_mult_8_32_q ;
wire Xd_0__inst_mult_8_33_q ;
wire Xd_0__inst_mult_11_32_q ;
wire Xd_0__inst_mult_11_33_q ;
wire Xd_0__inst_mult_10_32_q ;
wire Xd_0__inst_mult_10_33_q ;
wire Xd_0__inst_mult_5_32_q ;
wire Xd_0__inst_mult_5_33_q ;
wire Xd_0__inst_mult_4_32_q ;
wire Xd_0__inst_mult_4_33_q ;
wire Xd_0__inst_mult_7_32_q ;
wire Xd_0__inst_mult_7_33_q ;
wire Xd_0__inst_mult_6_32_q ;
wire Xd_0__inst_mult_6_33_q ;
wire Xd_0__inst_mult_1_32_q ;
wire Xd_0__inst_mult_1_33_q ;
wire Xd_0__inst_mult_0_32_q ;
wire Xd_0__inst_mult_0_33_q ;
wire Xd_0__inst_mult_3_32_q ;
wire Xd_0__inst_mult_3_33_q ;
wire Xd_0__inst_mult_2_32_q ;
wire Xd_0__inst_mult_2_33_q ;
wire [0:31] Xd_0__inst_sign ;
wire [0:31] Xd_0__inst_sign1 ;
wire [0:15] Xd_0__inst_r_sign ;
wire [27:0] Xd_0__inst_inst_inst_inst_dout ;


fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__16__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__18__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__19__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__20__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__21__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__22__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__23__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_121 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__24__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__24__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_121_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_126 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_inst_first_level_1__25__q ),
	.datad(!Xd_0__inst_inst_inst_first_level_0__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_126_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_127 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_131 (
// Equation(s):

	.dataa(!Xd_0__inst_inst_inst_first_level_1__26__q ),
	.datab(!Xd_0__inst_inst_inst_first_level_0__26__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_127 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_131_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_132 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_136 (
// Equation(s):

	.dataa(!Xd_0__inst_inst_inst_first_level_1__26__q ),
	.datab(!Xd_0__inst_inst_inst_first_level_0__26__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_132 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_136_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_204 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_205 ),
	.cout(Xd_0__inst_mult_2_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__0__q ),
	.datad(!Xd_0__inst_inst_first_level_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_210 ),
	.cout(Xd_0__inst_mult_2_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__1__q ),
	.datad(!Xd_0__inst_inst_first_level_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_6_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__2__q ),
	.datad(!Xd_0__inst_inst_first_level_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_11_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__3__q ),
	.datad(!Xd_0__inst_inst_first_level_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_16_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__4__q ),
	.datad(!Xd_0__inst_inst_first_level_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__5__q ),
	.datad(!Xd_0__inst_inst_first_level_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_26_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__6__q ),
	.datad(!Xd_0__inst_inst_first_level_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_31_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__7__q ),
	.datad(!Xd_0__inst_inst_first_level_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_36_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__8__q ),
	.datad(!Xd_0__inst_inst_first_level_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__9__q ),
	.datad(!Xd_0__inst_inst_first_level_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_46_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__10__q ),
	.datad(!Xd_0__inst_inst_first_level_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_51_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__11__q ),
	.datad(!Xd_0__inst_inst_first_level_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_56_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__12__q ),
	.datad(!Xd_0__inst_inst_first_level_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_66_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__14__q ),
	.datad(!Xd_0__inst_inst_first_level_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_71_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__15__q ),
	.datad(!Xd_0__inst_inst_first_level_2__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_76_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__16__q ),
	.datad(!Xd_0__inst_inst_first_level_2__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_81_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__16__q ),
	.datad(!Xd_0__inst_inst_first_level_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__17__q ),
	.datad(!Xd_0__inst_inst_first_level_2__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_86_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__17__q ),
	.datad(!Xd_0__inst_inst_first_level_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__18__q ),
	.datad(!Xd_0__inst_inst_first_level_2__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_91_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__18__q ),
	.datad(!Xd_0__inst_inst_first_level_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__19__q ),
	.datad(!Xd_0__inst_inst_first_level_2__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_96_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__19__q ),
	.datad(!Xd_0__inst_inst_first_level_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__20__q ),
	.datad(!Xd_0__inst_inst_first_level_2__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_101_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__20__q ),
	.datad(!Xd_0__inst_inst_first_level_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__21__q ),
	.datad(!Xd_0__inst_inst_first_level_2__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_106_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__21__q ),
	.datad(!Xd_0__inst_inst_first_level_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__22__q ),
	.datad(!Xd_0__inst_inst_first_level_2__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_111_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__22__q ),
	.datad(!Xd_0__inst_inst_first_level_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__23__q ),
	.datad(!Xd_0__inst_inst_first_level_2__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_116_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__23__q ),
	.datad(!Xd_0__inst_inst_first_level_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_121 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__24__q ),
	.datad(!Xd_0__inst_inst_first_level_2__24__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_121_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_121 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__24__q ),
	.datad(!Xd_0__inst_inst_first_level_0__24__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_121_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_126 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__25__q ),
	.datad(!Xd_0__inst_inst_first_level_2__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_126_sumout ),
	.cout(Xd_0__inst_inst_inst_add_1_127 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_126 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__25__q ),
	.datad(!Xd_0__inst_inst_first_level_0__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_126_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_127 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_1_131 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_3__25__q ),
	.datad(!Xd_0__inst_inst_first_level_2__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_1_127 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_1_131_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_inst_inst_add_0_131 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_inst_first_level_1__25__q ),
	.datad(!Xd_0__inst_inst_first_level_0__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_127 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_131_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_210 ),
	.datab(!Xd_0__inst_mult_26_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_205 ),
	.cout(Xd_0__inst_mult_26_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_210 ),
	.datab(!Xd_0__inst_mult_24_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_205 ),
	.cout(Xd_0__inst_mult_24_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_84 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[30]),
	.datac(!din_a[31]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_214 ),
	.cout(Xd_0__inst_mult_2_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__0__q ),
	.datad(!Xd_0__inst_r_sum2_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_1_sumout ),
	.cout(Xd_0__inst_inst_add_3_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__0__q ),
	.datad(!Xd_0__inst_r_sum2_4__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_1_sumout ),
	.cout(Xd_0__inst_inst_add_2_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_35 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[322]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_35_sumout ),
	.cout(Xd_0__inst_mult_26_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_210 ),
	.datab(!Xd_0__inst_mult_26_35_sumout ),
	.datac(!Xd_0__inst_mult_26_219 ),
	.datad(!Xd_0__inst_mult_26_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_214 ),
	.cout(Xd_0__inst_mult_26_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__0__q ),
	.datad(!Xd_0__inst_r_sum2_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_1_sumout ),
	.cout(Xd_0__inst_inst_add_1_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__0__q ),
	.datad(!Xd_0__inst_r_sum2_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_35 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[298]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_35_sumout ),
	.cout(Xd_0__inst_mult_24_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_210 ),
	.datab(!Xd_0__inst_mult_24_35_sumout ),
	.datac(!Xd_0__inst_mult_24_224 ),
	.datad(!Xd_0__inst_mult_24_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_214 ),
	.cout(Xd_0__inst_mult_24_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_85 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[30]),
	.datac(!din_a[30]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_219 ),
	.cout(Xd_0__inst_mult_2_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__1__q ),
	.datad(!Xd_0__inst_r_sum2_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_6_sumout ),
	.cout(Xd_0__inst_inst_add_3_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__1__q ),
	.datad(!Xd_0__inst_r_sum2_4__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_6_sumout ),
	.cout(Xd_0__inst_inst_add_2_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__1__q ),
	.datad(!Xd_0__inst_r_sum2_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_6_sumout ),
	.cout(Xd_0__inst_inst_add_1_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_6 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__1__q ),
	.datad(!Xd_0__inst_r_sum2_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__2__q ),
	.datad(!Xd_0__inst_r_sum2_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_11_sumout ),
	.cout(Xd_0__inst_inst_add_3_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__2__q ),
	.datad(!Xd_0__inst_r_sum2_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_11_sumout ),
	.cout(Xd_0__inst_inst_add_2_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__2__q ),
	.datad(!Xd_0__inst_r_sum2_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_11_sumout ),
	.cout(Xd_0__inst_inst_add_1_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_11 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__2__q ),
	.datad(!Xd_0__inst_r_sum2_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__3__q ),
	.datad(!Xd_0__inst_r_sum2_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_16_sumout ),
	.cout(Xd_0__inst_inst_add_3_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__3__q ),
	.datad(!Xd_0__inst_r_sum2_4__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_16_sumout ),
	.cout(Xd_0__inst_inst_add_2_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__3__q ),
	.datad(!Xd_0__inst_r_sum2_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_16_sumout ),
	.cout(Xd_0__inst_inst_add_1_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__3__q ),
	.datad(!Xd_0__inst_r_sum2_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__4__q ),
	.datad(!Xd_0__inst_r_sum2_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_21_sumout ),
	.cout(Xd_0__inst_inst_add_3_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__4__q ),
	.datad(!Xd_0__inst_r_sum2_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_21_sumout ),
	.cout(Xd_0__inst_inst_add_2_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__4__q ),
	.datad(!Xd_0__inst_r_sum2_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_21_sumout ),
	.cout(Xd_0__inst_inst_add_1_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__4__q ),
	.datad(!Xd_0__inst_r_sum2_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__5__q ),
	.datad(!Xd_0__inst_r_sum2_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_26_sumout ),
	.cout(Xd_0__inst_inst_add_3_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__5__q ),
	.datad(!Xd_0__inst_r_sum2_4__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_26_sumout ),
	.cout(Xd_0__inst_inst_add_2_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__5__q ),
	.datad(!Xd_0__inst_r_sum2_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_26_sumout ),
	.cout(Xd_0__inst_inst_add_1_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_26 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__5__q ),
	.datad(!Xd_0__inst_r_sum2_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__6__q ),
	.datad(!Xd_0__inst_r_sum2_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_31_sumout ),
	.cout(Xd_0__inst_inst_add_3_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__6__q ),
	.datad(!Xd_0__inst_r_sum2_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_31_sumout ),
	.cout(Xd_0__inst_inst_add_2_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__6__q ),
	.datad(!Xd_0__inst_r_sum2_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_31_sumout ),
	.cout(Xd_0__inst_inst_add_1_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_31 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__6__q ),
	.datad(!Xd_0__inst_r_sum2_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__7__q ),
	.datad(!Xd_0__inst_r_sum2_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_36_sumout ),
	.cout(Xd_0__inst_inst_add_3_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__7__q ),
	.datad(!Xd_0__inst_r_sum2_4__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_36_sumout ),
	.cout(Xd_0__inst_inst_add_2_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__7__q ),
	.datad(!Xd_0__inst_r_sum2_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_36_sumout ),
	.cout(Xd_0__inst_inst_add_1_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_36 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__7__q ),
	.datad(!Xd_0__inst_r_sum2_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__8__q ),
	.datad(!Xd_0__inst_r_sum2_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_41_sumout ),
	.cout(Xd_0__inst_inst_add_3_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__8__q ),
	.datad(!Xd_0__inst_r_sum2_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_41_sumout ),
	.cout(Xd_0__inst_inst_add_2_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__8__q ),
	.datad(!Xd_0__inst_r_sum2_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_41_sumout ),
	.cout(Xd_0__inst_inst_add_1_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__8__q ),
	.datad(!Xd_0__inst_r_sum2_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__9__q ),
	.datad(!Xd_0__inst_r_sum2_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_46_sumout ),
	.cout(Xd_0__inst_inst_add_3_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__9__q ),
	.datad(!Xd_0__inst_r_sum2_4__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_46_sumout ),
	.cout(Xd_0__inst_inst_add_2_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__9__q ),
	.datad(!Xd_0__inst_r_sum2_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_46_sumout ),
	.cout(Xd_0__inst_inst_add_1_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_46 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__9__q ),
	.datad(!Xd_0__inst_r_sum2_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__10__q ),
	.datad(!Xd_0__inst_r_sum2_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_51_sumout ),
	.cout(Xd_0__inst_inst_add_3_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__10__q ),
	.datad(!Xd_0__inst_r_sum2_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_51_sumout ),
	.cout(Xd_0__inst_inst_add_2_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__10__q ),
	.datad(!Xd_0__inst_r_sum2_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_51_sumout ),
	.cout(Xd_0__inst_inst_add_1_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_51 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__10__q ),
	.datad(!Xd_0__inst_r_sum2_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__11__q ),
	.datad(!Xd_0__inst_r_sum2_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_56_sumout ),
	.cout(Xd_0__inst_inst_add_3_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__11__q ),
	.datad(!Xd_0__inst_r_sum2_4__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_56_sumout ),
	.cout(Xd_0__inst_inst_add_2_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__11__q ),
	.datad(!Xd_0__inst_r_sum2_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_56_sumout ),
	.cout(Xd_0__inst_inst_add_1_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_56 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__11__q ),
	.datad(!Xd_0__inst_r_sum2_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__12__q ),
	.datad(!Xd_0__inst_r_sum2_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_61_sumout ),
	.cout(Xd_0__inst_inst_add_3_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__12__q ),
	.datad(!Xd_0__inst_r_sum2_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_61_sumout ),
	.cout(Xd_0__inst_inst_add_2_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__12__q ),
	.datad(!Xd_0__inst_r_sum2_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_61_sumout ),
	.cout(Xd_0__inst_inst_add_1_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_61 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__12__q ),
	.datad(!Xd_0__inst_r_sum2_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__13__q ),
	.datad(!Xd_0__inst_r_sum2_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_66_sumout ),
	.cout(Xd_0__inst_inst_add_3_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__13__q ),
	.datad(!Xd_0__inst_r_sum2_4__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_66_sumout ),
	.cout(Xd_0__inst_inst_add_2_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__13__q ),
	.datad(!Xd_0__inst_r_sum2_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_66_sumout ),
	.cout(Xd_0__inst_inst_add_1_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_66 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__13__q ),
	.datad(!Xd_0__inst_r_sum2_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__14__q ),
	.datad(!Xd_0__inst_r_sum2_6__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_71_sumout ),
	.cout(Xd_0__inst_inst_add_3_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__14__q ),
	.datad(!Xd_0__inst_r_sum2_4__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_71_sumout ),
	.cout(Xd_0__inst_inst_add_2_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__14__q ),
	.datad(!Xd_0__inst_r_sum2_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_71_sumout ),
	.cout(Xd_0__inst_inst_add_1_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_71 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__14__q ),
	.datad(!Xd_0__inst_r_sum2_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__15__q ),
	.datad(!Xd_0__inst_r_sum2_6__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_76_sumout ),
	.cout(Xd_0__inst_inst_add_3_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__15__q ),
	.datad(!Xd_0__inst_r_sum2_4__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_76_sumout ),
	.cout(Xd_0__inst_inst_add_2_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__15__q ),
	.datad(!Xd_0__inst_r_sum2_2__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_76_sumout ),
	.cout(Xd_0__inst_inst_add_1_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_76 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__15__q ),
	.datad(!Xd_0__inst_r_sum2_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__16__q ),
	.datad(!Xd_0__inst_r_sum2_6__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_81_sumout ),
	.cout(Xd_0__inst_inst_add_3_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__16__q ),
	.datad(!Xd_0__inst_r_sum2_4__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_81_sumout ),
	.cout(Xd_0__inst_inst_add_2_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__16__q ),
	.datad(!Xd_0__inst_r_sum2_2__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_81_sumout ),
	.cout(Xd_0__inst_inst_add_1_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_81 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__16__q ),
	.datad(!Xd_0__inst_r_sum2_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__17__q ),
	.datad(!Xd_0__inst_r_sum2_6__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_86_sumout ),
	.cout(Xd_0__inst_inst_add_3_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__17__q ),
	.datad(!Xd_0__inst_r_sum2_4__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_86_sumout ),
	.cout(Xd_0__inst_inst_add_2_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__17__q ),
	.datad(!Xd_0__inst_r_sum2_2__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_86_sumout ),
	.cout(Xd_0__inst_inst_add_1_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_86 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__17__q ),
	.datad(!Xd_0__inst_r_sum2_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__18__q ),
	.datad(!Xd_0__inst_r_sum2_6__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_91_sumout ),
	.cout(Xd_0__inst_inst_add_3_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__18__q ),
	.datad(!Xd_0__inst_r_sum2_4__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_91_sumout ),
	.cout(Xd_0__inst_inst_add_2_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__18__q ),
	.datad(!Xd_0__inst_r_sum2_2__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_91_sumout ),
	.cout(Xd_0__inst_inst_add_1_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_91 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__18__q ),
	.datad(!Xd_0__inst_r_sum2_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__19__q ),
	.datad(!Xd_0__inst_r_sum2_6__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_96_sumout ),
	.cout(Xd_0__inst_inst_add_3_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__19__q ),
	.datad(!Xd_0__inst_r_sum2_4__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_96_sumout ),
	.cout(Xd_0__inst_inst_add_2_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__19__q ),
	.datad(!Xd_0__inst_r_sum2_2__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_96_sumout ),
	.cout(Xd_0__inst_inst_add_1_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_96 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__19__q ),
	.datad(!Xd_0__inst_r_sum2_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__20__q ),
	.datad(!Xd_0__inst_r_sum2_6__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_101_sumout ),
	.cout(Xd_0__inst_inst_add_3_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__20__q ),
	.datad(!Xd_0__inst_r_sum2_4__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_101_sumout ),
	.cout(Xd_0__inst_inst_add_2_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__20__q ),
	.datad(!Xd_0__inst_r_sum2_2__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_101_sumout ),
	.cout(Xd_0__inst_inst_add_1_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_101 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__20__q ),
	.datad(!Xd_0__inst_r_sum2_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__21__q ),
	.datad(!Xd_0__inst_r_sum2_6__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_106_sumout ),
	.cout(Xd_0__inst_inst_add_3_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__21__q ),
	.datad(!Xd_0__inst_r_sum2_4__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_106_sumout ),
	.cout(Xd_0__inst_inst_add_2_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__21__q ),
	.datad(!Xd_0__inst_r_sum2_2__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_106_sumout ),
	.cout(Xd_0__inst_inst_add_1_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__21__q ),
	.datad(!Xd_0__inst_r_sum2_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__22__q ),
	.datad(!Xd_0__inst_r_sum2_6__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_111_sumout ),
	.cout(Xd_0__inst_inst_add_3_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__22__q ),
	.datad(!Xd_0__inst_r_sum2_4__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_111_sumout ),
	.cout(Xd_0__inst_inst_add_2_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__22__q ),
	.datad(!Xd_0__inst_r_sum2_2__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_111_sumout ),
	.cout(Xd_0__inst_inst_add_1_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_111 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__22__q ),
	.datad(!Xd_0__inst_r_sum2_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_7__23__q ),
	.datad(!Xd_0__inst_r_sum2_6__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_116_sumout ),
	.cout(Xd_0__inst_inst_add_3_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_5__23__q ),
	.datad(!Xd_0__inst_r_sum2_4__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_116_sumout ),
	.cout(Xd_0__inst_inst_add_2_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_3__23__q ),
	.datad(!Xd_0__inst_r_sum2_2__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_116_sumout ),
	.cout(Xd_0__inst_inst_add_1_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000F0FF0),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum2_1__23__q ),
	.datad(!Xd_0__inst_r_sum2_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_7__24__q ),
	.datab(!Xd_0__inst_r_sum2_6__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_121_sumout ),
	.cout(Xd_0__inst_inst_add_3_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_5__24__q ),
	.datab(!Xd_0__inst_r_sum2_4__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_121_sumout ),
	.cout(Xd_0__inst_inst_add_2_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_3__24__q ),
	.datab(!Xd_0__inst_r_sum2_2__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_121_sumout ),
	.cout(Xd_0__inst_inst_add_1_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_1__24__q ),
	.datab(!Xd_0__inst_r_sum2_0__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_121_sumout ),
	.cout(Xd_0__inst_inst_add_0_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_3_126 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_7__24__q ),
	.datab(!Xd_0__inst_r_sum2_6__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_3_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_3_126_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_2_126 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_5__24__q ),
	.datab(!Xd_0__inst_r_sum2_4__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_2_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_126_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_1_126 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_3__24__q ),
	.datab(!Xd_0__inst_r_sum2_2__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_1_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_1_126_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_inst_add_0_126 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum2_1__24__q ),
	.datab(!Xd_0__inst_r_sum2_0__24__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_inst_add_0_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_126_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_210 ),
	.datab(!Xd_0__inst_mult_25_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_205 ),
	.cout(Xd_0__inst_mult_25_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_234 ),
	.datab(!Xd_0__inst_mult_24_45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_219 ),
	.cout(Xd_0__inst_mult_24_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_85 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[322]),
	.datac(!Xd_0__inst_mult_26_234 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_219 ),
	.cout(Xd_0__inst_mult_26_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_35 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[334]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_35_sumout ),
	.cout(Xd_0__inst_mult_27_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_40 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[321]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_40_sumout ),
	.cout(Xd_0__inst_mult_26_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_219 ),
	.datab(!Xd_0__inst_mult_26_40_sumout ),
	.datac(!Xd_0__inst_mult_26_244 ),
	.datad(!Xd_0__inst_mult_26_239 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_224 ),
	.cout(Xd_0__inst_mult_26_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_210 ),
	.datab(!Xd_0__inst_mult_27_45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_205 ),
	.cout(Xd_0__inst_mult_27_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_254 ),
	.datab(!Xd_0__inst_mult_26_45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_229 ),
	.cout(Xd_0__inst_mult_26_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_86 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[298]),
	.datac(!Xd_0__inst_mult_24_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_224 ),
	.cout(Xd_0__inst_mult_24_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_40 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[297]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_40_sumout ),
	.cout(Xd_0__inst_mult_24_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_224 ),
	.datab(!Xd_0__inst_mult_24_40_sumout ),
	.datac(!Xd_0__inst_mult_24_254 ),
	.datad(!Xd_0__inst_mult_24_249 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_229 ),
	.cout(Xd_0__inst_mult_24_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_86 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(!din_a[29]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_224 ),
	.cout(Xd_0__inst_mult_2_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_15__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_14__0__q ),
	.datad(!Xd_0__inst_r_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_13__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_12__0__q ),
	.datad(!Xd_0__inst_r_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_35 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[304]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_35_sumout ),
	.cout(Xd_0__inst_mult_25_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_210 ),
	.datab(!Xd_0__inst_mult_25_35_sumout ),
	.datac(!Xd_0__inst_mult_25_219 ),
	.datad(!Xd_0__inst_mult_25_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_214 ),
	.cout(Xd_0__inst_mult_25_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_11__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_10__0__q ),
	.datad(!Xd_0__inst_r_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_9__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_8__0__q ),
	.datad(!Xd_0__inst_r_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_88 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_234 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_45 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[292]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_45_sumout ),
	.cout(Xd_0__inst_mult_24_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_234 ),
	.datab(!Xd_0__inst_mult_24_45_sumout ),
	.datac(!Xd_0__inst_mult_24_264 ),
	.datad(!Xd_0__inst_mult_24_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_239 ),
	.cout(Xd_0__inst_mult_24_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_26_88 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[321]),
	.datac(!din_a[313]),
	.datad(!din_b[320]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_234 ),
	.cout(Xd_0__inst_mult_26_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_89 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[321]),
	.datac(!Xd_0__inst_mult_26_264 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_239 ),
	.cout(Xd_0__inst_mult_26_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_40 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[333]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_40_sumout ),
	.cout(Xd_0__inst_mult_27_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_90 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_244 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_244 ),
	.datab(!Xd_0__inst_mult_26_239 ),
	.datac(!din_a[321]),
	.datad(!din_b[320]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_249 ),
	.cout(Xd_0__inst_mult_26_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_7__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_6__0__q ),
	.datad(!Xd_0__inst_r_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_5__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_45 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[328]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_45_sumout ),
	.cout(Xd_0__inst_mult_27_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_210 ),
	.datab(!Xd_0__inst_mult_27_45_sumout ),
	.datac(!Xd_0__inst_mult_27_219 ),
	.datad(!Xd_0__inst_mult_27_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_214 ),
	.cout(Xd_0__inst_mult_27_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_3__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_2__0__q ),
	.datad(!Xd_0__inst_r_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000005A5AA5),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_1__0__q ),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sum1_0__0__q ),
	.datad(!Xd_0__inst_r_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_127_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_92 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_254 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_45 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[316]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_45_sumout ),
	.cout(Xd_0__inst_mult_26_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_254 ),
	.datab(!Xd_0__inst_mult_26_45_sumout ),
	.datac(!Xd_0__inst_mult_26_284 ),
	.datad(!Xd_0__inst_mult_26_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_259 ),
	.cout(Xd_0__inst_mult_26_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_24_90 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[297]),
	.datac(!din_a[289]),
	.datad(!din_b[296]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_244 ),
	.cout(Xd_0__inst_mult_24_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_91 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[297]),
	.datac(!Xd_0__inst_mult_24_274 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_249 ),
	.cout(Xd_0__inst_mult_24_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_40 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[309]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_40_sumout ),
	.cout(Xd_0__inst_mult_25_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_92 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_254 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_254 ),
	.datab(!Xd_0__inst_mult_24_249 ),
	.datac(!din_a[297]),
	.datad(!din_b[296]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_259 ),
	.cout(Xd_0__inst_mult_24_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_87 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[30]),
	.datac(!din_a[28]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_229 ),
	.cout(Xd_0__inst_mult_2_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__1__q ),
	.datab(!Xd_0__inst_r_sum1_15__1__q ),
	.datac(!Xd_0__inst_r_sum1_15__0__q ),
	.datad(!Xd_0__inst_r_sum1_14__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__1__q ),
	.datab(!Xd_0__inst_r_sum1_13__1__q ),
	.datac(!Xd_0__inst_r_sum1_13__0__q ),
	.datad(!Xd_0__inst_r_sum1_12__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__1__q ),
	.datab(!Xd_0__inst_r_sum1_11__1__q ),
	.datac(!Xd_0__inst_r_sum1_11__0__q ),
	.datad(!Xd_0__inst_r_sum1_10__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__1__q ),
	.datab(!Xd_0__inst_r_sum1_9__1__q ),
	.datac(!Xd_0__inst_r_sum1_9__0__q ),
	.datad(!Xd_0__inst_r_sum1_8__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__1__q ),
	.datab(!Xd_0__inst_r_sum1_7__1__q ),
	.datac(!Xd_0__inst_r_sum1_7__0__q ),
	.datad(!Xd_0__inst_r_sum1_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__1__q ),
	.datab(!Xd_0__inst_r_sum1_5__1__q ),
	.datac(!Xd_0__inst_r_sum1_5__0__q ),
	.datad(!Xd_0__inst_r_sum1_4__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__1__q ),
	.datab(!Xd_0__inst_r_sum1_3__1__q ),
	.datac(!Xd_0__inst_r_sum1_3__0__q ),
	.datad(!Xd_0__inst_r_sum1_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__1__q ),
	.datab(!Xd_0__inst_r_sum1_1__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__0__q ),
	.datad(!Xd_0__inst_r_sum1_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__1__q ),
	.datab(!Xd_0__inst_r_sum1_15__1__q ),
	.datac(!Xd_0__inst_r_sum1_14__2__q ),
	.datad(!Xd_0__inst_r_sum1_15__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__1__q ),
	.datab(!Xd_0__inst_r_sum1_13__1__q ),
	.datac(!Xd_0__inst_r_sum1_12__2__q ),
	.datad(!Xd_0__inst_r_sum1_13__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__1__q ),
	.datab(!Xd_0__inst_r_sum1_11__1__q ),
	.datac(!Xd_0__inst_r_sum1_10__2__q ),
	.datad(!Xd_0__inst_r_sum1_11__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__1__q ),
	.datab(!Xd_0__inst_r_sum1_9__1__q ),
	.datac(!Xd_0__inst_r_sum1_8__2__q ),
	.datad(!Xd_0__inst_r_sum1_9__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__1__q ),
	.datab(!Xd_0__inst_r_sum1_7__1__q ),
	.datac(!Xd_0__inst_r_sum1_6__2__q ),
	.datad(!Xd_0__inst_r_sum1_7__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__1__q ),
	.datab(!Xd_0__inst_r_sum1_5__1__q ),
	.datac(!Xd_0__inst_r_sum1_4__2__q ),
	.datad(!Xd_0__inst_r_sum1_5__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__1__q ),
	.datab(!Xd_0__inst_r_sum1_3__1__q ),
	.datac(!Xd_0__inst_r_sum1_2__2__q ),
	.datad(!Xd_0__inst_r_sum1_3__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__1__q ),
	.datab(!Xd_0__inst_r_sum1_1__1__q ),
	.datac(!Xd_0__inst_r_sum1_0__2__q ),
	.datad(!Xd_0__inst_r_sum1_1__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__3__q ),
	.datab(!Xd_0__inst_r_sum1_15__3__q ),
	.datac(!Xd_0__inst_r_sum1_15__2__q ),
	.datad(!Xd_0__inst_r_sum1_14__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__3__q ),
	.datab(!Xd_0__inst_r_sum1_13__3__q ),
	.datac(!Xd_0__inst_r_sum1_13__2__q ),
	.datad(!Xd_0__inst_r_sum1_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__3__q ),
	.datab(!Xd_0__inst_r_sum1_11__3__q ),
	.datac(!Xd_0__inst_r_sum1_11__2__q ),
	.datad(!Xd_0__inst_r_sum1_10__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__3__q ),
	.datab(!Xd_0__inst_r_sum1_9__3__q ),
	.datac(!Xd_0__inst_r_sum1_9__2__q ),
	.datad(!Xd_0__inst_r_sum1_8__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__3__q ),
	.datab(!Xd_0__inst_r_sum1_7__3__q ),
	.datac(!Xd_0__inst_r_sum1_7__2__q ),
	.datad(!Xd_0__inst_r_sum1_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__3__q ),
	.datab(!Xd_0__inst_r_sum1_5__3__q ),
	.datac(!Xd_0__inst_r_sum1_5__2__q ),
	.datad(!Xd_0__inst_r_sum1_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__3__q ),
	.datab(!Xd_0__inst_r_sum1_3__3__q ),
	.datac(!Xd_0__inst_r_sum1_3__2__q ),
	.datad(!Xd_0__inst_r_sum1_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__3__q ),
	.datab(!Xd_0__inst_r_sum1_1__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__3__q ),
	.datab(!Xd_0__inst_r_sum1_15__3__q ),
	.datac(!Xd_0__inst_r_sum1_14__4__q ),
	.datad(!Xd_0__inst_r_sum1_15__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__3__q ),
	.datab(!Xd_0__inst_r_sum1_13__3__q ),
	.datac(!Xd_0__inst_r_sum1_12__4__q ),
	.datad(!Xd_0__inst_r_sum1_13__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__3__q ),
	.datab(!Xd_0__inst_r_sum1_11__3__q ),
	.datac(!Xd_0__inst_r_sum1_10__4__q ),
	.datad(!Xd_0__inst_r_sum1_11__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__3__q ),
	.datab(!Xd_0__inst_r_sum1_9__3__q ),
	.datac(!Xd_0__inst_r_sum1_8__4__q ),
	.datad(!Xd_0__inst_r_sum1_9__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__3__q ),
	.datab(!Xd_0__inst_r_sum1_7__3__q ),
	.datac(!Xd_0__inst_r_sum1_6__4__q ),
	.datad(!Xd_0__inst_r_sum1_7__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__3__q ),
	.datab(!Xd_0__inst_r_sum1_5__3__q ),
	.datac(!Xd_0__inst_r_sum1_4__4__q ),
	.datad(!Xd_0__inst_r_sum1_5__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__3__q ),
	.datab(!Xd_0__inst_r_sum1_3__3__q ),
	.datac(!Xd_0__inst_r_sum1_2__4__q ),
	.datad(!Xd_0__inst_r_sum1_3__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__3__q ),
	.datab(!Xd_0__inst_r_sum1_1__3__q ),
	.datac(!Xd_0__inst_r_sum1_0__4__q ),
	.datad(!Xd_0__inst_r_sum1_1__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__5__q ),
	.datab(!Xd_0__inst_r_sum1_15__5__q ),
	.datac(!Xd_0__inst_r_sum1_15__4__q ),
	.datad(!Xd_0__inst_r_sum1_14__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__5__q ),
	.datab(!Xd_0__inst_r_sum1_13__5__q ),
	.datac(!Xd_0__inst_r_sum1_13__4__q ),
	.datad(!Xd_0__inst_r_sum1_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__5__q ),
	.datab(!Xd_0__inst_r_sum1_11__5__q ),
	.datac(!Xd_0__inst_r_sum1_11__4__q ),
	.datad(!Xd_0__inst_r_sum1_10__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__5__q ),
	.datab(!Xd_0__inst_r_sum1_9__5__q ),
	.datac(!Xd_0__inst_r_sum1_9__4__q ),
	.datad(!Xd_0__inst_r_sum1_8__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__5__q ),
	.datab(!Xd_0__inst_r_sum1_7__5__q ),
	.datac(!Xd_0__inst_r_sum1_7__4__q ),
	.datad(!Xd_0__inst_r_sum1_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__5__q ),
	.datab(!Xd_0__inst_r_sum1_5__5__q ),
	.datac(!Xd_0__inst_r_sum1_5__4__q ),
	.datad(!Xd_0__inst_r_sum1_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__5__q ),
	.datab(!Xd_0__inst_r_sum1_3__5__q ),
	.datac(!Xd_0__inst_r_sum1_3__4__q ),
	.datad(!Xd_0__inst_r_sum1_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__5__q ),
	.datab(!Xd_0__inst_r_sum1_1__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__5__q ),
	.datab(!Xd_0__inst_r_sum1_15__5__q ),
	.datac(!Xd_0__inst_r_sum1_14__6__q ),
	.datad(!Xd_0__inst_r_sum1_15__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__5__q ),
	.datab(!Xd_0__inst_r_sum1_13__5__q ),
	.datac(!Xd_0__inst_r_sum1_12__6__q ),
	.datad(!Xd_0__inst_r_sum1_13__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__5__q ),
	.datab(!Xd_0__inst_r_sum1_11__5__q ),
	.datac(!Xd_0__inst_r_sum1_10__6__q ),
	.datad(!Xd_0__inst_r_sum1_11__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__5__q ),
	.datab(!Xd_0__inst_r_sum1_9__5__q ),
	.datac(!Xd_0__inst_r_sum1_8__6__q ),
	.datad(!Xd_0__inst_r_sum1_9__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__5__q ),
	.datab(!Xd_0__inst_r_sum1_7__5__q ),
	.datac(!Xd_0__inst_r_sum1_6__6__q ),
	.datad(!Xd_0__inst_r_sum1_7__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__5__q ),
	.datab(!Xd_0__inst_r_sum1_5__5__q ),
	.datac(!Xd_0__inst_r_sum1_4__6__q ),
	.datad(!Xd_0__inst_r_sum1_5__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__5__q ),
	.datab(!Xd_0__inst_r_sum1_3__5__q ),
	.datac(!Xd_0__inst_r_sum1_2__6__q ),
	.datad(!Xd_0__inst_r_sum1_3__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__5__q ),
	.datab(!Xd_0__inst_r_sum1_1__5__q ),
	.datac(!Xd_0__inst_r_sum1_0__6__q ),
	.datad(!Xd_0__inst_r_sum1_1__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__7__q ),
	.datab(!Xd_0__inst_r_sum1_15__7__q ),
	.datac(!Xd_0__inst_r_sum1_15__6__q ),
	.datad(!Xd_0__inst_r_sum1_14__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__7__q ),
	.datab(!Xd_0__inst_r_sum1_13__7__q ),
	.datac(!Xd_0__inst_r_sum1_13__6__q ),
	.datad(!Xd_0__inst_r_sum1_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__7__q ),
	.datab(!Xd_0__inst_r_sum1_11__7__q ),
	.datac(!Xd_0__inst_r_sum1_11__6__q ),
	.datad(!Xd_0__inst_r_sum1_10__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__7__q ),
	.datab(!Xd_0__inst_r_sum1_9__7__q ),
	.datac(!Xd_0__inst_r_sum1_9__6__q ),
	.datad(!Xd_0__inst_r_sum1_8__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__7__q ),
	.datab(!Xd_0__inst_r_sum1_7__7__q ),
	.datac(!Xd_0__inst_r_sum1_7__6__q ),
	.datad(!Xd_0__inst_r_sum1_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__7__q ),
	.datab(!Xd_0__inst_r_sum1_5__7__q ),
	.datac(!Xd_0__inst_r_sum1_5__6__q ),
	.datad(!Xd_0__inst_r_sum1_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__7__q ),
	.datab(!Xd_0__inst_r_sum1_3__7__q ),
	.datac(!Xd_0__inst_r_sum1_3__6__q ),
	.datad(!Xd_0__inst_r_sum1_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__7__q ),
	.datab(!Xd_0__inst_r_sum1_1__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__7__q ),
	.datab(!Xd_0__inst_r_sum1_15__7__q ),
	.datac(!Xd_0__inst_r_sum1_14__8__q ),
	.datad(!Xd_0__inst_r_sum1_15__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__7__q ),
	.datab(!Xd_0__inst_r_sum1_13__7__q ),
	.datac(!Xd_0__inst_r_sum1_12__8__q ),
	.datad(!Xd_0__inst_r_sum1_13__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__7__q ),
	.datab(!Xd_0__inst_r_sum1_11__7__q ),
	.datac(!Xd_0__inst_r_sum1_10__8__q ),
	.datad(!Xd_0__inst_r_sum1_11__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__7__q ),
	.datab(!Xd_0__inst_r_sum1_9__7__q ),
	.datac(!Xd_0__inst_r_sum1_8__8__q ),
	.datad(!Xd_0__inst_r_sum1_9__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__7__q ),
	.datab(!Xd_0__inst_r_sum1_7__7__q ),
	.datac(!Xd_0__inst_r_sum1_6__8__q ),
	.datad(!Xd_0__inst_r_sum1_7__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__7__q ),
	.datab(!Xd_0__inst_r_sum1_5__7__q ),
	.datac(!Xd_0__inst_r_sum1_4__8__q ),
	.datad(!Xd_0__inst_r_sum1_5__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__7__q ),
	.datab(!Xd_0__inst_r_sum1_3__7__q ),
	.datac(!Xd_0__inst_r_sum1_2__8__q ),
	.datad(!Xd_0__inst_r_sum1_3__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__7__q ),
	.datab(!Xd_0__inst_r_sum1_1__7__q ),
	.datac(!Xd_0__inst_r_sum1_0__8__q ),
	.datad(!Xd_0__inst_r_sum1_1__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__9__q ),
	.datab(!Xd_0__inst_r_sum1_15__9__q ),
	.datac(!Xd_0__inst_r_sum1_15__8__q ),
	.datad(!Xd_0__inst_r_sum1_14__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__9__q ),
	.datab(!Xd_0__inst_r_sum1_13__9__q ),
	.datac(!Xd_0__inst_r_sum1_13__8__q ),
	.datad(!Xd_0__inst_r_sum1_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__9__q ),
	.datab(!Xd_0__inst_r_sum1_11__9__q ),
	.datac(!Xd_0__inst_r_sum1_11__8__q ),
	.datad(!Xd_0__inst_r_sum1_10__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__9__q ),
	.datab(!Xd_0__inst_r_sum1_9__9__q ),
	.datac(!Xd_0__inst_r_sum1_9__8__q ),
	.datad(!Xd_0__inst_r_sum1_8__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__9__q ),
	.datab(!Xd_0__inst_r_sum1_7__9__q ),
	.datac(!Xd_0__inst_r_sum1_7__8__q ),
	.datad(!Xd_0__inst_r_sum1_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__9__q ),
	.datab(!Xd_0__inst_r_sum1_5__9__q ),
	.datac(!Xd_0__inst_r_sum1_5__8__q ),
	.datad(!Xd_0__inst_r_sum1_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__9__q ),
	.datab(!Xd_0__inst_r_sum1_3__9__q ),
	.datac(!Xd_0__inst_r_sum1_3__8__q ),
	.datad(!Xd_0__inst_r_sum1_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__9__q ),
	.datab(!Xd_0__inst_r_sum1_1__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__9__q ),
	.datab(!Xd_0__inst_r_sum1_15__9__q ),
	.datac(!Xd_0__inst_r_sum1_14__10__q ),
	.datad(!Xd_0__inst_r_sum1_15__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__9__q ),
	.datab(!Xd_0__inst_r_sum1_13__9__q ),
	.datac(!Xd_0__inst_r_sum1_12__10__q ),
	.datad(!Xd_0__inst_r_sum1_13__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__9__q ),
	.datab(!Xd_0__inst_r_sum1_11__9__q ),
	.datac(!Xd_0__inst_r_sum1_10__10__q ),
	.datad(!Xd_0__inst_r_sum1_11__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__9__q ),
	.datab(!Xd_0__inst_r_sum1_9__9__q ),
	.datac(!Xd_0__inst_r_sum1_8__10__q ),
	.datad(!Xd_0__inst_r_sum1_9__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__9__q ),
	.datab(!Xd_0__inst_r_sum1_7__9__q ),
	.datac(!Xd_0__inst_r_sum1_6__10__q ),
	.datad(!Xd_0__inst_r_sum1_7__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__9__q ),
	.datab(!Xd_0__inst_r_sum1_5__9__q ),
	.datac(!Xd_0__inst_r_sum1_4__10__q ),
	.datad(!Xd_0__inst_r_sum1_5__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__9__q ),
	.datab(!Xd_0__inst_r_sum1_3__9__q ),
	.datac(!Xd_0__inst_r_sum1_2__10__q ),
	.datad(!Xd_0__inst_r_sum1_3__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__9__q ),
	.datab(!Xd_0__inst_r_sum1_1__9__q ),
	.datac(!Xd_0__inst_r_sum1_0__10__q ),
	.datad(!Xd_0__inst_r_sum1_1__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__11__q ),
	.datab(!Xd_0__inst_r_sum1_15__11__q ),
	.datac(!Xd_0__inst_r_sum1_15__10__q ),
	.datad(!Xd_0__inst_r_sum1_14__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__11__q ),
	.datab(!Xd_0__inst_r_sum1_13__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__10__q ),
	.datad(!Xd_0__inst_r_sum1_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__11__q ),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_11__10__q ),
	.datad(!Xd_0__inst_r_sum1_10__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__11__q ),
	.datab(!Xd_0__inst_r_sum1_9__11__q ),
	.datac(!Xd_0__inst_r_sum1_9__10__q ),
	.datad(!Xd_0__inst_r_sum1_8__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__11__q ),
	.datab(!Xd_0__inst_r_sum1_7__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__10__q ),
	.datad(!Xd_0__inst_r_sum1_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__11__q ),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_5__10__q ),
	.datad(!Xd_0__inst_r_sum1_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__11__q ),
	.datab(!Xd_0__inst_r_sum1_3__11__q ),
	.datac(!Xd_0__inst_r_sum1_3__10__q ),
	.datad(!Xd_0__inst_r_sum1_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__11__q ),
	.datab(!Xd_0__inst_r_sum1_1__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__11__q ),
	.datab(!Xd_0__inst_r_sum1_15__11__q ),
	.datac(!Xd_0__inst_r_sum1_14__12__q ),
	.datad(!Xd_0__inst_r_sum1_15__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__11__q ),
	.datab(!Xd_0__inst_r_sum1_13__11__q ),
	.datac(!Xd_0__inst_r_sum1_12__12__q ),
	.datad(!Xd_0__inst_r_sum1_13__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__11__q ),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__12__q ),
	.datad(!Xd_0__inst_r_sum1_11__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__11__q ),
	.datab(!Xd_0__inst_r_sum1_9__11__q ),
	.datac(!Xd_0__inst_r_sum1_8__12__q ),
	.datad(!Xd_0__inst_r_sum1_9__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__11__q ),
	.datab(!Xd_0__inst_r_sum1_7__11__q ),
	.datac(!Xd_0__inst_r_sum1_6__12__q ),
	.datad(!Xd_0__inst_r_sum1_7__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__11__q ),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__12__q ),
	.datad(!Xd_0__inst_r_sum1_5__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__11__q ),
	.datab(!Xd_0__inst_r_sum1_3__11__q ),
	.datac(!Xd_0__inst_r_sum1_2__12__q ),
	.datad(!Xd_0__inst_r_sum1_3__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__11__q ),
	.datab(!Xd_0__inst_r_sum1_1__11__q ),
	.datac(!Xd_0__inst_r_sum1_0__12__q ),
	.datad(!Xd_0__inst_r_sum1_1__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__13__q ),
	.datab(!Xd_0__inst_r_sum1_15__13__q ),
	.datac(!Xd_0__inst_r_sum1_15__12__q ),
	.datad(!Xd_0__inst_r_sum1_14__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__13__q ),
	.datab(!Xd_0__inst_r_sum1_13__13__q ),
	.datac(!Xd_0__inst_r_sum1_13__12__q ),
	.datad(!Xd_0__inst_r_sum1_12__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__13__q ),
	.datab(!Xd_0__inst_r_sum1_11__13__q ),
	.datac(!Xd_0__inst_r_sum1_11__12__q ),
	.datad(!Xd_0__inst_r_sum1_10__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__13__q ),
	.datab(!Xd_0__inst_r_sum1_9__13__q ),
	.datac(!Xd_0__inst_r_sum1_9__12__q ),
	.datad(!Xd_0__inst_r_sum1_8__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__13__q ),
	.datab(!Xd_0__inst_r_sum1_7__13__q ),
	.datac(!Xd_0__inst_r_sum1_7__12__q ),
	.datad(!Xd_0__inst_r_sum1_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__13__q ),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_5__12__q ),
	.datad(!Xd_0__inst_r_sum1_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__13__q ),
	.datab(!Xd_0__inst_r_sum1_3__13__q ),
	.datac(!Xd_0__inst_r_sum1_3__12__q ),
	.datad(!Xd_0__inst_r_sum1_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__13__q ),
	.datab(!Xd_0__inst_r_sum1_1__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__12__q ),
	.datad(!Xd_0__inst_r_sum1_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__13__q ),
	.datab(!Xd_0__inst_r_sum1_15__13__q ),
	.datac(!Xd_0__inst_r_sum1_14__14__q ),
	.datad(!Xd_0__inst_r_sum1_15__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__13__q ),
	.datab(!Xd_0__inst_r_sum1_13__13__q ),
	.datac(!Xd_0__inst_r_sum1_12__14__q ),
	.datad(!Xd_0__inst_r_sum1_13__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__13__q ),
	.datab(!Xd_0__inst_r_sum1_11__13__q ),
	.datac(!Xd_0__inst_r_sum1_10__14__q ),
	.datad(!Xd_0__inst_r_sum1_11__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__13__q ),
	.datab(!Xd_0__inst_r_sum1_9__13__q ),
	.datac(!Xd_0__inst_r_sum1_8__14__q ),
	.datad(!Xd_0__inst_r_sum1_9__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__13__q ),
	.datab(!Xd_0__inst_r_sum1_7__13__q ),
	.datac(!Xd_0__inst_r_sum1_6__14__q ),
	.datad(!Xd_0__inst_r_sum1_7__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__13__q ),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__14__q ),
	.datad(!Xd_0__inst_r_sum1_5__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__13__q ),
	.datab(!Xd_0__inst_r_sum1_3__13__q ),
	.datac(!Xd_0__inst_r_sum1_2__14__q ),
	.datad(!Xd_0__inst_r_sum1_3__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__13__q ),
	.datab(!Xd_0__inst_r_sum1_1__13__q ),
	.datac(!Xd_0__inst_r_sum1_0__14__q ),
	.datad(!Xd_0__inst_r_sum1_1__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__15__q ),
	.datab(!Xd_0__inst_r_sum1_15__15__q ),
	.datac(!Xd_0__inst_r_sum1_15__14__q ),
	.datad(!Xd_0__inst_r_sum1_14__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__15__q ),
	.datab(!Xd_0__inst_r_sum1_13__15__q ),
	.datac(!Xd_0__inst_r_sum1_13__14__q ),
	.datad(!Xd_0__inst_r_sum1_12__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__15__q ),
	.datab(!Xd_0__inst_r_sum1_11__15__q ),
	.datac(!Xd_0__inst_r_sum1_11__14__q ),
	.datad(!Xd_0__inst_r_sum1_10__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__15__q ),
	.datab(!Xd_0__inst_r_sum1_9__15__q ),
	.datac(!Xd_0__inst_r_sum1_9__14__q ),
	.datad(!Xd_0__inst_r_sum1_8__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__15__q ),
	.datab(!Xd_0__inst_r_sum1_7__15__q ),
	.datac(!Xd_0__inst_r_sum1_7__14__q ),
	.datad(!Xd_0__inst_r_sum1_6__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__15__q ),
	.datab(!Xd_0__inst_r_sum1_5__15__q ),
	.datac(!Xd_0__inst_r_sum1_5__14__q ),
	.datad(!Xd_0__inst_r_sum1_4__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__15__q ),
	.datab(!Xd_0__inst_r_sum1_3__15__q ),
	.datac(!Xd_0__inst_r_sum1_3__14__q ),
	.datad(!Xd_0__inst_r_sum1_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__15__q ),
	.datab(!Xd_0__inst_r_sum1_1__15__q ),
	.datac(!Xd_0__inst_r_sum1_1__14__q ),
	.datad(!Xd_0__inst_r_sum1_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__15__q ),
	.datab(!Xd_0__inst_r_sum1_15__15__q ),
	.datac(!Xd_0__inst_r_sum1_14__16__q ),
	.datad(!Xd_0__inst_r_sum1_15__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__15__q ),
	.datab(!Xd_0__inst_r_sum1_13__15__q ),
	.datac(!Xd_0__inst_r_sum1_12__16__q ),
	.datad(!Xd_0__inst_r_sum1_13__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__15__q ),
	.datab(!Xd_0__inst_r_sum1_11__15__q ),
	.datac(!Xd_0__inst_r_sum1_10__16__q ),
	.datad(!Xd_0__inst_r_sum1_11__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__15__q ),
	.datab(!Xd_0__inst_r_sum1_9__15__q ),
	.datac(!Xd_0__inst_r_sum1_8__16__q ),
	.datad(!Xd_0__inst_r_sum1_9__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__15__q ),
	.datab(!Xd_0__inst_r_sum1_7__15__q ),
	.datac(!Xd_0__inst_r_sum1_6__16__q ),
	.datad(!Xd_0__inst_r_sum1_7__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__15__q ),
	.datab(!Xd_0__inst_r_sum1_5__15__q ),
	.datac(!Xd_0__inst_r_sum1_4__16__q ),
	.datad(!Xd_0__inst_r_sum1_5__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__15__q ),
	.datab(!Xd_0__inst_r_sum1_3__15__q ),
	.datac(!Xd_0__inst_r_sum1_2__16__q ),
	.datad(!Xd_0__inst_r_sum1_3__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__15__q ),
	.datab(!Xd_0__inst_r_sum1_1__15__q ),
	.datac(!Xd_0__inst_r_sum1_0__16__q ),
	.datad(!Xd_0__inst_r_sum1_1__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__17__q ),
	.datab(!Xd_0__inst_r_sum1_15__17__q ),
	.datac(!Xd_0__inst_r_sum1_15__16__q ),
	.datad(!Xd_0__inst_r_sum1_14__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__17__q ),
	.datab(!Xd_0__inst_r_sum1_13__17__q ),
	.datac(!Xd_0__inst_r_sum1_13__16__q ),
	.datad(!Xd_0__inst_r_sum1_12__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__17__q ),
	.datab(!Xd_0__inst_r_sum1_11__17__q ),
	.datac(!Xd_0__inst_r_sum1_11__16__q ),
	.datad(!Xd_0__inst_r_sum1_10__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__17__q ),
	.datab(!Xd_0__inst_r_sum1_9__17__q ),
	.datac(!Xd_0__inst_r_sum1_9__16__q ),
	.datad(!Xd_0__inst_r_sum1_8__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__17__q ),
	.datab(!Xd_0__inst_r_sum1_7__17__q ),
	.datac(!Xd_0__inst_r_sum1_7__16__q ),
	.datad(!Xd_0__inst_r_sum1_6__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__17__q ),
	.datab(!Xd_0__inst_r_sum1_5__17__q ),
	.datac(!Xd_0__inst_r_sum1_5__16__q ),
	.datad(!Xd_0__inst_r_sum1_4__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__17__q ),
	.datab(!Xd_0__inst_r_sum1_3__17__q ),
	.datac(!Xd_0__inst_r_sum1_3__16__q ),
	.datad(!Xd_0__inst_r_sum1_2__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__17__q ),
	.datab(!Xd_0__inst_r_sum1_1__17__q ),
	.datac(!Xd_0__inst_r_sum1_1__16__q ),
	.datad(!Xd_0__inst_r_sum1_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__17__q ),
	.datab(!Xd_0__inst_r_sum1_15__17__q ),
	.datac(!Xd_0__inst_r_sum1_14__18__q ),
	.datad(!Xd_0__inst_r_sum1_15__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__17__q ),
	.datab(!Xd_0__inst_r_sum1_13__17__q ),
	.datac(!Xd_0__inst_r_sum1_12__18__q ),
	.datad(!Xd_0__inst_r_sum1_13__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__17__q ),
	.datab(!Xd_0__inst_r_sum1_11__17__q ),
	.datac(!Xd_0__inst_r_sum1_10__18__q ),
	.datad(!Xd_0__inst_r_sum1_11__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__17__q ),
	.datab(!Xd_0__inst_r_sum1_9__17__q ),
	.datac(!Xd_0__inst_r_sum1_8__18__q ),
	.datad(!Xd_0__inst_r_sum1_9__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__17__q ),
	.datab(!Xd_0__inst_r_sum1_7__17__q ),
	.datac(!Xd_0__inst_r_sum1_6__18__q ),
	.datad(!Xd_0__inst_r_sum1_7__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__17__q ),
	.datab(!Xd_0__inst_r_sum1_5__17__q ),
	.datac(!Xd_0__inst_r_sum1_4__18__q ),
	.datad(!Xd_0__inst_r_sum1_5__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__17__q ),
	.datab(!Xd_0__inst_r_sum1_3__17__q ),
	.datac(!Xd_0__inst_r_sum1_2__18__q ),
	.datad(!Xd_0__inst_r_sum1_3__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__17__q ),
	.datab(!Xd_0__inst_r_sum1_1__17__q ),
	.datac(!Xd_0__inst_r_sum1_0__18__q ),
	.datad(!Xd_0__inst_r_sum1_1__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__19__q ),
	.datab(!Xd_0__inst_r_sum1_15__19__q ),
	.datac(!Xd_0__inst_r_sum1_15__18__q ),
	.datad(!Xd_0__inst_r_sum1_14__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__19__q ),
	.datab(!Xd_0__inst_r_sum1_13__19__q ),
	.datac(!Xd_0__inst_r_sum1_13__18__q ),
	.datad(!Xd_0__inst_r_sum1_12__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__19__q ),
	.datab(!Xd_0__inst_r_sum1_11__19__q ),
	.datac(!Xd_0__inst_r_sum1_11__18__q ),
	.datad(!Xd_0__inst_r_sum1_10__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__19__q ),
	.datab(!Xd_0__inst_r_sum1_9__19__q ),
	.datac(!Xd_0__inst_r_sum1_9__18__q ),
	.datad(!Xd_0__inst_r_sum1_8__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__19__q ),
	.datab(!Xd_0__inst_r_sum1_7__19__q ),
	.datac(!Xd_0__inst_r_sum1_7__18__q ),
	.datad(!Xd_0__inst_r_sum1_6__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__19__q ),
	.datab(!Xd_0__inst_r_sum1_5__19__q ),
	.datac(!Xd_0__inst_r_sum1_5__18__q ),
	.datad(!Xd_0__inst_r_sum1_4__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__19__q ),
	.datab(!Xd_0__inst_r_sum1_3__19__q ),
	.datac(!Xd_0__inst_r_sum1_3__18__q ),
	.datad(!Xd_0__inst_r_sum1_2__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__19__q ),
	.datab(!Xd_0__inst_r_sum1_1__19__q ),
	.datac(!Xd_0__inst_r_sum1_1__18__q ),
	.datad(!Xd_0__inst_r_sum1_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__19__q ),
	.datab(!Xd_0__inst_r_sum1_15__19__q ),
	.datac(!Xd_0__inst_r_sum1_14__20__q ),
	.datad(!Xd_0__inst_r_sum1_15__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__19__q ),
	.datab(!Xd_0__inst_r_sum1_13__19__q ),
	.datac(!Xd_0__inst_r_sum1_12__20__q ),
	.datad(!Xd_0__inst_r_sum1_13__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__19__q ),
	.datab(!Xd_0__inst_r_sum1_11__19__q ),
	.datac(!Xd_0__inst_r_sum1_10__20__q ),
	.datad(!Xd_0__inst_r_sum1_11__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__19__q ),
	.datab(!Xd_0__inst_r_sum1_9__19__q ),
	.datac(!Xd_0__inst_r_sum1_8__20__q ),
	.datad(!Xd_0__inst_r_sum1_9__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__19__q ),
	.datab(!Xd_0__inst_r_sum1_7__19__q ),
	.datac(!Xd_0__inst_r_sum1_6__20__q ),
	.datad(!Xd_0__inst_r_sum1_7__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__19__q ),
	.datab(!Xd_0__inst_r_sum1_5__19__q ),
	.datac(!Xd_0__inst_r_sum1_4__20__q ),
	.datad(!Xd_0__inst_r_sum1_5__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__19__q ),
	.datab(!Xd_0__inst_r_sum1_3__19__q ),
	.datac(!Xd_0__inst_r_sum1_2__20__q ),
	.datad(!Xd_0__inst_r_sum1_3__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__19__q ),
	.datab(!Xd_0__inst_r_sum1_1__19__q ),
	.datac(!Xd_0__inst_r_sum1_0__20__q ),
	.datad(!Xd_0__inst_r_sum1_1__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__21__q ),
	.datab(!Xd_0__inst_r_sum1_15__21__q ),
	.datac(!Xd_0__inst_r_sum1_15__20__q ),
	.datad(!Xd_0__inst_r_sum1_14__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__21__q ),
	.datab(!Xd_0__inst_r_sum1_13__21__q ),
	.datac(!Xd_0__inst_r_sum1_13__20__q ),
	.datad(!Xd_0__inst_r_sum1_12__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__21__q ),
	.datab(!Xd_0__inst_r_sum1_11__21__q ),
	.datac(!Xd_0__inst_r_sum1_11__20__q ),
	.datad(!Xd_0__inst_r_sum1_10__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__21__q ),
	.datab(!Xd_0__inst_r_sum1_9__21__q ),
	.datac(!Xd_0__inst_r_sum1_9__20__q ),
	.datad(!Xd_0__inst_r_sum1_8__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__21__q ),
	.datab(!Xd_0__inst_r_sum1_7__21__q ),
	.datac(!Xd_0__inst_r_sum1_7__20__q ),
	.datad(!Xd_0__inst_r_sum1_6__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__21__q ),
	.datab(!Xd_0__inst_r_sum1_5__21__q ),
	.datac(!Xd_0__inst_r_sum1_5__20__q ),
	.datad(!Xd_0__inst_r_sum1_4__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__21__q ),
	.datab(!Xd_0__inst_r_sum1_3__21__q ),
	.datac(!Xd_0__inst_r_sum1_3__20__q ),
	.datad(!Xd_0__inst_r_sum1_2__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__21__q ),
	.datab(!Xd_0__inst_r_sum1_1__21__q ),
	.datac(!Xd_0__inst_r_sum1_1__20__q ),
	.datad(!Xd_0__inst_r_sum1_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__21__q ),
	.datab(!Xd_0__inst_r_sum1_15__21__q ),
	.datac(!Xd_0__inst_r_sum1_14__22__q ),
	.datad(!Xd_0__inst_r_sum1_15__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__21__q ),
	.datab(!Xd_0__inst_r_sum1_13__21__q ),
	.datac(!Xd_0__inst_r_sum1_12__22__q ),
	.datad(!Xd_0__inst_r_sum1_13__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__21__q ),
	.datab(!Xd_0__inst_r_sum1_11__21__q ),
	.datac(!Xd_0__inst_r_sum1_10__22__q ),
	.datad(!Xd_0__inst_r_sum1_11__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__21__q ),
	.datab(!Xd_0__inst_r_sum1_9__21__q ),
	.datac(!Xd_0__inst_r_sum1_8__22__q ),
	.datad(!Xd_0__inst_r_sum1_9__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__21__q ),
	.datab(!Xd_0__inst_r_sum1_7__21__q ),
	.datac(!Xd_0__inst_r_sum1_6__22__q ),
	.datad(!Xd_0__inst_r_sum1_7__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__21__q ),
	.datab(!Xd_0__inst_r_sum1_5__21__q ),
	.datac(!Xd_0__inst_r_sum1_4__22__q ),
	.datad(!Xd_0__inst_r_sum1_5__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__21__q ),
	.datab(!Xd_0__inst_r_sum1_3__21__q ),
	.datac(!Xd_0__inst_r_sum1_2__22__q ),
	.datad(!Xd_0__inst_r_sum1_3__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001101EE1),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__21__q ),
	.datab(!Xd_0__inst_r_sum1_1__21__q ),
	.datac(!Xd_0__inst_r_sum1_0__22__q ),
	.datad(!Xd_0__inst_r_sum1_1__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__23__q ),
	.datab(!Xd_0__inst_r_sum1_15__23__q ),
	.datac(!Xd_0__inst_r_sum1_15__22__q ),
	.datad(!Xd_0__inst_r_sum1_14__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__23__q ),
	.datab(!Xd_0__inst_r_sum1_13__23__q ),
	.datac(!Xd_0__inst_r_sum1_13__22__q ),
	.datad(!Xd_0__inst_r_sum1_12__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__23__q ),
	.datab(!Xd_0__inst_r_sum1_11__23__q ),
	.datac(!Xd_0__inst_r_sum1_11__22__q ),
	.datad(!Xd_0__inst_r_sum1_10__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__23__q ),
	.datab(!Xd_0__inst_r_sum1_9__23__q ),
	.datac(!Xd_0__inst_r_sum1_9__22__q ),
	.datad(!Xd_0__inst_r_sum1_8__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__23__q ),
	.datab(!Xd_0__inst_r_sum1_7__23__q ),
	.datac(!Xd_0__inst_r_sum1_7__22__q ),
	.datad(!Xd_0__inst_r_sum1_6__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__23__q ),
	.datab(!Xd_0__inst_r_sum1_5__23__q ),
	.datac(!Xd_0__inst_r_sum1_5__22__q ),
	.datad(!Xd_0__inst_r_sum1_4__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__23__q ),
	.datab(!Xd_0__inst_r_sum1_3__23__q ),
	.datac(!Xd_0__inst_r_sum1_3__22__q ),
	.datad(!Xd_0__inst_r_sum1_2__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__23__q ),
	.datab(!Xd_0__inst_r_sum1_1__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__22__q ),
	.datad(!Xd_0__inst_r_sum1_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_116_sumout ),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_14__23__q ),
	.datab(!Xd_0__inst_r_sum1_15__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_7__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_7__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_12__23__q ),
	.datab(!Xd_0__inst_r_sum1_13__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_6__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_6__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_10__23__q ),
	.datab(!Xd_0__inst_r_sum1_11__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_5__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_5__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_8__23__q ),
	.datab(!Xd_0__inst_r_sum1_9__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_4__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_4__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_6__23__q ),
	.datab(!Xd_0__inst_r_sum1_7__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_3__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_3__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_4__23__q ),
	.datab(!Xd_0__inst_r_sum1_5__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_2__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_2__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_2__23__q ),
	.datab(!Xd_0__inst_r_sum1_3__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_1__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_1__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000007777),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_r_sum1_0__23__q ),
	.datab(!Xd_0__inst_r_sum1_1__23__q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a2_0__adder2_inst_add_0_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a2_0__adder2_inst_add_0_121_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_7__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_7__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_6__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [12]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_6__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_85 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[304]),
	.datac(!Xd_0__inst_mult_25_229 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_219 ),
	.cout(Xd_0__inst_mult_25_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_35 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[364]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_35_sumout ),
	.cout(Xd_0__inst_mult_30_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_45 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[303]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_45_sumout ),
	.cout(Xd_0__inst_mult_25_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_219 ),
	.datab(!Xd_0__inst_mult_25_45_sumout ),
	.datac(!Xd_0__inst_mult_25_239 ),
	.datad(!Xd_0__inst_mult_25_234 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_224 ),
	.cout(Xd_0__inst_mult_25_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_5__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_5__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_4__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [8]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_4__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_94 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[292]),
	.datac(!Xd_0__inst_mult_24_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_264 ),
	.cout(Xd_0__inst_mult_24_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_50 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[291]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_50_sumout ),
	.cout(Xd_0__inst_mult_24_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_264 ),
	.datab(!Xd_0__inst_mult_24_50_sumout ),
	.datac(!Xd_0__inst_mult_24_304 ),
	.datad(!Xd_0__inst_mult_24_299 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_269 ),
	.cout(Xd_0__inst_mult_24_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_94 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[322]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_264 ),
	.cout(Xd_0__inst_mult_26_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_95 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_294 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_269 ),
	.cout(Xd_0__inst_mult_26_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_96 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[319]),
	.datac(!Xd_0__inst_mult_26_304 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_274 ),
	.cout(Xd_0__inst_mult_26_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_274 ),
	.datab(!Xd_0__inst_mult_26_269 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_279 ),
	.cout(Xd_0__inst_mult_26_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_3__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_3__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_2__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_2__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_85 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[328]),
	.datac(!Xd_0__inst_mult_27_229 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_219 ),
	.cout(Xd_0__inst_mult_27_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_50 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[327]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_50_sumout ),
	.cout(Xd_0__inst_mult_27_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_219 ),
	.datab(!Xd_0__inst_mult_27_50_sumout ),
	.datac(!Xd_0__inst_mult_27_239 ),
	.datad(!Xd_0__inst_mult_27_234 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_224 ),
	.cout(Xd_0__inst_mult_27_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_1__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_1__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000F0F0000),
	.shared_arith("off")
) Xd_0__inst_a2_0__adder2_inst_add_0_127 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_r_sign [0]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a2_0__adder2_inst_add_0_127_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_98 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[316]),
	.datac(!Xd_0__inst_mult_26_319 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_284 ),
	.cout(Xd_0__inst_mult_26_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_50 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[315]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_50_sumout ),
	.cout(Xd_0__inst_mult_26_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_284 ),
	.datab(!Xd_0__inst_mult_26_50_sumout ),
	.datac(!Xd_0__inst_mult_26_329 ),
	.datad(!Xd_0__inst_mult_26_324 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_289 ),
	.cout(Xd_0__inst_mult_26_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_96 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[298]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_274 ),
	.cout(Xd_0__inst_mult_24_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_97 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_279 ),
	.cout(Xd_0__inst_mult_24_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_98 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[295]),
	.datac(!Xd_0__inst_mult_24_324 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_284 ),
	.cout(Xd_0__inst_mult_24_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_284 ),
	.datab(!Xd_0__inst_mult_24_279 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_289 ),
	.cout(Xd_0__inst_mult_24_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_88 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[30]),
	.datac(!din_a[27]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_234 ),
	.cout(Xd_0__inst_mult_2_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [30]),
	.datab(!Xd_0__inst_sign [31]),
	.datac(!Xd_0__inst_product_31__0__q ),
	.datad(!Xd_0__inst_product_30__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [28]),
	.datab(!Xd_0__inst_sign [29]),
	.datac(!Xd_0__inst_product_29__0__q ),
	.datad(!Xd_0__inst_product_28__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_210 ),
	.datab(!Xd_0__inst_mult_21_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_205 ),
	.cout(Xd_0__inst_mult_21_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [26]),
	.datab(!Xd_0__inst_sign [27]),
	.datac(!Xd_0__inst_product_27__0__q ),
	.datad(!Xd_0__inst_product_26__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [24]),
	.datab(!Xd_0__inst_sign [25]),
	.datac(!Xd_0__inst_product_25__0__q ),
	.datad(!Xd_0__inst_product_24__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_210 ),
	.datab(!Xd_0__inst_mult_20_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_205 ),
	.cout(Xd_0__inst_mult_20_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_229 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_88 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[303]),
	.datac(!Xd_0__inst_mult_25_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_234 ),
	.cout(Xd_0__inst_mult_25_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_89 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_239 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_239 ),
	.datab(!Xd_0__inst_mult_25_234 ),
	.datac(!din_a[310]),
	.datad(!din_b[302]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_244 ),
	.cout(Xd_0__inst_mult_25_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [22]),
	.datab(!Xd_0__inst_sign [23]),
	.datac(!Xd_0__inst_product_23__0__q ),
	.datad(!Xd_0__inst_product_22__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [20]),
	.datab(!Xd_0__inst_sign [21]),
	.datac(!Xd_0__inst_product_21__0__q ),
	.datad(!Xd_0__inst_product_20__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_210 ),
	.datab(!Xd_0__inst_mult_23_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_205 ),
	.cout(Xd_0__inst_mult_23_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [18]),
	.datab(!Xd_0__inst_sign [19]),
	.datac(!Xd_0__inst_product_19__0__q ),
	.datad(!Xd_0__inst_product_18__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [16]),
	.datab(!Xd_0__inst_sign [17]),
	.datac(!Xd_0__inst_product_17__0__q ),
	.datad(!Xd_0__inst_product_16__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_210 ),
	.datab(!Xd_0__inst_mult_22_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_205 ),
	.cout(Xd_0__inst_mult_22_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_101 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[291]),
	.datac(!Xd_0__inst_mult_24_339 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_299 ),
	.cout(Xd_0__inst_mult_24_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_102 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_304 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_304 ),
	.datab(!Xd_0__inst_mult_24_299 ),
	.datac(!din_a[298]),
	.datad(!din_b[290]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_309 ),
	.cout(Xd_0__inst_mult_24_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_100 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[321]),
	.datac(!din_a[318]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_294 ),
	.cout(Xd_0__inst_mult_26_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_101 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_339 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_299 ),
	.cout(Xd_0__inst_mult_26_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_102 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_304 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_103 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[318]),
	.datac(!Xd_0__inst_mult_26_349 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_309 ),
	.cout(Xd_0__inst_mult_26_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_309 ),
	.datab(!Xd_0__inst_mult_26_299 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_314 ),
	.cout(Xd_0__inst_mult_26_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [14]),
	.datab(!Xd_0__inst_sign [15]),
	.datac(!Xd_0__inst_product_15__0__q ),
	.datad(!Xd_0__inst_product_14__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [12]),
	.datab(!Xd_0__inst_sign [13]),
	.datac(!Xd_0__inst_product_13__0__q ),
	.datad(!Xd_0__inst_product_12__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_210 ),
	.datab(!Xd_0__inst_mult_19_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_205 ),
	.cout(Xd_0__inst_mult_19_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [10]),
	.datab(!Xd_0__inst_sign [11]),
	.datac(!Xd_0__inst_product_11__0__q ),
	.datad(!Xd_0__inst_product_10__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [8]),
	.datab(!Xd_0__inst_sign [9]),
	.datac(!Xd_0__inst_product_9__0__q ),
	.datad(!Xd_0__inst_product_8__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_210 ),
	.datab(!Xd_0__inst_mult_17_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_205 ),
	.cout(Xd_0__inst_mult_17_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_87 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_229 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_88 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[327]),
	.datac(!Xd_0__inst_mult_27_249 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_234 ),
	.cout(Xd_0__inst_mult_27_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_89 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_239 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_239 ),
	.datab(!Xd_0__inst_mult_27_234 ),
	.datac(!din_a[334]),
	.datad(!din_b[326]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_244 ),
	.cout(Xd_0__inst_mult_27_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [6]),
	.datab(!Xd_0__inst_sign [7]),
	.datac(!Xd_0__inst_product_7__0__q ),
	.datad(!Xd_0__inst_product_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [4]),
	.datab(!Xd_0__inst_sign [5]),
	.datac(!Xd_0__inst_product_5__0__q ),
	.datad(!Xd_0__inst_product_4__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_210 ),
	.datab(!Xd_0__inst_mult_16_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_205 ),
	.cout(Xd_0__inst_mult_16_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [2]),
	.datab(!Xd_0__inst_sign [3]),
	.datac(!Xd_0__inst_product_3__0__q ),
	.datad(!Xd_0__inst_product_2__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000014286996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_1 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [0]),
	.datab(!Xd_0__inst_sign [1]),
	.datac(!Xd_0__inst_product_1__0__q ),
	.datad(!Xd_0__inst_product_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_122_cout ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_210 ),
	.datab(!Xd_0__inst_mult_29_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_205 ),
	.cout(Xd_0__inst_mult_29_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_105 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_319 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_106 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[315]),
	.datac(!Xd_0__inst_mult_26_364 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_324 ),
	.cout(Xd_0__inst_mult_26_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_26_107 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_329 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_108 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_329 ),
	.datab(!Xd_0__inst_mult_26_324 ),
	.datac(!din_a[322]),
	.datad(!din_b[314]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_334 ),
	.cout(Xd_0__inst_mult_26_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_104 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[297]),
	.datac(!din_a[294]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_314 ),
	.cout(Xd_0__inst_mult_24_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_105 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_359 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_319 ),
	.cout(Xd_0__inst_mult_24_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_24_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_107 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[294]),
	.datac(!Xd_0__inst_mult_24_369 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_329 ),
	.cout(Xd_0__inst_mult_24_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_108 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_329 ),
	.datab(!Xd_0__inst_mult_24_319 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_334 ),
	.cout(Xd_0__inst_mult_24_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_89 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[30]),
	.datac(!din_a[26]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_239 ),
	.cout(Xd_0__inst_mult_2_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__1__q ),
	.datad(!Xd_0__inst_product_28__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__1__q ),
	.datad(!Xd_0__inst_product_30__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__1__q ),
	.datad(!Xd_0__inst_product_24__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__1__q ),
	.datad(!Xd_0__inst_product_26__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__1__q ),
	.datad(!Xd_0__inst_product_20__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__1__q ),
	.datad(!Xd_0__inst_product_22__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__1__q ),
	.datad(!Xd_0__inst_product_16__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__1__q ),
	.datad(!Xd_0__inst_product_18__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__1__q ),
	.datad(!Xd_0__inst_product_12__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__1__q ),
	.datad(!Xd_0__inst_product_14__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__1__q ),
	.datad(!Xd_0__inst_product_8__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__1__q ),
	.datad(!Xd_0__inst_product_10__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__1__q ),
	.datad(!Xd_0__inst_product_4__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__1__q ),
	.datad(!Xd_0__inst_product_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__1__q ),
	.datad(!Xd_0__inst_product_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_6 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__1__q ),
	.datad(!Xd_0__inst_product_2__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__2__q ),
	.datad(!Xd_0__inst_product_28__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__2__q ),
	.datad(!Xd_0__inst_product_30__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__2__q ),
	.datad(!Xd_0__inst_product_24__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__2__q ),
	.datad(!Xd_0__inst_product_26__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__2__q ),
	.datad(!Xd_0__inst_product_20__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__2__q ),
	.datad(!Xd_0__inst_product_22__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__2__q ),
	.datad(!Xd_0__inst_product_16__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__2__q ),
	.datad(!Xd_0__inst_product_18__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__2__q ),
	.datad(!Xd_0__inst_product_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__2__q ),
	.datad(!Xd_0__inst_product_14__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__2__q ),
	.datad(!Xd_0__inst_product_8__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__2__q ),
	.datad(!Xd_0__inst_product_10__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__2__q ),
	.datad(!Xd_0__inst_product_4__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__2__q ),
	.datad(!Xd_0__inst_product_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__2__q ),
	.datad(!Xd_0__inst_product_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_11 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__2__q ),
	.datad(!Xd_0__inst_product_2__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__3__q ),
	.datad(!Xd_0__inst_product_28__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__3__q ),
	.datad(!Xd_0__inst_product_30__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__3__q ),
	.datad(!Xd_0__inst_product_24__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__3__q ),
	.datad(!Xd_0__inst_product_26__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__3__q ),
	.datad(!Xd_0__inst_product_20__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__3__q ),
	.datad(!Xd_0__inst_product_22__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__3__q ),
	.datad(!Xd_0__inst_product_16__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__3__q ),
	.datad(!Xd_0__inst_product_18__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__3__q ),
	.datad(!Xd_0__inst_product_12__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__3__q ),
	.datad(!Xd_0__inst_product_14__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__3__q ),
	.datad(!Xd_0__inst_product_8__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__3__q ),
	.datad(!Xd_0__inst_product_10__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__3__q ),
	.datad(!Xd_0__inst_product_4__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__3__q ),
	.datad(!Xd_0__inst_product_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__3__q ),
	.datad(!Xd_0__inst_product_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_16 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__3__q ),
	.datad(!Xd_0__inst_product_2__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__4__q ),
	.datad(!Xd_0__inst_product_28__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__4__q ),
	.datad(!Xd_0__inst_product_30__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__4__q ),
	.datad(!Xd_0__inst_product_24__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__4__q ),
	.datad(!Xd_0__inst_product_26__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__4__q ),
	.datad(!Xd_0__inst_product_20__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__4__q ),
	.datad(!Xd_0__inst_product_22__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__4__q ),
	.datad(!Xd_0__inst_product_16__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__4__q ),
	.datad(!Xd_0__inst_product_18__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__4__q ),
	.datad(!Xd_0__inst_product_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__4__q ),
	.datad(!Xd_0__inst_product_14__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__4__q ),
	.datad(!Xd_0__inst_product_8__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__4__q ),
	.datad(!Xd_0__inst_product_10__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__4__q ),
	.datad(!Xd_0__inst_product_4__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__4__q ),
	.datad(!Xd_0__inst_product_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__4__q ),
	.datad(!Xd_0__inst_product_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_21 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__4__q ),
	.datad(!Xd_0__inst_product_2__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__5__q ),
	.datad(!Xd_0__inst_product_28__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__5__q ),
	.datad(!Xd_0__inst_product_30__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__5__q ),
	.datad(!Xd_0__inst_product_24__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__5__q ),
	.datad(!Xd_0__inst_product_26__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__5__q ),
	.datad(!Xd_0__inst_product_20__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__5__q ),
	.datad(!Xd_0__inst_product_22__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__5__q ),
	.datad(!Xd_0__inst_product_16__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__5__q ),
	.datad(!Xd_0__inst_product_18__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__5__q ),
	.datad(!Xd_0__inst_product_12__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__5__q ),
	.datad(!Xd_0__inst_product_14__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__5__q ),
	.datad(!Xd_0__inst_product_8__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__5__q ),
	.datad(!Xd_0__inst_product_10__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__5__q ),
	.datad(!Xd_0__inst_product_4__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__5__q ),
	.datad(!Xd_0__inst_product_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__5__q ),
	.datad(!Xd_0__inst_product_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_26 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__5__q ),
	.datad(!Xd_0__inst_product_2__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__6__q ),
	.datad(!Xd_0__inst_product_28__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__6__q ),
	.datad(!Xd_0__inst_product_30__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__6__q ),
	.datad(!Xd_0__inst_product_24__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__6__q ),
	.datad(!Xd_0__inst_product_26__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__6__q ),
	.datad(!Xd_0__inst_product_20__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__6__q ),
	.datad(!Xd_0__inst_product_22__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__6__q ),
	.datad(!Xd_0__inst_product_16__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__6__q ),
	.datad(!Xd_0__inst_product_18__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__6__q ),
	.datad(!Xd_0__inst_product_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__6__q ),
	.datad(!Xd_0__inst_product_14__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__6__q ),
	.datad(!Xd_0__inst_product_8__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__6__q ),
	.datad(!Xd_0__inst_product_10__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__6__q ),
	.datad(!Xd_0__inst_product_4__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__6__q ),
	.datad(!Xd_0__inst_product_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__6__q ),
	.datad(!Xd_0__inst_product_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_31 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__6__q ),
	.datad(!Xd_0__inst_product_2__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__7__q ),
	.datad(!Xd_0__inst_product_28__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__7__q ),
	.datad(!Xd_0__inst_product_30__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__7__q ),
	.datad(!Xd_0__inst_product_24__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__7__q ),
	.datad(!Xd_0__inst_product_26__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__7__q ),
	.datad(!Xd_0__inst_product_20__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__7__q ),
	.datad(!Xd_0__inst_product_22__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__7__q ),
	.datad(!Xd_0__inst_product_16__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__7__q ),
	.datad(!Xd_0__inst_product_18__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__7__q ),
	.datad(!Xd_0__inst_product_12__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__7__q ),
	.datad(!Xd_0__inst_product_14__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__7__q ),
	.datad(!Xd_0__inst_product_8__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__7__q ),
	.datad(!Xd_0__inst_product_10__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__7__q ),
	.datad(!Xd_0__inst_product_4__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__7__q ),
	.datad(!Xd_0__inst_product_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__7__q ),
	.datad(!Xd_0__inst_product_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_36 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__7__q ),
	.datad(!Xd_0__inst_product_2__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__8__q ),
	.datad(!Xd_0__inst_product_28__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__8__q ),
	.datad(!Xd_0__inst_product_30__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__8__q ),
	.datad(!Xd_0__inst_product_24__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__8__q ),
	.datad(!Xd_0__inst_product_26__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__8__q ),
	.datad(!Xd_0__inst_product_20__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__8__q ),
	.datad(!Xd_0__inst_product_22__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__8__q ),
	.datad(!Xd_0__inst_product_16__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__8__q ),
	.datad(!Xd_0__inst_product_18__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__8__q ),
	.datad(!Xd_0__inst_product_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__8__q ),
	.datad(!Xd_0__inst_product_14__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__8__q ),
	.datad(!Xd_0__inst_product_8__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__8__q ),
	.datad(!Xd_0__inst_product_10__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__8__q ),
	.datad(!Xd_0__inst_product_4__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__8__q ),
	.datad(!Xd_0__inst_product_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__8__q ),
	.datad(!Xd_0__inst_product_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_41 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__8__q ),
	.datad(!Xd_0__inst_product_2__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__9__q ),
	.datad(!Xd_0__inst_product_28__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__9__q ),
	.datad(!Xd_0__inst_product_30__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__9__q ),
	.datad(!Xd_0__inst_product_24__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__9__q ),
	.datad(!Xd_0__inst_product_26__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__9__q ),
	.datad(!Xd_0__inst_product_20__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__9__q ),
	.datad(!Xd_0__inst_product_22__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__9__q ),
	.datad(!Xd_0__inst_product_16__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__9__q ),
	.datad(!Xd_0__inst_product_18__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__9__q ),
	.datad(!Xd_0__inst_product_12__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__9__q ),
	.datad(!Xd_0__inst_product_14__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__9__q ),
	.datad(!Xd_0__inst_product_8__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__9__q ),
	.datad(!Xd_0__inst_product_10__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__9__q ),
	.datad(!Xd_0__inst_product_4__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__9__q ),
	.datad(!Xd_0__inst_product_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__9__q ),
	.datad(!Xd_0__inst_product_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_46 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__9__q ),
	.datad(!Xd_0__inst_product_2__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__10__q ),
	.datad(!Xd_0__inst_product_28__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__10__q ),
	.datad(!Xd_0__inst_product_30__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__10__q ),
	.datad(!Xd_0__inst_product_24__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__10__q ),
	.datad(!Xd_0__inst_product_26__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__10__q ),
	.datad(!Xd_0__inst_product_20__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__10__q ),
	.datad(!Xd_0__inst_product_22__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__10__q ),
	.datad(!Xd_0__inst_product_16__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__10__q ),
	.datad(!Xd_0__inst_product_18__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__10__q ),
	.datad(!Xd_0__inst_product_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__10__q ),
	.datad(!Xd_0__inst_product_14__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__10__q ),
	.datad(!Xd_0__inst_product_8__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__10__q ),
	.datad(!Xd_0__inst_product_10__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__10__q ),
	.datad(!Xd_0__inst_product_4__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__10__q ),
	.datad(!Xd_0__inst_product_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__10__q ),
	.datad(!Xd_0__inst_product_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_51 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__10__q ),
	.datad(!Xd_0__inst_product_2__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__11__q ),
	.datad(!Xd_0__inst_product_28__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__11__q ),
	.datad(!Xd_0__inst_product_30__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__11__q ),
	.datad(!Xd_0__inst_product_24__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__11__q ),
	.datad(!Xd_0__inst_product_26__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__11__q ),
	.datad(!Xd_0__inst_product_20__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__11__q ),
	.datad(!Xd_0__inst_product_22__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__11__q ),
	.datad(!Xd_0__inst_product_16__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__11__q ),
	.datad(!Xd_0__inst_product_18__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__11__q ),
	.datad(!Xd_0__inst_product_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__11__q ),
	.datad(!Xd_0__inst_product_14__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__11__q ),
	.datad(!Xd_0__inst_product_8__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__11__q ),
	.datad(!Xd_0__inst_product_10__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__11__q ),
	.datad(!Xd_0__inst_product_4__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__11__q ),
	.datad(!Xd_0__inst_product_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__11__q ),
	.datad(!Xd_0__inst_product_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_56 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__11__q ),
	.datad(!Xd_0__inst_product_2__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__12__q ),
	.datad(!Xd_0__inst_product_28__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__12__q ),
	.datad(!Xd_0__inst_product_30__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__12__q ),
	.datad(!Xd_0__inst_product_24__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__12__q ),
	.datad(!Xd_0__inst_product_26__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__12__q ),
	.datad(!Xd_0__inst_product_20__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__12__q ),
	.datad(!Xd_0__inst_product_22__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__12__q ),
	.datad(!Xd_0__inst_product_16__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__12__q ),
	.datad(!Xd_0__inst_product_18__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__12__q ),
	.datad(!Xd_0__inst_product_12__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__12__q ),
	.datad(!Xd_0__inst_product_14__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__12__q ),
	.datad(!Xd_0__inst_product_8__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__12__q ),
	.datad(!Xd_0__inst_product_10__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__12__q ),
	.datad(!Xd_0__inst_product_4__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__12__q ),
	.datad(!Xd_0__inst_product_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__12__q ),
	.datad(!Xd_0__inst_product_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_61 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__12__q ),
	.datad(!Xd_0__inst_product_2__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__13__q ),
	.datad(!Xd_0__inst_product_28__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__13__q ),
	.datad(!Xd_0__inst_product_30__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__13__q ),
	.datad(!Xd_0__inst_product_24__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__13__q ),
	.datad(!Xd_0__inst_product_26__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__13__q ),
	.datad(!Xd_0__inst_product_20__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__13__q ),
	.datad(!Xd_0__inst_product_22__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__13__q ),
	.datad(!Xd_0__inst_product_16__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__13__q ),
	.datad(!Xd_0__inst_product_18__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__13__q ),
	.datad(!Xd_0__inst_product_12__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__13__q ),
	.datad(!Xd_0__inst_product_14__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__13__q ),
	.datad(!Xd_0__inst_product_8__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__13__q ),
	.datad(!Xd_0__inst_product_10__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__13__q ),
	.datad(!Xd_0__inst_product_4__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__13__q ),
	.datad(!Xd_0__inst_product_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__13__q ),
	.datad(!Xd_0__inst_product_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_66 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__13__q ),
	.datad(!Xd_0__inst_product_2__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__14__q ),
	.datad(!Xd_0__inst_product_28__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__14__q ),
	.datad(!Xd_0__inst_product_30__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__14__q ),
	.datad(!Xd_0__inst_product_24__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__14__q ),
	.datad(!Xd_0__inst_product_26__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__14__q ),
	.datad(!Xd_0__inst_product_20__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__14__q ),
	.datad(!Xd_0__inst_product_22__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__14__q ),
	.datad(!Xd_0__inst_product_16__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__14__q ),
	.datad(!Xd_0__inst_product_18__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__14__q ),
	.datad(!Xd_0__inst_product_12__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__14__q ),
	.datad(!Xd_0__inst_product_14__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__14__q ),
	.datad(!Xd_0__inst_product_8__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__14__q ),
	.datad(!Xd_0__inst_product_10__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__14__q ),
	.datad(!Xd_0__inst_product_4__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__14__q ),
	.datad(!Xd_0__inst_product_6__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__14__q ),
	.datad(!Xd_0__inst_product_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_71 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__14__q ),
	.datad(!Xd_0__inst_product_2__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__15__q ),
	.datad(!Xd_0__inst_product_28__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__15__q ),
	.datad(!Xd_0__inst_product_30__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__15__q ),
	.datad(!Xd_0__inst_product_24__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__15__q ),
	.datad(!Xd_0__inst_product_26__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__15__q ),
	.datad(!Xd_0__inst_product_20__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__15__q ),
	.datad(!Xd_0__inst_product_22__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__15__q ),
	.datad(!Xd_0__inst_product_16__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__15__q ),
	.datad(!Xd_0__inst_product_18__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__15__q ),
	.datad(!Xd_0__inst_product_12__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__15__q ),
	.datad(!Xd_0__inst_product_14__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__15__q ),
	.datad(!Xd_0__inst_product_8__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__15__q ),
	.datad(!Xd_0__inst_product_10__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__15__q ),
	.datad(!Xd_0__inst_product_4__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__15__q ),
	.datad(!Xd_0__inst_product_6__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__15__q ),
	.datad(!Xd_0__inst_product_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_76 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__15__q ),
	.datad(!Xd_0__inst_product_2__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__16__q ),
	.datad(!Xd_0__inst_product_28__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__16__q ),
	.datad(!Xd_0__inst_product_30__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__16__q ),
	.datad(!Xd_0__inst_product_24__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__16__q ),
	.datad(!Xd_0__inst_product_26__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__16__q ),
	.datad(!Xd_0__inst_product_20__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__16__q ),
	.datad(!Xd_0__inst_product_22__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__16__q ),
	.datad(!Xd_0__inst_product_16__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__16__q ),
	.datad(!Xd_0__inst_product_18__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__16__q ),
	.datad(!Xd_0__inst_product_12__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__16__q ),
	.datad(!Xd_0__inst_product_14__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__16__q ),
	.datad(!Xd_0__inst_product_8__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__16__q ),
	.datad(!Xd_0__inst_product_10__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__16__q ),
	.datad(!Xd_0__inst_product_4__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__16__q ),
	.datad(!Xd_0__inst_product_6__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__16__q ),
	.datad(!Xd_0__inst_product_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_81 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__16__q ),
	.datad(!Xd_0__inst_product_2__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__17__q ),
	.datad(!Xd_0__inst_product_28__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__17__q ),
	.datad(!Xd_0__inst_product_30__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__17__q ),
	.datad(!Xd_0__inst_product_24__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__17__q ),
	.datad(!Xd_0__inst_product_26__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__17__q ),
	.datad(!Xd_0__inst_product_20__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__17__q ),
	.datad(!Xd_0__inst_product_22__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__17__q ),
	.datad(!Xd_0__inst_product_16__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__17__q ),
	.datad(!Xd_0__inst_product_18__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__17__q ),
	.datad(!Xd_0__inst_product_12__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__17__q ),
	.datad(!Xd_0__inst_product_14__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__17__q ),
	.datad(!Xd_0__inst_product_8__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__17__q ),
	.datad(!Xd_0__inst_product_10__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__17__q ),
	.datad(!Xd_0__inst_product_4__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__17__q ),
	.datad(!Xd_0__inst_product_6__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__17__q ),
	.datad(!Xd_0__inst_product_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__17__q ),
	.datad(!Xd_0__inst_product_2__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_86_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__18__q ),
	.datad(!Xd_0__inst_product_28__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__18__q ),
	.datad(!Xd_0__inst_product_30__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__18__q ),
	.datad(!Xd_0__inst_product_24__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__18__q ),
	.datad(!Xd_0__inst_product_26__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__18__q ),
	.datad(!Xd_0__inst_product_20__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__18__q ),
	.datad(!Xd_0__inst_product_22__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__18__q ),
	.datad(!Xd_0__inst_product_16__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__18__q ),
	.datad(!Xd_0__inst_product_18__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__18__q ),
	.datad(!Xd_0__inst_product_12__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__18__q ),
	.datad(!Xd_0__inst_product_14__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__18__q ),
	.datad(!Xd_0__inst_product_8__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__18__q ),
	.datad(!Xd_0__inst_product_10__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__18__q ),
	.datad(!Xd_0__inst_product_4__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__18__q ),
	.datad(!Xd_0__inst_product_6__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__18__q ),
	.datad(!Xd_0__inst_product_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__18__q ),
	.datad(!Xd_0__inst_product_2__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_91_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__19__q ),
	.datad(!Xd_0__inst_product_28__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__19__q ),
	.datad(!Xd_0__inst_product_30__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__19__q ),
	.datad(!Xd_0__inst_product_24__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__19__q ),
	.datad(!Xd_0__inst_product_26__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__19__q ),
	.datad(!Xd_0__inst_product_20__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__19__q ),
	.datad(!Xd_0__inst_product_22__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__19__q ),
	.datad(!Xd_0__inst_product_16__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__19__q ),
	.datad(!Xd_0__inst_product_18__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__19__q ),
	.datad(!Xd_0__inst_product_12__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__19__q ),
	.datad(!Xd_0__inst_product_14__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__19__q ),
	.datad(!Xd_0__inst_product_8__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__19__q ),
	.datad(!Xd_0__inst_product_10__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__19__q ),
	.datad(!Xd_0__inst_product_4__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__19__q ),
	.datad(!Xd_0__inst_product_6__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__19__q ),
	.datad(!Xd_0__inst_product_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__19__q ),
	.datad(!Xd_0__inst_product_2__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_96_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__20__q ),
	.datad(!Xd_0__inst_product_28__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__20__q ),
	.datad(!Xd_0__inst_product_30__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__20__q ),
	.datad(!Xd_0__inst_product_24__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__20__q ),
	.datad(!Xd_0__inst_product_26__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__20__q ),
	.datad(!Xd_0__inst_product_20__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__20__q ),
	.datad(!Xd_0__inst_product_22__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__20__q ),
	.datad(!Xd_0__inst_product_16__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__20__q ),
	.datad(!Xd_0__inst_product_18__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__20__q ),
	.datad(!Xd_0__inst_product_12__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__20__q ),
	.datad(!Xd_0__inst_product_14__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__20__q ),
	.datad(!Xd_0__inst_product_8__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__20__q ),
	.datad(!Xd_0__inst_product_10__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__20__q ),
	.datad(!Xd_0__inst_product_4__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__20__q ),
	.datad(!Xd_0__inst_product_6__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__20__q ),
	.datad(!Xd_0__inst_product_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__20__q ),
	.datad(!Xd_0__inst_product_2__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_101_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(!Xd_0__inst_product_29__21__q ),
	.datad(!Xd_0__inst_product_28__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(!Xd_0__inst_product_31__21__q ),
	.datad(!Xd_0__inst_product_30__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(!Xd_0__inst_product_25__21__q ),
	.datad(!Xd_0__inst_product_24__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(!Xd_0__inst_product_27__21__q ),
	.datad(!Xd_0__inst_product_26__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(!Xd_0__inst_product_21__21__q ),
	.datad(!Xd_0__inst_product_20__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(!Xd_0__inst_product_23__21__q ),
	.datad(!Xd_0__inst_product_22__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(!Xd_0__inst_product_17__21__q ),
	.datad(!Xd_0__inst_product_16__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(!Xd_0__inst_product_19__21__q ),
	.datad(!Xd_0__inst_product_18__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(!Xd_0__inst_product_13__21__q ),
	.datad(!Xd_0__inst_product_12__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(!Xd_0__inst_product_15__21__q ),
	.datad(!Xd_0__inst_product_14__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(!Xd_0__inst_product_9__21__q ),
	.datad(!Xd_0__inst_product_8__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(!Xd_0__inst_product_11__21__q ),
	.datad(!Xd_0__inst_product_10__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(!Xd_0__inst_product_5__21__q ),
	.datad(!Xd_0__inst_product_4__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(!Xd_0__inst_product_7__21__q ),
	.datad(!Xd_0__inst_product_6__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(!Xd_0__inst_product_1__21__q ),
	.datad(!Xd_0__inst_product_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000012486996),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_106 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(!Xd_0__inst_product_3__21__q ),
	.datad(!Xd_0__inst_product_2__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_106_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [29]),
	.datab(!Xd_0__inst_sign [28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [31]),
	.datab(!Xd_0__inst_sign [30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [25]),
	.datab(!Xd_0__inst_sign [24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [27]),
	.datab(!Xd_0__inst_sign [26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [21]),
	.datab(!Xd_0__inst_sign [20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [23]),
	.datab(!Xd_0__inst_sign [22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [17]),
	.datab(!Xd_0__inst_sign [16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [19]),
	.datab(!Xd_0__inst_sign [18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [13]),
	.datab(!Xd_0__inst_sign [12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [15]),
	.datab(!Xd_0__inst_sign [14]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [9]),
	.datab(!Xd_0__inst_sign [8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [11]),
	.datab(!Xd_0__inst_sign [10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [5]),
	.datab(!Xd_0__inst_sign [4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [7]),
	.datab(!Xd_0__inst_sign [6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [1]),
	.datab(!Xd_0__inst_sign [0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_111 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [3]),
	.datab(!Xd_0__inst_sign [2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_111_sumout ),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [29]),
	.datad(!Xd_0__inst_sign [28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [31]),
	.datad(!Xd_0__inst_sign [30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [25]),
	.datad(!Xd_0__inst_sign [24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [27]),
	.datad(!Xd_0__inst_sign [26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [21]),
	.datad(!Xd_0__inst_sign [20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [23]),
	.datad(!Xd_0__inst_sign [22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [17]),
	.datad(!Xd_0__inst_sign [16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [19]),
	.datad(!Xd_0__inst_sign [18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [13]),
	.datad(!Xd_0__inst_sign [12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [15]),
	.datad(!Xd_0__inst_sign [14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [9]),
	.datad(!Xd_0__inst_sign [8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [11]),
	.datad(!Xd_0__inst_sign [10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [5]),
	.datad(!Xd_0__inst_sign [4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [7]),
	.datad(!Xd_0__inst_sign [6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [1]),
	.datad(!Xd_0__inst_sign [0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_116 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [3]),
	.datad(!Xd_0__inst_sign [2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_add_0_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_add_0_116_sumout ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_15__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [30]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_15__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_14__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [28]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_14__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_35 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[256]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_35_sumout ),
	.cout(Xd_0__inst_mult_21_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_210 ),
	.datab(!Xd_0__inst_mult_21_35_sumout ),
	.datac(!Xd_0__inst_mult_21_219 ),
	.datad(!Xd_0__inst_mult_21_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_214 ),
	.cout(Xd_0__inst_mult_21_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_13__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [26]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_13__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_12__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [24]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_12__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_35 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[244]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_35_sumout ),
	.cout(Xd_0__inst_mult_20_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_210 ),
	.datab(!Xd_0__inst_mult_20_35_sumout ),
	.datac(!Xd_0__inst_mult_20_219 ),
	.datad(!Xd_0__inst_mult_20_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_214 ),
	.cout(Xd_0__inst_mult_20_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_91 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[304]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_249 ),
	.cout(Xd_0__inst_mult_25_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_92 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_254 ),
	.cout(Xd_0__inst_mult_25_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_93 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[301]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_259 ),
	.cout(Xd_0__inst_mult_25_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_259 ),
	.datab(!Xd_0__inst_mult_25_254 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_264 ),
	.cout(Xd_0__inst_mult_25_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_11__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [22]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_11__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_10__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [20]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_10__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_35 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[280]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_35_sumout ),
	.cout(Xd_0__inst_mult_23_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_210 ),
	.datab(!Xd_0__inst_mult_23_35_sumout ),
	.datac(!Xd_0__inst_mult_23_219 ),
	.datad(!Xd_0__inst_mult_23_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_214 ),
	.cout(Xd_0__inst_mult_23_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_9__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [18]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_9__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_8__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [16]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_8__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_35 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[268]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_35_sumout ),
	.cout(Xd_0__inst_mult_22_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_210 ),
	.datab(!Xd_0__inst_mult_22_35_sumout ),
	.datac(!Xd_0__inst_mult_22_219 ),
	.datad(!Xd_0__inst_mult_22_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_214 ),
	.cout(Xd_0__inst_mult_22_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_109 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[292]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_339 ),
	.cout(Xd_0__inst_mult_24_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_110 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_344 ),
	.cout(Xd_0__inst_mult_24_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_111 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[289]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_349 ),
	.cout(Xd_0__inst_mult_24_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_112 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_349 ),
	.datab(!Xd_0__inst_mult_24_344 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_354 ),
	.cout(Xd_0__inst_mult_24_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_109 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[321]),
	.datac(!din_a[317]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_339 ),
	.cout(Xd_0__inst_mult_26_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_110 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_344 ),
	.cout(Xd_0__inst_mult_26_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_111 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[319]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_349 ),
	.cout(Xd_0__inst_mult_26_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_112 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_394 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_354 ),
	.cout(Xd_0__inst_mult_26_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_354 ),
	.datab(!Xd_0__inst_mult_26_344 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_359 ),
	.cout(Xd_0__inst_mult_26_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_7__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [14]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_7__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_6__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [12]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_6__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_35 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[232]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_35_sumout ),
	.cout(Xd_0__inst_mult_19_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_210 ),
	.datab(!Xd_0__inst_mult_19_35_sumout ),
	.datac(!Xd_0__inst_mult_19_219 ),
	.datad(!Xd_0__inst_mult_19_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_214 ),
	.cout(Xd_0__inst_mult_19_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_5__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [10]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_5__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_4__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [8]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_4__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_35 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[208]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_35_sumout ),
	.cout(Xd_0__inst_mult_17_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_210 ),
	.datab(!Xd_0__inst_mult_17_35_sumout ),
	.datac(!Xd_0__inst_mult_17_219 ),
	.datad(!Xd_0__inst_mult_17_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_214 ),
	.cout(Xd_0__inst_mult_17_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_91 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[328]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_249 ),
	.cout(Xd_0__inst_mult_27_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_92 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_269 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_254 ),
	.cout(Xd_0__inst_mult_27_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_93 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[325]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_259 ),
	.cout(Xd_0__inst_mult_27_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_259 ),
	.datab(!Xd_0__inst_mult_27_254 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_264 ),
	.cout(Xd_0__inst_mult_27_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_3__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [6]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_3__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_2__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [4]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_250 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_2__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_35 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[196]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_35_sumout ),
	.cout(Xd_0__inst_mult_16_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_210 ),
	.datab(!Xd_0__inst_mult_16_35_sumout ),
	.datac(!Xd_0__inst_mult_16_219 ),
	.datad(!Xd_0__inst_mult_16_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_214 ),
	.cout(Xd_0__inst_mult_16_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_1__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [2]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_1__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000055550000),
	.shared_arith("off")
) Xd_0__inst_a1_0__adder1_inst_add_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_sign [0]),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_206 ),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_a1_0__adder1_inst_add_0_122_cout ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_210 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_35 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[352]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_35_sumout ),
	.cout(Xd_0__inst_mult_29_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_210 ),
	.datab(!Xd_0__inst_mult_29_35_sumout ),
	.datac(!Xd_0__inst_mult_29_219 ),
	.datad(!Xd_0__inst_mult_29_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_214 ),
	.cout(Xd_0__inst_mult_29_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_114 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[316]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_364 ),
	.cout(Xd_0__inst_mult_26_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_115 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_409 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_369 ),
	.cout(Xd_0__inst_mult_26_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_116 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[313]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_374 ),
	.cout(Xd_0__inst_mult_26_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_374 ),
	.datab(!Xd_0__inst_mult_26_369 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_379 ),
	.cout(Xd_0__inst_mult_26_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_113 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[297]),
	.datac(!din_a[293]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_359 ),
	.cout(Xd_0__inst_mult_24_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_114 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_404 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_364 ),
	.cout(Xd_0__inst_mult_24_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_115 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[295]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_369 ),
	.cout(Xd_0__inst_mult_24_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_116 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_414 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_374 ),
	.cout(Xd_0__inst_mult_24_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_374 ),
	.datab(!Xd_0__inst_mult_24_364 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_379 ),
	.cout(Xd_0__inst_mult_24_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_90 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[30]),
	.datac(!din_a[25]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_244 ),
	.cout(Xd_0__inst_mult_2_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_294 ),
	.datab(!Xd_0__inst_mult_9_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_205 ),
	.cout(Xd_0__inst_mult_9_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_294 ),
	.datab(!Xd_0__inst_mult_8_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_205 ),
	.cout(Xd_0__inst_mult_8_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_1 (
// Equation(s):

	.dataa(!din_a[383]),
	.datab(!din_b[383]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_7 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_1_sumout ),
	.cout(Xd_0__inst_i29_2 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_85 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[256]),
	.datac(!Xd_0__inst_mult_21_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_219 ),
	.cout(Xd_0__inst_mult_21_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_35 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_35_sumout ),
	.cout(Xd_0__inst_mult_13_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_40 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[255]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_40_sumout ),
	.cout(Xd_0__inst_mult_21_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_219 ),
	.datab(!Xd_0__inst_mult_21_40_sumout ),
	.datac(!Xd_0__inst_mult_21_324 ),
	.datad(!Xd_0__inst_mult_21_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_224 ),
	.cout(Xd_0__inst_mult_21_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_294 ),
	.datab(!Xd_0__inst_mult_11_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_205 ),
	.cout(Xd_0__inst_mult_11_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_294 ),
	.datab(!Xd_0__inst_mult_10_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_205 ),
	.cout(Xd_0__inst_mult_10_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_6 (
// Equation(s):

	.dataa(!din_a[335]),
	.datab(!din_b[335]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_12 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_6_sumout ),
	.cout(Xd_0__inst_i29_7 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_85 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[244]),
	.datac(!Xd_0__inst_mult_20_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_219 ),
	.cout(Xd_0__inst_mult_20_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_40 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[249]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_40_sumout ),
	.cout(Xd_0__inst_mult_20_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_45 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[243]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_45_sumout ),
	.cout(Xd_0__inst_mult_20_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_219 ),
	.datab(!Xd_0__inst_mult_20_45_sumout ),
	.datac(!Xd_0__inst_mult_20_324 ),
	.datad(!Xd_0__inst_mult_20_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_224 ),
	.cout(Xd_0__inst_mult_20_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_95 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[303]),
	.datac(!din_a[307]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_269 ),
	.cout(Xd_0__inst_mult_25_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_96 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_374 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_274 ),
	.cout(Xd_0__inst_mult_25_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_97 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[301]),
	.datac(!din_a[310]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_279 ),
	.cout(Xd_0__inst_mult_25_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_279 ),
	.datab(!Xd_0__inst_mult_25_274 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_284 ),
	.cout(Xd_0__inst_mult_25_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_294 ),
	.datab(!Xd_0__inst_mult_3_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_205 ),
	.cout(Xd_0__inst_mult_3_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_294 ),
	.datab(!Xd_0__inst_mult_0_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_205 ),
	.cout(Xd_0__inst_mult_0_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_11 (
// Equation(s):

	.dataa(!din_a[287]),
	.datab(!din_b[287]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_17 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_11_sumout ),
	.cout(Xd_0__inst_i29_12 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_85 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[280]),
	.datac(!Xd_0__inst_mult_23_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_219 ),
	.cout(Xd_0__inst_mult_23_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_40 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[279]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_40_sumout ),
	.cout(Xd_0__inst_mult_23_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_219 ),
	.datab(!Xd_0__inst_mult_23_40_sumout ),
	.datac(!Xd_0__inst_mult_23_324 ),
	.datad(!Xd_0__inst_mult_23_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_224 ),
	.cout(Xd_0__inst_mult_23_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_294 ),
	.datab(!Xd_0__inst_mult_6_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_205 ),
	.cout(Xd_0__inst_mult_6_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_294 ),
	.datab(!Xd_0__inst_mult_1_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_205 ),
	.cout(Xd_0__inst_mult_1_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_16 (
// Equation(s):

	.dataa(!din_a[239]),
	.datab(!din_b[239]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_22 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_16_sumout ),
	.cout(Xd_0__inst_i29_17 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_85 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[268]),
	.datac(!Xd_0__inst_mult_22_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_219 ),
	.cout(Xd_0__inst_mult_22_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_40 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[267]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_40_sumout ),
	.cout(Xd_0__inst_mult_22_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_219 ),
	.datab(!Xd_0__inst_mult_22_40_sumout ),
	.datac(!Xd_0__inst_mult_22_324 ),
	.datad(!Xd_0__inst_mult_22_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_224 ),
	.cout(Xd_0__inst_mult_22_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_118 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[291]),
	.datac(!din_a[295]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_384 ),
	.cout(Xd_0__inst_mult_24_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_119 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_389 ),
	.cout(Xd_0__inst_mult_24_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_120 (
// Equation(s):

	.dataa(!din_a[297]),
	.datab(!din_b[289]),
	.datac(!din_a[298]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_394 ),
	.cout(Xd_0__inst_mult_24_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_394 ),
	.datab(!Xd_0__inst_mult_24_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_399 ),
	.cout(Xd_0__inst_mult_24_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_118 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[321]),
	.datac(!din_a[316]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_384 ),
	.cout(Xd_0__inst_mult_26_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_119 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_389 ),
	.cout(Xd_0__inst_mult_26_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_120 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[318]),
	.datac(!din_a[319]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_394 ),
	.cout(Xd_0__inst_mult_26_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_121 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_399 ),
	.cout(Xd_0__inst_mult_26_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_399 ),
	.datab(!Xd_0__inst_mult_26_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_404 ),
	.cout(Xd_0__inst_mult_26_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_294 ),
	.datab(!Xd_0__inst_mult_7_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_205 ),
	.cout(Xd_0__inst_mult_7_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_294 ),
	.datab(!Xd_0__inst_mult_4_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_205 ),
	.cout(Xd_0__inst_mult_4_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_21 (
// Equation(s):

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_27 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_21_sumout ),
	.cout(Xd_0__inst_i29_22 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_85 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[232]),
	.datac(!Xd_0__inst_mult_19_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_219 ),
	.cout(Xd_0__inst_mult_19_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_40 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[231]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_40_sumout ),
	.cout(Xd_0__inst_mult_19_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_219 ),
	.datab(!Xd_0__inst_mult_19_40_sumout ),
	.datac(!Xd_0__inst_mult_19_324 ),
	.datad(!Xd_0__inst_mult_19_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_224 ),
	.cout(Xd_0__inst_mult_19_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_294 ),
	.datab(!Xd_0__inst_mult_30_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_205 ),
	.cout(Xd_0__inst_mult_30_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_294 ),
	.datab(!Xd_0__inst_mult_5_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_205 ),
	.cout(Xd_0__inst_mult_5_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_26 (
// Equation(s):

	.dataa(!din_a[143]),
	.datab(!din_b[143]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_32 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_26_sumout ),
	.cout(Xd_0__inst_i29_27 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_85 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[208]),
	.datac(!Xd_0__inst_mult_17_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_219 ),
	.cout(Xd_0__inst_mult_17_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_40 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[207]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_40_sumout ),
	.cout(Xd_0__inst_mult_17_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_219 ),
	.datab(!Xd_0__inst_mult_17_40_sumout ),
	.datac(!Xd_0__inst_mult_17_324 ),
	.datad(!Xd_0__inst_mult_17_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_224 ),
	.cout(Xd_0__inst_mult_17_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_95 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[327]),
	.datac(!din_a[331]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_269 ),
	.cout(Xd_0__inst_mult_27_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_96 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_374 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_274 ),
	.cout(Xd_0__inst_mult_27_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_97 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[325]),
	.datac(!din_a[334]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_279 ),
	.cout(Xd_0__inst_mult_27_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_279 ),
	.datab(!Xd_0__inst_mult_27_274 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_284 ),
	.cout(Xd_0__inst_mult_27_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_294 ),
	.datab(!Xd_0__inst_mult_13_45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_205 ),
	.cout(Xd_0__inst_mult_13_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_344 ),
	.datab(!Xd_0__inst_mult_2_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_249 ),
	.cout(Xd_0__inst_mult_2_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_31 (
// Equation(s):

	.dataa(!din_a[95]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_31_sumout ),
	.cout(Xd_0__inst_i29_32 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_85 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[196]),
	.datac(!Xd_0__inst_mult_16_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_219 ),
	.cout(Xd_0__inst_mult_16_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_40 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[195]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_40_sumout ),
	.cout(Xd_0__inst_mult_16_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_219 ),
	.datab(!Xd_0__inst_mult_16_40_sumout ),
	.datac(!Xd_0__inst_mult_16_324 ),
	.datad(!Xd_0__inst_mult_16_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_224 ),
	.cout(Xd_0__inst_mult_16_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_294 ),
	.datab(!Xd_0__inst_mult_28_40_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_205 ),
	.cout(Xd_0__inst_mult_28_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_294 ),
	.datab(!Xd_0__inst_mult_31_40_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_205 ),
	.cout(Xd_0__inst_mult_31_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_36 (
// Equation(s):

	.dataa(!din_a[47]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_42 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_36_sumout ),
	.cout(Xd_0__inst_i29_37 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_85 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[352]),
	.datac(!Xd_0__inst_mult_29_314 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_219 ),
	.cout(Xd_0__inst_mult_29_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_40 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[351]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_40_sumout ),
	.cout(Xd_0__inst_mult_29_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_219 ),
	.datab(!Xd_0__inst_mult_29_40_sumout ),
	.datac(!Xd_0__inst_mult_29_324 ),
	.datad(!Xd_0__inst_mult_29_319 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_224 ),
	.cout(Xd_0__inst_mult_29_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_123 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[315]),
	.datac(!din_a[319]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_409 ),
	.cout(Xd_0__inst_mult_26_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_124 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_539 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_414 ),
	.cout(Xd_0__inst_mult_26_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_125 (
// Equation(s):

	.dataa(!din_a[321]),
	.datab(!din_b[313]),
	.datac(!din_a[322]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_419 ),
	.cout(Xd_0__inst_mult_26_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_419 ),
	.datab(!Xd_0__inst_mult_26_414 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_424 ),
	.cout(Xd_0__inst_mult_26_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_122 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[297]),
	.datac(!din_a[292]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_404 ),
	.cout(Xd_0__inst_mult_24_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_123 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_534 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_409 ),
	.cout(Xd_0__inst_mult_24_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_124 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[294]),
	.datac(!din_a[295]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_414 ),
	.cout(Xd_0__inst_mult_24_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_125 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_419 ),
	.cout(Xd_0__inst_mult_24_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_419 ),
	.datab(!Xd_0__inst_mult_24_409 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_424 ),
	.cout(Xd_0__inst_mult_24_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_92 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[29]),
	.datac(!din_a[24]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_254 ),
	.cout(Xd_0__inst_mult_2_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_0_q ),
	.datab(!Xd_0__inst_mult_29_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_229 ),
	.cout(Xd_0__inst_mult_29_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_0_q ),
	.datab(!Xd_0__inst_mult_28_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_210 ),
	.cout(Xd_0__inst_mult_28_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_0_q ),
	.datab(!Xd_0__inst_mult_31_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_210 ),
	.cout(Xd_0__inst_mult_31_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_0_q ),
	.datab(!Xd_0__inst_mult_30_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_210 ),
	.cout(Xd_0__inst_mult_30_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_0_q ),
	.datab(!Xd_0__inst_mult_25_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_289 ),
	.cout(Xd_0__inst_mult_25_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_0_q ),
	.datab(!Xd_0__inst_mult_24_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_429 ),
	.cout(Xd_0__inst_mult_24_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_0_q ),
	.datab(!Xd_0__inst_mult_27_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_289 ),
	.cout(Xd_0__inst_mult_27_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_0_q ),
	.datab(!Xd_0__inst_mult_26_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_429 ),
	.cout(Xd_0__inst_mult_26_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_0_q ),
	.datab(!Xd_0__inst_mult_21_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_229 ),
	.cout(Xd_0__inst_mult_21_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_0_q ),
	.datab(!Xd_0__inst_mult_20_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_229 ),
	.cout(Xd_0__inst_mult_20_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_0_q ),
	.datab(!Xd_0__inst_mult_23_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_229 ),
	.cout(Xd_0__inst_mult_23_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_0_q ),
	.datab(!Xd_0__inst_mult_22_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_229 ),
	.cout(Xd_0__inst_mult_22_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_0_q ),
	.datab(!Xd_0__inst_mult_17_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_229 ),
	.cout(Xd_0__inst_mult_17_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_0_q ),
	.datab(!Xd_0__inst_mult_16_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_229 ),
	.cout(Xd_0__inst_mult_16_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_0_q ),
	.datab(!Xd_0__inst_mult_19_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_229 ),
	.cout(Xd_0__inst_mult_19_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_0_q ),
	.datab(!Xd_0__inst_mult_18_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_205 ),
	.cout(Xd_0__inst_mult_18_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_210 ),
	.cout(Xd_0__inst_mult_13_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_205 ),
	.cout(Xd_0__inst_mult_12_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_205 ),
	.cout(Xd_0__inst_mult_15_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_204 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_205 ),
	.cout(Xd_0__inst_mult_14_206 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_210 ),
	.cout(Xd_0__inst_mult_9_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_210 ),
	.cout(Xd_0__inst_mult_8_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_0_q ),
	.datab(!Xd_0__inst_mult_11_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_210 ),
	.cout(Xd_0__inst_mult_11_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_210 ),
	.cout(Xd_0__inst_mult_10_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_210 ),
	.cout(Xd_0__inst_mult_5_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_210 ),
	.cout(Xd_0__inst_mult_4_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_210 ),
	.cout(Xd_0__inst_mult_7_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_210 ),
	.cout(Xd_0__inst_mult_6_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_210 ),
	.cout(Xd_0__inst_mult_1_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_210 ),
	.cout(Xd_0__inst_mult_0_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_210 ),
	.cout(Xd_0__inst_mult_3_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_259 ),
	.cout(Xd_0__inst_mult_2_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_2_q ),
	.datab(!Xd_0__inst_mult_29_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_234 ),
	.cout(Xd_0__inst_mult_29_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_2_q ),
	.datab(!Xd_0__inst_mult_28_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_214 ),
	.cout(Xd_0__inst_mult_28_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_2_q ),
	.datab(!Xd_0__inst_mult_31_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_214 ),
	.cout(Xd_0__inst_mult_31_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_2_q ),
	.datab(!Xd_0__inst_mult_30_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_214 ),
	.cout(Xd_0__inst_mult_30_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_2_q ),
	.datab(!Xd_0__inst_mult_25_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_294 ),
	.cout(Xd_0__inst_mult_25_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_2_q ),
	.datab(!Xd_0__inst_mult_24_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_434 ),
	.cout(Xd_0__inst_mult_24_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_2_q ),
	.datab(!Xd_0__inst_mult_27_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_294 ),
	.cout(Xd_0__inst_mult_27_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_2_q ),
	.datab(!Xd_0__inst_mult_26_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_434 ),
	.cout(Xd_0__inst_mult_26_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_2_q ),
	.datab(!Xd_0__inst_mult_21_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_234 ),
	.cout(Xd_0__inst_mult_21_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_2_q ),
	.datab(!Xd_0__inst_mult_20_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_234 ),
	.cout(Xd_0__inst_mult_20_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_2_q ),
	.datab(!Xd_0__inst_mult_23_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_234 ),
	.cout(Xd_0__inst_mult_23_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_2_q ),
	.datab(!Xd_0__inst_mult_22_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_234 ),
	.cout(Xd_0__inst_mult_22_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_2_q ),
	.datab(!Xd_0__inst_mult_17_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_234 ),
	.cout(Xd_0__inst_mult_17_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_2_q ),
	.datab(!Xd_0__inst_mult_16_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_234 ),
	.cout(Xd_0__inst_mult_16_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_2_q ),
	.datab(!Xd_0__inst_mult_19_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_234 ),
	.cout(Xd_0__inst_mult_19_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_2_q ),
	.datab(!Xd_0__inst_mult_18_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_210 ),
	.cout(Xd_0__inst_mult_18_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_2_q ),
	.datab(!Xd_0__inst_mult_13_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_214 ),
	.cout(Xd_0__inst_mult_13_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_2_q ),
	.datab(!Xd_0__inst_mult_12_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_210 ),
	.cout(Xd_0__inst_mult_12_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_2_q ),
	.datab(!Xd_0__inst_mult_15_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_210 ),
	.cout(Xd_0__inst_mult_15_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_2_q ),
	.datab(!Xd_0__inst_mult_14_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_206 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_210 ),
	.cout(Xd_0__inst_mult_14_211 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_2_q ),
	.datab(!Xd_0__inst_mult_9_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_214 ),
	.cout(Xd_0__inst_mult_9_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_2_q ),
	.datab(!Xd_0__inst_mult_8_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_214 ),
	.cout(Xd_0__inst_mult_8_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_2_q ),
	.datab(!Xd_0__inst_mult_11_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_214 ),
	.cout(Xd_0__inst_mult_11_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_2_q ),
	.datab(!Xd_0__inst_mult_10_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_214 ),
	.cout(Xd_0__inst_mult_10_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_2_q ),
	.datab(!Xd_0__inst_mult_5_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_214 ),
	.cout(Xd_0__inst_mult_5_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_2_q ),
	.datab(!Xd_0__inst_mult_4_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_214 ),
	.cout(Xd_0__inst_mult_4_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_2_q ),
	.datab(!Xd_0__inst_mult_7_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_214 ),
	.cout(Xd_0__inst_mult_7_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_2_q ),
	.datab(!Xd_0__inst_mult_6_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_214 ),
	.cout(Xd_0__inst_mult_6_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_2_q ),
	.datab(!Xd_0__inst_mult_1_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_214 ),
	.cout(Xd_0__inst_mult_1_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_2_q ),
	.datab(!Xd_0__inst_mult_0_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_214 ),
	.cout(Xd_0__inst_mult_0_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_2_q ),
	.datab(!Xd_0__inst_mult_3_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_214 ),
	.cout(Xd_0__inst_mult_3_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_2_q ),
	.datab(!Xd_0__inst_mult_2_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_264 ),
	.cout(Xd_0__inst_mult_2_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_239 ),
	.cout(Xd_0__inst_mult_29_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_219 ),
	.cout(Xd_0__inst_mult_28_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_219 ),
	.cout(Xd_0__inst_mult_31_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_219 ),
	.cout(Xd_0__inst_mult_30_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_299 ),
	.cout(Xd_0__inst_mult_25_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_439 ),
	.cout(Xd_0__inst_mult_24_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_299 ),
	.cout(Xd_0__inst_mult_27_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_439 ),
	.cout(Xd_0__inst_mult_26_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_239 ),
	.cout(Xd_0__inst_mult_21_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_239 ),
	.cout(Xd_0__inst_mult_20_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_239 ),
	.cout(Xd_0__inst_mult_23_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_239 ),
	.cout(Xd_0__inst_mult_22_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_239 ),
	.cout(Xd_0__inst_mult_17_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_239 ),
	.cout(Xd_0__inst_mult_16_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_239 ),
	.cout(Xd_0__inst_mult_19_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_214 ),
	.cout(Xd_0__inst_mult_18_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_219 ),
	.cout(Xd_0__inst_mult_13_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_214 ),
	.cout(Xd_0__inst_mult_12_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_214 ),
	.cout(Xd_0__inst_mult_15_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_84 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_211 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_214 ),
	.cout(Xd_0__inst_mult_14_215 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_219 ),
	.cout(Xd_0__inst_mult_9_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_219 ),
	.cout(Xd_0__inst_mult_8_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_219 ),
	.cout(Xd_0__inst_mult_11_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_219 ),
	.cout(Xd_0__inst_mult_10_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_219 ),
	.cout(Xd_0__inst_mult_5_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_219 ),
	.cout(Xd_0__inst_mult_4_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_219 ),
	.cout(Xd_0__inst_mult_7_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_219 ),
	.cout(Xd_0__inst_mult_6_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_219 ),
	.cout(Xd_0__inst_mult_1_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_219 ),
	.cout(Xd_0__inst_mult_0_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_219 ),
	.cout(Xd_0__inst_mult_3_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_269 ),
	.cout(Xd_0__inst_mult_2_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_6_q ),
	.datab(!Xd_0__inst_mult_29_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_244 ),
	.cout(Xd_0__inst_mult_29_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_6_q ),
	.datab(!Xd_0__inst_mult_28_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_224 ),
	.cout(Xd_0__inst_mult_28_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_6_q ),
	.datab(!Xd_0__inst_mult_31_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_224 ),
	.cout(Xd_0__inst_mult_31_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_6_q ),
	.datab(!Xd_0__inst_mult_30_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_224 ),
	.cout(Xd_0__inst_mult_30_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_6_q ),
	.datab(!Xd_0__inst_mult_25_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_304 ),
	.cout(Xd_0__inst_mult_25_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_6_q ),
	.datab(!Xd_0__inst_mult_24_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_444 ),
	.cout(Xd_0__inst_mult_24_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_6_q ),
	.datab(!Xd_0__inst_mult_27_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_304 ),
	.cout(Xd_0__inst_mult_27_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_6_q ),
	.datab(!Xd_0__inst_mult_26_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_444 ),
	.cout(Xd_0__inst_mult_26_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_6_q ),
	.datab(!Xd_0__inst_mult_21_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_244 ),
	.cout(Xd_0__inst_mult_21_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_6_q ),
	.datab(!Xd_0__inst_mult_20_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_244 ),
	.cout(Xd_0__inst_mult_20_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_6_q ),
	.datab(!Xd_0__inst_mult_23_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_244 ),
	.cout(Xd_0__inst_mult_23_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_6_q ),
	.datab(!Xd_0__inst_mult_22_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_244 ),
	.cout(Xd_0__inst_mult_22_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_6_q ),
	.datab(!Xd_0__inst_mult_17_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_244 ),
	.cout(Xd_0__inst_mult_17_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_6_q ),
	.datab(!Xd_0__inst_mult_16_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_244 ),
	.cout(Xd_0__inst_mult_16_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_6_q ),
	.datab(!Xd_0__inst_mult_19_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_244 ),
	.cout(Xd_0__inst_mult_19_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_6_q ),
	.datab(!Xd_0__inst_mult_18_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_219 ),
	.cout(Xd_0__inst_mult_18_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_6_q ),
	.datab(!Xd_0__inst_mult_13_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_224 ),
	.cout(Xd_0__inst_mult_13_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_6_q ),
	.datab(!Xd_0__inst_mult_12_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_219 ),
	.cout(Xd_0__inst_mult_12_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_6_q ),
	.datab(!Xd_0__inst_mult_15_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_219 ),
	.cout(Xd_0__inst_mult_15_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_85 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_6_q ),
	.datab(!Xd_0__inst_mult_14_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_215 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_219 ),
	.cout(Xd_0__inst_mult_14_220 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_6_q ),
	.datab(!Xd_0__inst_mult_9_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_224 ),
	.cout(Xd_0__inst_mult_9_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_6_q ),
	.datab(!Xd_0__inst_mult_8_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_224 ),
	.cout(Xd_0__inst_mult_8_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_6_q ),
	.datab(!Xd_0__inst_mult_11_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_224 ),
	.cout(Xd_0__inst_mult_11_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_6_q ),
	.datab(!Xd_0__inst_mult_10_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_224 ),
	.cout(Xd_0__inst_mult_10_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_6_q ),
	.datab(!Xd_0__inst_mult_5_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_224 ),
	.cout(Xd_0__inst_mult_5_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_6_q ),
	.datab(!Xd_0__inst_mult_4_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_224 ),
	.cout(Xd_0__inst_mult_4_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_6_q ),
	.datab(!Xd_0__inst_mult_7_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_224 ),
	.cout(Xd_0__inst_mult_7_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_6_q ),
	.datab(!Xd_0__inst_mult_6_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_224 ),
	.cout(Xd_0__inst_mult_6_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_6_q ),
	.datab(!Xd_0__inst_mult_1_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_224 ),
	.cout(Xd_0__inst_mult_1_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_6_q ),
	.datab(!Xd_0__inst_mult_0_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_224 ),
	.cout(Xd_0__inst_mult_0_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_6_q ),
	.datab(!Xd_0__inst_mult_3_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_224 ),
	.cout(Xd_0__inst_mult_3_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_6_q ),
	.datab(!Xd_0__inst_mult_2_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_274 ),
	.cout(Xd_0__inst_mult_2_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_8_q ),
	.datab(!Xd_0__inst_mult_29_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_249 ),
	.cout(Xd_0__inst_mult_29_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_8_q ),
	.datab(!Xd_0__inst_mult_28_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_229 ),
	.cout(Xd_0__inst_mult_28_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_8_q ),
	.datab(!Xd_0__inst_mult_31_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_229 ),
	.cout(Xd_0__inst_mult_31_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_8_q ),
	.datab(!Xd_0__inst_mult_30_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_229 ),
	.cout(Xd_0__inst_mult_30_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_8_q ),
	.datab(!Xd_0__inst_mult_25_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_309 ),
	.cout(Xd_0__inst_mult_25_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_8_q ),
	.datab(!Xd_0__inst_mult_24_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_449 ),
	.cout(Xd_0__inst_mult_24_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_8_q ),
	.datab(!Xd_0__inst_mult_27_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_309 ),
	.cout(Xd_0__inst_mult_27_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_8_q ),
	.datab(!Xd_0__inst_mult_26_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_449 ),
	.cout(Xd_0__inst_mult_26_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_8_q ),
	.datab(!Xd_0__inst_mult_21_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_249 ),
	.cout(Xd_0__inst_mult_21_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_8_q ),
	.datab(!Xd_0__inst_mult_20_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_249 ),
	.cout(Xd_0__inst_mult_20_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_8_q ),
	.datab(!Xd_0__inst_mult_23_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_249 ),
	.cout(Xd_0__inst_mult_23_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_8_q ),
	.datab(!Xd_0__inst_mult_22_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_249 ),
	.cout(Xd_0__inst_mult_22_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_8_q ),
	.datab(!Xd_0__inst_mult_17_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_249 ),
	.cout(Xd_0__inst_mult_17_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_8_q ),
	.datab(!Xd_0__inst_mult_16_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_249 ),
	.cout(Xd_0__inst_mult_16_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_8_q ),
	.datab(!Xd_0__inst_mult_19_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_249 ),
	.cout(Xd_0__inst_mult_19_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_8_q ),
	.datab(!Xd_0__inst_mult_18_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_224 ),
	.cout(Xd_0__inst_mult_18_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_8_q ),
	.datab(!Xd_0__inst_mult_13_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_229 ),
	.cout(Xd_0__inst_mult_13_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_8_q ),
	.datab(!Xd_0__inst_mult_12_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_224 ),
	.cout(Xd_0__inst_mult_12_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_8_q ),
	.datab(!Xd_0__inst_mult_15_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_224 ),
	.cout(Xd_0__inst_mult_15_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_86 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_8_q ),
	.datab(!Xd_0__inst_mult_14_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_220 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_224 ),
	.cout(Xd_0__inst_mult_14_225 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_8_q ),
	.datab(!Xd_0__inst_mult_9_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_229 ),
	.cout(Xd_0__inst_mult_9_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_8_q ),
	.datab(!Xd_0__inst_mult_8_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_229 ),
	.cout(Xd_0__inst_mult_8_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_8_q ),
	.datab(!Xd_0__inst_mult_11_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_229 ),
	.cout(Xd_0__inst_mult_11_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_8_q ),
	.datab(!Xd_0__inst_mult_10_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_229 ),
	.cout(Xd_0__inst_mult_10_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_229 ),
	.cout(Xd_0__inst_mult_5_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_229 ),
	.cout(Xd_0__inst_mult_4_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_229 ),
	.cout(Xd_0__inst_mult_7_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_229 ),
	.cout(Xd_0__inst_mult_6_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_229 ),
	.cout(Xd_0__inst_mult_1_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_229 ),
	.cout(Xd_0__inst_mult_0_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_229 ),
	.cout(Xd_0__inst_mult_3_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_279 ),
	.cout(Xd_0__inst_mult_2_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_10_q ),
	.datab(!Xd_0__inst_mult_29_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_254 ),
	.cout(Xd_0__inst_mult_29_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_10_q ),
	.datab(!Xd_0__inst_mult_28_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_234 ),
	.cout(Xd_0__inst_mult_28_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_10_q ),
	.datab(!Xd_0__inst_mult_31_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_234 ),
	.cout(Xd_0__inst_mult_31_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_10_q ),
	.datab(!Xd_0__inst_mult_30_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_234 ),
	.cout(Xd_0__inst_mult_30_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_10_q ),
	.datab(!Xd_0__inst_mult_25_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_314 ),
	.cout(Xd_0__inst_mult_25_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_10_q ),
	.datab(!Xd_0__inst_mult_24_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_454 ),
	.cout(Xd_0__inst_mult_24_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_10_q ),
	.datab(!Xd_0__inst_mult_27_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_314 ),
	.cout(Xd_0__inst_mult_27_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_10_q ),
	.datab(!Xd_0__inst_mult_26_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_454 ),
	.cout(Xd_0__inst_mult_26_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_10_q ),
	.datab(!Xd_0__inst_mult_21_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_254 ),
	.cout(Xd_0__inst_mult_21_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_10_q ),
	.datab(!Xd_0__inst_mult_20_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_254 ),
	.cout(Xd_0__inst_mult_20_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_10_q ),
	.datab(!Xd_0__inst_mult_23_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_254 ),
	.cout(Xd_0__inst_mult_23_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_10_q ),
	.datab(!Xd_0__inst_mult_22_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_254 ),
	.cout(Xd_0__inst_mult_22_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_10_q ),
	.datab(!Xd_0__inst_mult_17_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_254 ),
	.cout(Xd_0__inst_mult_17_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_10_q ),
	.datab(!Xd_0__inst_mult_16_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_254 ),
	.cout(Xd_0__inst_mult_16_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_10_q ),
	.datab(!Xd_0__inst_mult_19_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_254 ),
	.cout(Xd_0__inst_mult_19_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_10_q ),
	.datab(!Xd_0__inst_mult_18_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_229 ),
	.cout(Xd_0__inst_mult_18_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_10_q ),
	.datab(!Xd_0__inst_mult_13_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_234 ),
	.cout(Xd_0__inst_mult_13_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_10_q ),
	.datab(!Xd_0__inst_mult_12_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_229 ),
	.cout(Xd_0__inst_mult_12_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_10_q ),
	.datab(!Xd_0__inst_mult_15_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_229 ),
	.cout(Xd_0__inst_mult_15_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_87 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_10_q ),
	.datab(!Xd_0__inst_mult_14_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_225 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_229 ),
	.cout(Xd_0__inst_mult_14_230 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_10_q ),
	.datab(!Xd_0__inst_mult_9_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_234 ),
	.cout(Xd_0__inst_mult_9_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_10_q ),
	.datab(!Xd_0__inst_mult_8_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_234 ),
	.cout(Xd_0__inst_mult_8_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_10_q ),
	.datab(!Xd_0__inst_mult_11_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_234 ),
	.cout(Xd_0__inst_mult_11_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_10_q ),
	.datab(!Xd_0__inst_mult_10_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_234 ),
	.cout(Xd_0__inst_mult_10_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_10_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_234 ),
	.cout(Xd_0__inst_mult_5_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_10_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_234 ),
	.cout(Xd_0__inst_mult_4_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_10_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_234 ),
	.cout(Xd_0__inst_mult_7_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_10_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_234 ),
	.cout(Xd_0__inst_mult_6_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_10_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_234 ),
	.cout(Xd_0__inst_mult_1_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_10_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_234 ),
	.cout(Xd_0__inst_mult_0_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_10_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_234 ),
	.cout(Xd_0__inst_mult_3_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_10_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_284 ),
	.cout(Xd_0__inst_mult_2_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_12_q ),
	.datab(!Xd_0__inst_mult_29_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_259 ),
	.cout(Xd_0__inst_mult_29_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_12_q ),
	.datab(!Xd_0__inst_mult_28_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_239 ),
	.cout(Xd_0__inst_mult_28_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_12_q ),
	.datab(!Xd_0__inst_mult_31_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_239 ),
	.cout(Xd_0__inst_mult_31_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_12_q ),
	.datab(!Xd_0__inst_mult_30_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_239 ),
	.cout(Xd_0__inst_mult_30_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_12_q ),
	.datab(!Xd_0__inst_mult_25_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_319 ),
	.cout(Xd_0__inst_mult_25_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_12_q ),
	.datab(!Xd_0__inst_mult_24_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_459 ),
	.cout(Xd_0__inst_mult_24_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_12_q ),
	.datab(!Xd_0__inst_mult_27_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_319 ),
	.cout(Xd_0__inst_mult_27_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_12_q ),
	.datab(!Xd_0__inst_mult_26_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_459 ),
	.cout(Xd_0__inst_mult_26_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_12_q ),
	.datab(!Xd_0__inst_mult_21_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_259 ),
	.cout(Xd_0__inst_mult_21_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_12_q ),
	.datab(!Xd_0__inst_mult_20_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_259 ),
	.cout(Xd_0__inst_mult_20_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_12_q ),
	.datab(!Xd_0__inst_mult_23_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_259 ),
	.cout(Xd_0__inst_mult_23_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_12_q ),
	.datab(!Xd_0__inst_mult_22_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_259 ),
	.cout(Xd_0__inst_mult_22_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_12_q ),
	.datab(!Xd_0__inst_mult_17_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_259 ),
	.cout(Xd_0__inst_mult_17_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_12_q ),
	.datab(!Xd_0__inst_mult_16_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_259 ),
	.cout(Xd_0__inst_mult_16_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_12_q ),
	.datab(!Xd_0__inst_mult_19_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_259 ),
	.cout(Xd_0__inst_mult_19_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_12_q ),
	.datab(!Xd_0__inst_mult_18_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_234 ),
	.cout(Xd_0__inst_mult_18_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_12_q ),
	.datab(!Xd_0__inst_mult_13_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_239 ),
	.cout(Xd_0__inst_mult_13_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_12_q ),
	.datab(!Xd_0__inst_mult_12_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_234 ),
	.cout(Xd_0__inst_mult_12_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_12_q ),
	.datab(!Xd_0__inst_mult_15_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_234 ),
	.cout(Xd_0__inst_mult_15_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_88 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_12_q ),
	.datab(!Xd_0__inst_mult_14_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_230 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_234 ),
	.cout(Xd_0__inst_mult_14_235 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_12_q ),
	.datab(!Xd_0__inst_mult_9_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_239 ),
	.cout(Xd_0__inst_mult_9_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_12_q ),
	.datab(!Xd_0__inst_mult_8_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_239 ),
	.cout(Xd_0__inst_mult_8_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_12_q ),
	.datab(!Xd_0__inst_mult_11_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_239 ),
	.cout(Xd_0__inst_mult_11_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_12_q ),
	.datab(!Xd_0__inst_mult_10_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_239 ),
	.cout(Xd_0__inst_mult_10_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_12_q ),
	.datab(!Xd_0__inst_mult_5_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_239 ),
	.cout(Xd_0__inst_mult_5_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_12_q ),
	.datab(!Xd_0__inst_mult_4_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_239 ),
	.cout(Xd_0__inst_mult_4_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_12_q ),
	.datab(!Xd_0__inst_mult_7_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_239 ),
	.cout(Xd_0__inst_mult_7_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_12_q ),
	.datab(!Xd_0__inst_mult_6_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_239 ),
	.cout(Xd_0__inst_mult_6_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_12_q ),
	.datab(!Xd_0__inst_mult_1_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_239 ),
	.cout(Xd_0__inst_mult_1_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_12_q ),
	.datab(!Xd_0__inst_mult_0_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_239 ),
	.cout(Xd_0__inst_mult_0_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_12_q ),
	.datab(!Xd_0__inst_mult_3_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_239 ),
	.cout(Xd_0__inst_mult_3_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_12_q ),
	.datab(!Xd_0__inst_mult_2_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_289 ),
	.cout(Xd_0__inst_mult_2_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_14_q ),
	.datab(!Xd_0__inst_mult_29_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_264 ),
	.cout(Xd_0__inst_mult_29_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_14_q ),
	.datab(!Xd_0__inst_mult_28_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_244 ),
	.cout(Xd_0__inst_mult_28_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_14_q ),
	.datab(!Xd_0__inst_mult_31_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_244 ),
	.cout(Xd_0__inst_mult_31_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_14_q ),
	.datab(!Xd_0__inst_mult_30_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_244 ),
	.cout(Xd_0__inst_mult_30_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_106 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_14_q ),
	.datab(!Xd_0__inst_mult_25_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_324 ),
	.cout(Xd_0__inst_mult_25_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_14_q ),
	.datab(!Xd_0__inst_mult_24_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_464 ),
	.cout(Xd_0__inst_mult_24_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_106 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_14_q ),
	.datab(!Xd_0__inst_mult_27_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_324 ),
	.cout(Xd_0__inst_mult_27_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_14_q ),
	.datab(!Xd_0__inst_mult_26_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_464 ),
	.cout(Xd_0__inst_mult_26_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_14_q ),
	.datab(!Xd_0__inst_mult_21_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_264 ),
	.cout(Xd_0__inst_mult_21_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_14_q ),
	.datab(!Xd_0__inst_mult_20_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_264 ),
	.cout(Xd_0__inst_mult_20_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_14_q ),
	.datab(!Xd_0__inst_mult_23_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_264 ),
	.cout(Xd_0__inst_mult_23_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_14_q ),
	.datab(!Xd_0__inst_mult_22_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_264 ),
	.cout(Xd_0__inst_mult_22_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_14_q ),
	.datab(!Xd_0__inst_mult_17_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_264 ),
	.cout(Xd_0__inst_mult_17_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_14_q ),
	.datab(!Xd_0__inst_mult_16_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_264 ),
	.cout(Xd_0__inst_mult_16_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_14_q ),
	.datab(!Xd_0__inst_mult_19_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_264 ),
	.cout(Xd_0__inst_mult_19_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_14_q ),
	.datab(!Xd_0__inst_mult_18_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_239 ),
	.cout(Xd_0__inst_mult_18_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_14_q ),
	.datab(!Xd_0__inst_mult_13_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_244 ),
	.cout(Xd_0__inst_mult_13_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_14_q ),
	.datab(!Xd_0__inst_mult_12_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_239 ),
	.cout(Xd_0__inst_mult_12_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_14_q ),
	.datab(!Xd_0__inst_mult_15_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_239 ),
	.cout(Xd_0__inst_mult_15_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_89 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_14_q ),
	.datab(!Xd_0__inst_mult_14_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_239 ),
	.cout(Xd_0__inst_mult_14_240 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_14_q ),
	.datab(!Xd_0__inst_mult_9_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_244 ),
	.cout(Xd_0__inst_mult_9_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_14_q ),
	.datab(!Xd_0__inst_mult_8_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_244 ),
	.cout(Xd_0__inst_mult_8_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_14_q ),
	.datab(!Xd_0__inst_mult_11_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_244 ),
	.cout(Xd_0__inst_mult_11_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_14_q ),
	.datab(!Xd_0__inst_mult_10_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_244 ),
	.cout(Xd_0__inst_mult_10_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_14_q ),
	.datab(!Xd_0__inst_mult_5_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_244 ),
	.cout(Xd_0__inst_mult_5_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_14_q ),
	.datab(!Xd_0__inst_mult_4_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_244 ),
	.cout(Xd_0__inst_mult_4_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_14_q ),
	.datab(!Xd_0__inst_mult_7_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_244 ),
	.cout(Xd_0__inst_mult_7_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_14_q ),
	.datab(!Xd_0__inst_mult_6_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_244 ),
	.cout(Xd_0__inst_mult_6_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_14_q ),
	.datab(!Xd_0__inst_mult_1_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_244 ),
	.cout(Xd_0__inst_mult_1_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_14_q ),
	.datab(!Xd_0__inst_mult_0_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_244 ),
	.cout(Xd_0__inst_mult_0_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_14_q ),
	.datab(!Xd_0__inst_mult_3_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_244 ),
	.cout(Xd_0__inst_mult_3_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_14_q ),
	.datab(!Xd_0__inst_mult_2_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_294 ),
	.cout(Xd_0__inst_mult_2_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_16_q ),
	.datab(!Xd_0__inst_mult_29_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_269 ),
	.cout(Xd_0__inst_mult_29_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_16_q ),
	.datab(!Xd_0__inst_mult_28_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_249 ),
	.cout(Xd_0__inst_mult_28_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_16_q ),
	.datab(!Xd_0__inst_mult_31_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_249 ),
	.cout(Xd_0__inst_mult_31_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_16_q ),
	.datab(!Xd_0__inst_mult_30_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_249 ),
	.cout(Xd_0__inst_mult_30_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_16_q ),
	.datab(!Xd_0__inst_mult_25_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_329 ),
	.cout(Xd_0__inst_mult_25_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_16_q ),
	.datab(!Xd_0__inst_mult_24_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_469 ),
	.cout(Xd_0__inst_mult_24_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_16_q ),
	.datab(!Xd_0__inst_mult_27_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_329 ),
	.cout(Xd_0__inst_mult_27_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_16_q ),
	.datab(!Xd_0__inst_mult_26_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_469 ),
	.cout(Xd_0__inst_mult_26_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_16_q ),
	.datab(!Xd_0__inst_mult_21_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_269 ),
	.cout(Xd_0__inst_mult_21_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_16_q ),
	.datab(!Xd_0__inst_mult_20_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_269 ),
	.cout(Xd_0__inst_mult_20_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_16_q ),
	.datab(!Xd_0__inst_mult_23_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_269 ),
	.cout(Xd_0__inst_mult_23_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_16_q ),
	.datab(!Xd_0__inst_mult_22_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_269 ),
	.cout(Xd_0__inst_mult_22_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_16_q ),
	.datab(!Xd_0__inst_mult_17_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_269 ),
	.cout(Xd_0__inst_mult_17_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_16_q ),
	.datab(!Xd_0__inst_mult_16_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_269 ),
	.cout(Xd_0__inst_mult_16_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_16_q ),
	.datab(!Xd_0__inst_mult_19_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_269 ),
	.cout(Xd_0__inst_mult_19_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_16_q ),
	.datab(!Xd_0__inst_mult_18_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_244 ),
	.cout(Xd_0__inst_mult_18_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_16_q ),
	.datab(!Xd_0__inst_mult_13_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_249 ),
	.cout(Xd_0__inst_mult_13_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_16_q ),
	.datab(!Xd_0__inst_mult_12_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_244 ),
	.cout(Xd_0__inst_mult_12_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_16_q ),
	.datab(!Xd_0__inst_mult_15_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_244 ),
	.cout(Xd_0__inst_mult_15_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_90 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_16_q ),
	.datab(!Xd_0__inst_mult_14_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_240 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_244 ),
	.cout(Xd_0__inst_mult_14_245 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_16_q ),
	.datab(!Xd_0__inst_mult_9_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_249 ),
	.cout(Xd_0__inst_mult_9_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_16_q ),
	.datab(!Xd_0__inst_mult_8_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_249 ),
	.cout(Xd_0__inst_mult_8_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_16_q ),
	.datab(!Xd_0__inst_mult_11_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_249 ),
	.cout(Xd_0__inst_mult_11_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_16_q ),
	.datab(!Xd_0__inst_mult_10_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_249 ),
	.cout(Xd_0__inst_mult_10_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_16_q ),
	.datab(!Xd_0__inst_mult_5_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_249 ),
	.cout(Xd_0__inst_mult_5_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_16_q ),
	.datab(!Xd_0__inst_mult_4_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_249 ),
	.cout(Xd_0__inst_mult_4_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_16_q ),
	.datab(!Xd_0__inst_mult_7_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_249 ),
	.cout(Xd_0__inst_mult_7_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_16_q ),
	.datab(!Xd_0__inst_mult_6_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_249 ),
	.cout(Xd_0__inst_mult_6_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_16_q ),
	.datab(!Xd_0__inst_mult_1_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_249 ),
	.cout(Xd_0__inst_mult_1_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_16_q ),
	.datab(!Xd_0__inst_mult_0_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_249 ),
	.cout(Xd_0__inst_mult_0_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_16_q ),
	.datab(!Xd_0__inst_mult_3_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_249 ),
	.cout(Xd_0__inst_mult_3_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_16_q ),
	.datab(!Xd_0__inst_mult_2_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_299 ),
	.cout(Xd_0__inst_mult_2_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_18_q ),
	.datab(!Xd_0__inst_mult_29_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_274 ),
	.cout(Xd_0__inst_mult_29_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_18_q ),
	.datab(!Xd_0__inst_mult_28_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_254 ),
	.cout(Xd_0__inst_mult_28_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_18_q ),
	.datab(!Xd_0__inst_mult_31_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_254 ),
	.cout(Xd_0__inst_mult_31_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_18_q ),
	.datab(!Xd_0__inst_mult_30_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_254 ),
	.cout(Xd_0__inst_mult_30_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_108 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_18_q ),
	.datab(!Xd_0__inst_mult_25_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_334 ),
	.cout(Xd_0__inst_mult_25_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_18_q ),
	.datab(!Xd_0__inst_mult_24_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_474 ),
	.cout(Xd_0__inst_mult_24_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_108 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_18_q ),
	.datab(!Xd_0__inst_mult_27_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_334 ),
	.cout(Xd_0__inst_mult_27_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_18_q ),
	.datab(!Xd_0__inst_mult_26_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_474 ),
	.cout(Xd_0__inst_mult_26_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_18_q ),
	.datab(!Xd_0__inst_mult_21_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_274 ),
	.cout(Xd_0__inst_mult_21_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_18_q ),
	.datab(!Xd_0__inst_mult_20_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_274 ),
	.cout(Xd_0__inst_mult_20_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_18_q ),
	.datab(!Xd_0__inst_mult_23_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_274 ),
	.cout(Xd_0__inst_mult_23_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_18_q ),
	.datab(!Xd_0__inst_mult_22_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_274 ),
	.cout(Xd_0__inst_mult_22_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_18_q ),
	.datab(!Xd_0__inst_mult_17_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_274 ),
	.cout(Xd_0__inst_mult_17_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_18_q ),
	.datab(!Xd_0__inst_mult_16_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_274 ),
	.cout(Xd_0__inst_mult_16_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_18_q ),
	.datab(!Xd_0__inst_mult_19_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_274 ),
	.cout(Xd_0__inst_mult_19_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_18_q ),
	.datab(!Xd_0__inst_mult_18_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_249 ),
	.cout(Xd_0__inst_mult_18_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_18_q ),
	.datab(!Xd_0__inst_mult_13_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_254 ),
	.cout(Xd_0__inst_mult_13_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_18_q ),
	.datab(!Xd_0__inst_mult_12_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_249 ),
	.cout(Xd_0__inst_mult_12_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_18_q ),
	.datab(!Xd_0__inst_mult_15_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_249 ),
	.cout(Xd_0__inst_mult_15_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_91 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_18_q ),
	.datab(!Xd_0__inst_mult_14_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_249 ),
	.cout(Xd_0__inst_mult_14_250 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_18_q ),
	.datab(!Xd_0__inst_mult_9_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_254 ),
	.cout(Xd_0__inst_mult_9_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_18_q ),
	.datab(!Xd_0__inst_mult_8_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_254 ),
	.cout(Xd_0__inst_mult_8_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_18_q ),
	.datab(!Xd_0__inst_mult_11_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_254 ),
	.cout(Xd_0__inst_mult_11_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_18_q ),
	.datab(!Xd_0__inst_mult_10_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_254 ),
	.cout(Xd_0__inst_mult_10_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_18_q ),
	.datab(!Xd_0__inst_mult_5_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_254 ),
	.cout(Xd_0__inst_mult_5_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_18_q ),
	.datab(!Xd_0__inst_mult_4_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_254 ),
	.cout(Xd_0__inst_mult_4_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_18_q ),
	.datab(!Xd_0__inst_mult_7_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_254 ),
	.cout(Xd_0__inst_mult_7_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_18_q ),
	.datab(!Xd_0__inst_mult_6_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_254 ),
	.cout(Xd_0__inst_mult_6_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_18_q ),
	.datab(!Xd_0__inst_mult_1_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_254 ),
	.cout(Xd_0__inst_mult_1_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_18_q ),
	.datab(!Xd_0__inst_mult_0_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_254 ),
	.cout(Xd_0__inst_mult_0_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_18_q ),
	.datab(!Xd_0__inst_mult_3_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_254 ),
	.cout(Xd_0__inst_mult_3_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_18_q ),
	.datab(!Xd_0__inst_mult_2_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_304 ),
	.cout(Xd_0__inst_mult_2_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_20_q ),
	.datab(!Xd_0__inst_mult_29_21_q ),
	.datac(!Xd_0__inst_mult_29_22_q ),
	.datad(!Xd_0__inst_mult_29_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_279 ),
	.cout(Xd_0__inst_mult_29_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_20_q ),
	.datab(!Xd_0__inst_mult_28_21_q ),
	.datac(!Xd_0__inst_mult_28_22_q ),
	.datad(!Xd_0__inst_mult_28_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_259 ),
	.cout(Xd_0__inst_mult_28_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_20_q ),
	.datab(!Xd_0__inst_mult_31_21_q ),
	.datac(!Xd_0__inst_mult_31_22_q ),
	.datad(!Xd_0__inst_mult_31_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_259 ),
	.cout(Xd_0__inst_mult_31_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_20_q ),
	.datab(!Xd_0__inst_mult_30_21_q ),
	.datac(!Xd_0__inst_mult_30_22_q ),
	.datad(!Xd_0__inst_mult_30_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_259 ),
	.cout(Xd_0__inst_mult_30_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_20_q ),
	.datab(!Xd_0__inst_mult_25_21_q ),
	.datac(!Xd_0__inst_mult_25_22_q ),
	.datad(!Xd_0__inst_mult_25_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_339 ),
	.cout(Xd_0__inst_mult_25_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_20_q ),
	.datab(!Xd_0__inst_mult_24_21_q ),
	.datac(!Xd_0__inst_mult_24_22_q ),
	.datad(!Xd_0__inst_mult_24_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_479 ),
	.cout(Xd_0__inst_mult_24_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_20_q ),
	.datab(!Xd_0__inst_mult_27_21_q ),
	.datac(!Xd_0__inst_mult_27_22_q ),
	.datad(!Xd_0__inst_mult_27_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_339 ),
	.cout(Xd_0__inst_mult_27_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_20_q ),
	.datab(!Xd_0__inst_mult_26_21_q ),
	.datac(!Xd_0__inst_mult_26_22_q ),
	.datad(!Xd_0__inst_mult_26_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_479 ),
	.cout(Xd_0__inst_mult_26_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_20_q ),
	.datab(!Xd_0__inst_mult_21_21_q ),
	.datac(!Xd_0__inst_mult_21_22_q ),
	.datad(!Xd_0__inst_mult_21_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_279 ),
	.cout(Xd_0__inst_mult_21_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_20_q ),
	.datab(!Xd_0__inst_mult_20_21_q ),
	.datac(!Xd_0__inst_mult_20_22_q ),
	.datad(!Xd_0__inst_mult_20_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_279 ),
	.cout(Xd_0__inst_mult_20_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_20_q ),
	.datab(!Xd_0__inst_mult_23_21_q ),
	.datac(!Xd_0__inst_mult_23_22_q ),
	.datad(!Xd_0__inst_mult_23_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_279 ),
	.cout(Xd_0__inst_mult_23_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_20_q ),
	.datab(!Xd_0__inst_mult_22_21_q ),
	.datac(!Xd_0__inst_mult_22_22_q ),
	.datad(!Xd_0__inst_mult_22_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_279 ),
	.cout(Xd_0__inst_mult_22_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_20_q ),
	.datab(!Xd_0__inst_mult_17_21_q ),
	.datac(!Xd_0__inst_mult_17_22_q ),
	.datad(!Xd_0__inst_mult_17_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_279 ),
	.cout(Xd_0__inst_mult_17_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_20_q ),
	.datab(!Xd_0__inst_mult_16_21_q ),
	.datac(!Xd_0__inst_mult_16_22_q ),
	.datad(!Xd_0__inst_mult_16_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_279 ),
	.cout(Xd_0__inst_mult_16_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_20_q ),
	.datab(!Xd_0__inst_mult_19_21_q ),
	.datac(!Xd_0__inst_mult_19_22_q ),
	.datad(!Xd_0__inst_mult_19_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_279 ),
	.cout(Xd_0__inst_mult_19_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_20_q ),
	.datab(!Xd_0__inst_mult_18_21_q ),
	.datac(!Xd_0__inst_mult_18_22_q ),
	.datad(!Xd_0__inst_mult_18_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_254 ),
	.cout(Xd_0__inst_mult_18_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_20_q ),
	.datab(!Xd_0__inst_mult_13_21_q ),
	.datac(!Xd_0__inst_mult_13_22_q ),
	.datad(!Xd_0__inst_mult_13_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_259 ),
	.cout(Xd_0__inst_mult_13_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_20_q ),
	.datab(!Xd_0__inst_mult_12_21_q ),
	.datac(!Xd_0__inst_mult_12_22_q ),
	.datad(!Xd_0__inst_mult_12_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_254 ),
	.cout(Xd_0__inst_mult_12_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_20_q ),
	.datab(!Xd_0__inst_mult_15_21_q ),
	.datac(!Xd_0__inst_mult_15_22_q ),
	.datad(!Xd_0__inst_mult_15_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_254 ),
	.cout(Xd_0__inst_mult_15_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_92 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_20_q ),
	.datab(!Xd_0__inst_mult_14_21_q ),
	.datac(!Xd_0__inst_mult_14_22_q ),
	.datad(!Xd_0__inst_mult_14_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_250 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_254 ),
	.cout(Xd_0__inst_mult_14_255 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_20_q ),
	.datab(!Xd_0__inst_mult_9_21_q ),
	.datac(!Xd_0__inst_mult_9_22_q ),
	.datad(!Xd_0__inst_mult_9_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_259 ),
	.cout(Xd_0__inst_mult_9_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_20_q ),
	.datab(!Xd_0__inst_mult_8_21_q ),
	.datac(!Xd_0__inst_mult_8_22_q ),
	.datad(!Xd_0__inst_mult_8_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_259 ),
	.cout(Xd_0__inst_mult_8_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_20_q ),
	.datab(!Xd_0__inst_mult_11_21_q ),
	.datac(!Xd_0__inst_mult_11_22_q ),
	.datad(!Xd_0__inst_mult_11_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_259 ),
	.cout(Xd_0__inst_mult_11_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_20_q ),
	.datab(!Xd_0__inst_mult_10_21_q ),
	.datac(!Xd_0__inst_mult_10_22_q ),
	.datad(!Xd_0__inst_mult_10_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_259 ),
	.cout(Xd_0__inst_mult_10_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_20_q ),
	.datab(!Xd_0__inst_mult_5_21_q ),
	.datac(!Xd_0__inst_mult_5_22_q ),
	.datad(!Xd_0__inst_mult_5_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_259 ),
	.cout(Xd_0__inst_mult_5_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_20_q ),
	.datab(!Xd_0__inst_mult_4_21_q ),
	.datac(!Xd_0__inst_mult_4_22_q ),
	.datad(!Xd_0__inst_mult_4_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_259 ),
	.cout(Xd_0__inst_mult_4_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_20_q ),
	.datab(!Xd_0__inst_mult_7_21_q ),
	.datac(!Xd_0__inst_mult_7_22_q ),
	.datad(!Xd_0__inst_mult_7_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_259 ),
	.cout(Xd_0__inst_mult_7_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_20_q ),
	.datab(!Xd_0__inst_mult_6_21_q ),
	.datac(!Xd_0__inst_mult_6_22_q ),
	.datad(!Xd_0__inst_mult_6_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_259 ),
	.cout(Xd_0__inst_mult_6_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_20_q ),
	.datab(!Xd_0__inst_mult_1_21_q ),
	.datac(!Xd_0__inst_mult_1_22_q ),
	.datad(!Xd_0__inst_mult_1_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_259 ),
	.cout(Xd_0__inst_mult_1_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_20_q ),
	.datab(!Xd_0__inst_mult_0_21_q ),
	.datac(!Xd_0__inst_mult_0_22_q ),
	.datad(!Xd_0__inst_mult_0_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_259 ),
	.cout(Xd_0__inst_mult_0_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_20_q ),
	.datab(!Xd_0__inst_mult_3_21_q ),
	.datac(!Xd_0__inst_mult_3_22_q ),
	.datad(!Xd_0__inst_mult_3_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_259 ),
	.cout(Xd_0__inst_mult_3_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_20_q ),
	.datab(!Xd_0__inst_mult_2_21_q ),
	.datac(!Xd_0__inst_mult_2_22_q ),
	.datad(!Xd_0__inst_mult_2_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_309 ),
	.cout(Xd_0__inst_mult_2_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_24_q ),
	.datab(!Xd_0__inst_mult_29_25_q ),
	.datac(!Xd_0__inst_mult_29_20_q ),
	.datad(!Xd_0__inst_mult_29_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_284 ),
	.cout(Xd_0__inst_mult_29_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_24_q ),
	.datab(!Xd_0__inst_mult_28_25_q ),
	.datac(!Xd_0__inst_mult_28_20_q ),
	.datad(!Xd_0__inst_mult_28_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_264 ),
	.cout(Xd_0__inst_mult_28_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_24_q ),
	.datab(!Xd_0__inst_mult_31_25_q ),
	.datac(!Xd_0__inst_mult_31_20_q ),
	.datad(!Xd_0__inst_mult_31_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_264 ),
	.cout(Xd_0__inst_mult_31_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_24_q ),
	.datab(!Xd_0__inst_mult_30_25_q ),
	.datac(!Xd_0__inst_mult_30_20_q ),
	.datad(!Xd_0__inst_mult_30_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_264 ),
	.cout(Xd_0__inst_mult_30_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_24_q ),
	.datab(!Xd_0__inst_mult_25_25_q ),
	.datac(!Xd_0__inst_mult_25_20_q ),
	.datad(!Xd_0__inst_mult_25_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_344 ),
	.cout(Xd_0__inst_mult_25_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_24_q ),
	.datab(!Xd_0__inst_mult_24_25_q ),
	.datac(!Xd_0__inst_mult_24_20_q ),
	.datad(!Xd_0__inst_mult_24_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_484 ),
	.cout(Xd_0__inst_mult_24_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_24_q ),
	.datab(!Xd_0__inst_mult_27_25_q ),
	.datac(!Xd_0__inst_mult_27_20_q ),
	.datad(!Xd_0__inst_mult_27_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_344 ),
	.cout(Xd_0__inst_mult_27_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_24_q ),
	.datab(!Xd_0__inst_mult_26_25_q ),
	.datac(!Xd_0__inst_mult_26_20_q ),
	.datad(!Xd_0__inst_mult_26_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_484 ),
	.cout(Xd_0__inst_mult_26_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_24_q ),
	.datab(!Xd_0__inst_mult_21_25_q ),
	.datac(!Xd_0__inst_mult_21_20_q ),
	.datad(!Xd_0__inst_mult_21_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_284 ),
	.cout(Xd_0__inst_mult_21_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_24_q ),
	.datab(!Xd_0__inst_mult_20_25_q ),
	.datac(!Xd_0__inst_mult_20_20_q ),
	.datad(!Xd_0__inst_mult_20_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_284 ),
	.cout(Xd_0__inst_mult_20_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_24_q ),
	.datab(!Xd_0__inst_mult_23_25_q ),
	.datac(!Xd_0__inst_mult_23_20_q ),
	.datad(!Xd_0__inst_mult_23_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_284 ),
	.cout(Xd_0__inst_mult_23_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_24_q ),
	.datab(!Xd_0__inst_mult_22_25_q ),
	.datac(!Xd_0__inst_mult_22_20_q ),
	.datad(!Xd_0__inst_mult_22_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_284 ),
	.cout(Xd_0__inst_mult_22_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_24_q ),
	.datab(!Xd_0__inst_mult_17_25_q ),
	.datac(!Xd_0__inst_mult_17_20_q ),
	.datad(!Xd_0__inst_mult_17_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_284 ),
	.cout(Xd_0__inst_mult_17_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_24_q ),
	.datab(!Xd_0__inst_mult_16_25_q ),
	.datac(!Xd_0__inst_mult_16_20_q ),
	.datad(!Xd_0__inst_mult_16_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_284 ),
	.cout(Xd_0__inst_mult_16_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_24_q ),
	.datab(!Xd_0__inst_mult_19_25_q ),
	.datac(!Xd_0__inst_mult_19_20_q ),
	.datad(!Xd_0__inst_mult_19_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_284 ),
	.cout(Xd_0__inst_mult_19_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_24_q ),
	.datab(!Xd_0__inst_mult_18_25_q ),
	.datac(!Xd_0__inst_mult_18_20_q ),
	.datad(!Xd_0__inst_mult_18_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_259 ),
	.cout(Xd_0__inst_mult_18_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_24_q ),
	.datab(!Xd_0__inst_mult_13_25_q ),
	.datac(!Xd_0__inst_mult_13_20_q ),
	.datad(!Xd_0__inst_mult_13_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_264 ),
	.cout(Xd_0__inst_mult_13_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_24_q ),
	.datab(!Xd_0__inst_mult_12_25_q ),
	.datac(!Xd_0__inst_mult_12_20_q ),
	.datad(!Xd_0__inst_mult_12_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_259 ),
	.cout(Xd_0__inst_mult_12_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_24_q ),
	.datab(!Xd_0__inst_mult_15_25_q ),
	.datac(!Xd_0__inst_mult_15_20_q ),
	.datad(!Xd_0__inst_mult_15_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_259 ),
	.cout(Xd_0__inst_mult_15_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_93 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_24_q ),
	.datab(!Xd_0__inst_mult_14_25_q ),
	.datac(!Xd_0__inst_mult_14_20_q ),
	.datad(!Xd_0__inst_mult_14_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_255 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_259 ),
	.cout(Xd_0__inst_mult_14_260 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_24_q ),
	.datab(!Xd_0__inst_mult_9_25_q ),
	.datac(!Xd_0__inst_mult_9_20_q ),
	.datad(!Xd_0__inst_mult_9_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_264 ),
	.cout(Xd_0__inst_mult_9_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_24_q ),
	.datab(!Xd_0__inst_mult_8_25_q ),
	.datac(!Xd_0__inst_mult_8_20_q ),
	.datad(!Xd_0__inst_mult_8_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_264 ),
	.cout(Xd_0__inst_mult_8_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_24_q ),
	.datab(!Xd_0__inst_mult_11_25_q ),
	.datac(!Xd_0__inst_mult_11_20_q ),
	.datad(!Xd_0__inst_mult_11_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_264 ),
	.cout(Xd_0__inst_mult_11_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_24_q ),
	.datab(!Xd_0__inst_mult_10_25_q ),
	.datac(!Xd_0__inst_mult_10_20_q ),
	.datad(!Xd_0__inst_mult_10_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_264 ),
	.cout(Xd_0__inst_mult_10_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_24_q ),
	.datab(!Xd_0__inst_mult_5_25_q ),
	.datac(!Xd_0__inst_mult_5_20_q ),
	.datad(!Xd_0__inst_mult_5_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_264 ),
	.cout(Xd_0__inst_mult_5_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_24_q ),
	.datab(!Xd_0__inst_mult_4_25_q ),
	.datac(!Xd_0__inst_mult_4_20_q ),
	.datad(!Xd_0__inst_mult_4_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_264 ),
	.cout(Xd_0__inst_mult_4_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_24_q ),
	.datab(!Xd_0__inst_mult_7_25_q ),
	.datac(!Xd_0__inst_mult_7_20_q ),
	.datad(!Xd_0__inst_mult_7_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_264 ),
	.cout(Xd_0__inst_mult_7_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_24_q ),
	.datab(!Xd_0__inst_mult_6_25_q ),
	.datac(!Xd_0__inst_mult_6_20_q ),
	.datad(!Xd_0__inst_mult_6_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_264 ),
	.cout(Xd_0__inst_mult_6_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_24_q ),
	.datab(!Xd_0__inst_mult_1_25_q ),
	.datac(!Xd_0__inst_mult_1_20_q ),
	.datad(!Xd_0__inst_mult_1_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_264 ),
	.cout(Xd_0__inst_mult_1_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_24_q ),
	.datab(!Xd_0__inst_mult_0_25_q ),
	.datac(!Xd_0__inst_mult_0_20_q ),
	.datad(!Xd_0__inst_mult_0_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_264 ),
	.cout(Xd_0__inst_mult_0_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_24_q ),
	.datab(!Xd_0__inst_mult_3_25_q ),
	.datac(!Xd_0__inst_mult_3_20_q ),
	.datad(!Xd_0__inst_mult_3_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_264 ),
	.cout(Xd_0__inst_mult_3_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_24_q ),
	.datab(!Xd_0__inst_mult_2_25_q ),
	.datac(!Xd_0__inst_mult_2_20_q ),
	.datad(!Xd_0__inst_mult_2_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_314 ),
	.cout(Xd_0__inst_mult_2_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_26_q ),
	.datab(!Xd_0__inst_mult_29_27_q ),
	.datac(!Xd_0__inst_mult_29_24_q ),
	.datad(!Xd_0__inst_mult_29_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_289 ),
	.cout(Xd_0__inst_mult_29_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_26_q ),
	.datab(!Xd_0__inst_mult_28_27_q ),
	.datac(!Xd_0__inst_mult_28_24_q ),
	.datad(!Xd_0__inst_mult_28_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_269 ),
	.cout(Xd_0__inst_mult_28_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_26_q ),
	.datab(!Xd_0__inst_mult_31_27_q ),
	.datac(!Xd_0__inst_mult_31_24_q ),
	.datad(!Xd_0__inst_mult_31_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_269 ),
	.cout(Xd_0__inst_mult_31_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_26_q ),
	.datab(!Xd_0__inst_mult_30_27_q ),
	.datac(!Xd_0__inst_mult_30_24_q ),
	.datad(!Xd_0__inst_mult_30_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_269 ),
	.cout(Xd_0__inst_mult_30_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_26_q ),
	.datab(!Xd_0__inst_mult_25_27_q ),
	.datac(!Xd_0__inst_mult_25_24_q ),
	.datad(!Xd_0__inst_mult_25_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_349 ),
	.cout(Xd_0__inst_mult_25_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_26_q ),
	.datab(!Xd_0__inst_mult_24_27_q ),
	.datac(!Xd_0__inst_mult_24_24_q ),
	.datad(!Xd_0__inst_mult_24_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_489 ),
	.cout(Xd_0__inst_mult_24_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_26_q ),
	.datab(!Xd_0__inst_mult_27_27_q ),
	.datac(!Xd_0__inst_mult_27_24_q ),
	.datad(!Xd_0__inst_mult_27_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_349 ),
	.cout(Xd_0__inst_mult_27_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_26_q ),
	.datab(!Xd_0__inst_mult_26_27_q ),
	.datac(!Xd_0__inst_mult_26_24_q ),
	.datad(!Xd_0__inst_mult_26_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_489 ),
	.cout(Xd_0__inst_mult_26_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_26_q ),
	.datab(!Xd_0__inst_mult_21_27_q ),
	.datac(!Xd_0__inst_mult_21_24_q ),
	.datad(!Xd_0__inst_mult_21_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_289 ),
	.cout(Xd_0__inst_mult_21_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_26_q ),
	.datab(!Xd_0__inst_mult_20_27_q ),
	.datac(!Xd_0__inst_mult_20_24_q ),
	.datad(!Xd_0__inst_mult_20_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_289 ),
	.cout(Xd_0__inst_mult_20_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_26_q ),
	.datab(!Xd_0__inst_mult_23_27_q ),
	.datac(!Xd_0__inst_mult_23_24_q ),
	.datad(!Xd_0__inst_mult_23_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_289 ),
	.cout(Xd_0__inst_mult_23_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_26_q ),
	.datab(!Xd_0__inst_mult_22_27_q ),
	.datac(!Xd_0__inst_mult_22_24_q ),
	.datad(!Xd_0__inst_mult_22_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_289 ),
	.cout(Xd_0__inst_mult_22_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_26_q ),
	.datab(!Xd_0__inst_mult_17_27_q ),
	.datac(!Xd_0__inst_mult_17_24_q ),
	.datad(!Xd_0__inst_mult_17_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_289 ),
	.cout(Xd_0__inst_mult_17_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_26_q ),
	.datab(!Xd_0__inst_mult_16_27_q ),
	.datac(!Xd_0__inst_mult_16_24_q ),
	.datad(!Xd_0__inst_mult_16_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_289 ),
	.cout(Xd_0__inst_mult_16_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_26_q ),
	.datab(!Xd_0__inst_mult_19_27_q ),
	.datac(!Xd_0__inst_mult_19_24_q ),
	.datad(!Xd_0__inst_mult_19_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_289 ),
	.cout(Xd_0__inst_mult_19_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_26_q ),
	.datab(!Xd_0__inst_mult_18_27_q ),
	.datac(!Xd_0__inst_mult_18_24_q ),
	.datad(!Xd_0__inst_mult_18_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_264 ),
	.cout(Xd_0__inst_mult_18_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_26_q ),
	.datab(!Xd_0__inst_mult_13_27_q ),
	.datac(!Xd_0__inst_mult_13_24_q ),
	.datad(!Xd_0__inst_mult_13_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_269 ),
	.cout(Xd_0__inst_mult_13_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_26_q ),
	.datab(!Xd_0__inst_mult_12_27_q ),
	.datac(!Xd_0__inst_mult_12_24_q ),
	.datad(!Xd_0__inst_mult_12_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_264 ),
	.cout(Xd_0__inst_mult_12_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_26_q ),
	.datab(!Xd_0__inst_mult_15_27_q ),
	.datac(!Xd_0__inst_mult_15_24_q ),
	.datad(!Xd_0__inst_mult_15_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_264 ),
	.cout(Xd_0__inst_mult_15_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_94 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_26_q ),
	.datab(!Xd_0__inst_mult_14_27_q ),
	.datac(!Xd_0__inst_mult_14_24_q ),
	.datad(!Xd_0__inst_mult_14_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_260 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_264 ),
	.cout(Xd_0__inst_mult_14_265 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_26_q ),
	.datab(!Xd_0__inst_mult_9_27_q ),
	.datac(!Xd_0__inst_mult_9_24_q ),
	.datad(!Xd_0__inst_mult_9_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_269 ),
	.cout(Xd_0__inst_mult_9_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_26_q ),
	.datab(!Xd_0__inst_mult_8_27_q ),
	.datac(!Xd_0__inst_mult_8_24_q ),
	.datad(!Xd_0__inst_mult_8_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_269 ),
	.cout(Xd_0__inst_mult_8_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_26_q ),
	.datab(!Xd_0__inst_mult_11_27_q ),
	.datac(!Xd_0__inst_mult_11_24_q ),
	.datad(!Xd_0__inst_mult_11_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_269 ),
	.cout(Xd_0__inst_mult_11_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_26_q ),
	.datab(!Xd_0__inst_mult_10_27_q ),
	.datac(!Xd_0__inst_mult_10_24_q ),
	.datad(!Xd_0__inst_mult_10_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_269 ),
	.cout(Xd_0__inst_mult_10_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_26_q ),
	.datab(!Xd_0__inst_mult_5_27_q ),
	.datac(!Xd_0__inst_mult_5_24_q ),
	.datad(!Xd_0__inst_mult_5_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_269 ),
	.cout(Xd_0__inst_mult_5_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_26_q ),
	.datab(!Xd_0__inst_mult_4_27_q ),
	.datac(!Xd_0__inst_mult_4_24_q ),
	.datad(!Xd_0__inst_mult_4_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_269 ),
	.cout(Xd_0__inst_mult_4_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_26_q ),
	.datab(!Xd_0__inst_mult_7_27_q ),
	.datac(!Xd_0__inst_mult_7_24_q ),
	.datad(!Xd_0__inst_mult_7_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_269 ),
	.cout(Xd_0__inst_mult_7_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_26_q ),
	.datab(!Xd_0__inst_mult_6_27_q ),
	.datac(!Xd_0__inst_mult_6_24_q ),
	.datad(!Xd_0__inst_mult_6_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_269 ),
	.cout(Xd_0__inst_mult_6_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_26_q ),
	.datab(!Xd_0__inst_mult_1_27_q ),
	.datac(!Xd_0__inst_mult_1_24_q ),
	.datad(!Xd_0__inst_mult_1_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_269 ),
	.cout(Xd_0__inst_mult_1_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_26_q ),
	.datab(!Xd_0__inst_mult_0_27_q ),
	.datac(!Xd_0__inst_mult_0_24_q ),
	.datad(!Xd_0__inst_mult_0_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_269 ),
	.cout(Xd_0__inst_mult_0_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_26_q ),
	.datab(!Xd_0__inst_mult_3_27_q ),
	.datac(!Xd_0__inst_mult_3_24_q ),
	.datad(!Xd_0__inst_mult_3_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_269 ),
	.cout(Xd_0__inst_mult_3_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_26_q ),
	.datab(!Xd_0__inst_mult_2_27_q ),
	.datac(!Xd_0__inst_mult_2_24_q ),
	.datad(!Xd_0__inst_mult_2_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_319 ),
	.cout(Xd_0__inst_mult_2_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_28_q ),
	.datab(!Xd_0__inst_mult_29_29_q ),
	.datac(!Xd_0__inst_mult_29_26_q ),
	.datad(!Xd_0__inst_mult_29_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_294 ),
	.cout(Xd_0__inst_mult_29_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_28_q ),
	.datab(!Xd_0__inst_mult_28_29_q ),
	.datac(!Xd_0__inst_mult_28_26_q ),
	.datad(!Xd_0__inst_mult_28_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_274 ),
	.cout(Xd_0__inst_mult_28_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_28_q ),
	.datab(!Xd_0__inst_mult_31_29_q ),
	.datac(!Xd_0__inst_mult_31_26_q ),
	.datad(!Xd_0__inst_mult_31_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_274 ),
	.cout(Xd_0__inst_mult_31_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_28_q ),
	.datab(!Xd_0__inst_mult_30_29_q ),
	.datac(!Xd_0__inst_mult_30_26_q ),
	.datad(!Xd_0__inst_mult_30_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_274 ),
	.cout(Xd_0__inst_mult_30_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_112 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_28_q ),
	.datab(!Xd_0__inst_mult_25_29_q ),
	.datac(!Xd_0__inst_mult_25_26_q ),
	.datad(!Xd_0__inst_mult_25_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_354 ),
	.cout(Xd_0__inst_mult_25_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_28_q ),
	.datab(!Xd_0__inst_mult_24_29_q ),
	.datac(!Xd_0__inst_mult_24_26_q ),
	.datad(!Xd_0__inst_mult_24_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_494 ),
	.cout(Xd_0__inst_mult_24_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_112 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_28_q ),
	.datab(!Xd_0__inst_mult_27_29_q ),
	.datac(!Xd_0__inst_mult_27_26_q ),
	.datad(!Xd_0__inst_mult_27_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_354 ),
	.cout(Xd_0__inst_mult_27_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_28_q ),
	.datab(!Xd_0__inst_mult_26_29_q ),
	.datac(!Xd_0__inst_mult_26_26_q ),
	.datad(!Xd_0__inst_mult_26_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_494 ),
	.cout(Xd_0__inst_mult_26_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_28_q ),
	.datab(!Xd_0__inst_mult_21_29_q ),
	.datac(!Xd_0__inst_mult_21_26_q ),
	.datad(!Xd_0__inst_mult_21_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_294 ),
	.cout(Xd_0__inst_mult_21_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_28_q ),
	.datab(!Xd_0__inst_mult_20_29_q ),
	.datac(!Xd_0__inst_mult_20_26_q ),
	.datad(!Xd_0__inst_mult_20_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_294 ),
	.cout(Xd_0__inst_mult_20_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_28_q ),
	.datab(!Xd_0__inst_mult_23_29_q ),
	.datac(!Xd_0__inst_mult_23_26_q ),
	.datad(!Xd_0__inst_mult_23_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_294 ),
	.cout(Xd_0__inst_mult_23_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_28_q ),
	.datab(!Xd_0__inst_mult_22_29_q ),
	.datac(!Xd_0__inst_mult_22_26_q ),
	.datad(!Xd_0__inst_mult_22_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_294 ),
	.cout(Xd_0__inst_mult_22_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_28_q ),
	.datab(!Xd_0__inst_mult_17_29_q ),
	.datac(!Xd_0__inst_mult_17_26_q ),
	.datad(!Xd_0__inst_mult_17_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_294 ),
	.cout(Xd_0__inst_mult_17_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_28_q ),
	.datab(!Xd_0__inst_mult_16_29_q ),
	.datac(!Xd_0__inst_mult_16_26_q ),
	.datad(!Xd_0__inst_mult_16_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_294 ),
	.cout(Xd_0__inst_mult_16_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_28_q ),
	.datab(!Xd_0__inst_mult_19_29_q ),
	.datac(!Xd_0__inst_mult_19_26_q ),
	.datad(!Xd_0__inst_mult_19_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_294 ),
	.cout(Xd_0__inst_mult_19_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_28_q ),
	.datab(!Xd_0__inst_mult_18_29_q ),
	.datac(!Xd_0__inst_mult_18_26_q ),
	.datad(!Xd_0__inst_mult_18_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_269 ),
	.cout(Xd_0__inst_mult_18_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_28_q ),
	.datab(!Xd_0__inst_mult_13_29_q ),
	.datac(!Xd_0__inst_mult_13_26_q ),
	.datad(!Xd_0__inst_mult_13_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_274 ),
	.cout(Xd_0__inst_mult_13_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_28_q ),
	.datab(!Xd_0__inst_mult_12_29_q ),
	.datac(!Xd_0__inst_mult_12_26_q ),
	.datad(!Xd_0__inst_mult_12_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_269 ),
	.cout(Xd_0__inst_mult_12_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_28_q ),
	.datab(!Xd_0__inst_mult_15_29_q ),
	.datac(!Xd_0__inst_mult_15_26_q ),
	.datad(!Xd_0__inst_mult_15_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_269 ),
	.cout(Xd_0__inst_mult_15_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_95 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_28_q ),
	.datab(!Xd_0__inst_mult_14_29_q ),
	.datac(!Xd_0__inst_mult_14_26_q ),
	.datad(!Xd_0__inst_mult_14_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_265 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_269 ),
	.cout(Xd_0__inst_mult_14_270 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_28_q ),
	.datab(!Xd_0__inst_mult_9_29_q ),
	.datac(!Xd_0__inst_mult_9_26_q ),
	.datad(!Xd_0__inst_mult_9_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_274 ),
	.cout(Xd_0__inst_mult_9_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_28_q ),
	.datab(!Xd_0__inst_mult_8_29_q ),
	.datac(!Xd_0__inst_mult_8_26_q ),
	.datad(!Xd_0__inst_mult_8_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_274 ),
	.cout(Xd_0__inst_mult_8_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_28_q ),
	.datab(!Xd_0__inst_mult_11_29_q ),
	.datac(!Xd_0__inst_mult_11_26_q ),
	.datad(!Xd_0__inst_mult_11_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_274 ),
	.cout(Xd_0__inst_mult_11_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_28_q ),
	.datab(!Xd_0__inst_mult_10_29_q ),
	.datac(!Xd_0__inst_mult_10_26_q ),
	.datad(!Xd_0__inst_mult_10_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_274 ),
	.cout(Xd_0__inst_mult_10_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_28_q ),
	.datab(!Xd_0__inst_mult_5_29_q ),
	.datac(!Xd_0__inst_mult_5_26_q ),
	.datad(!Xd_0__inst_mult_5_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_274 ),
	.cout(Xd_0__inst_mult_5_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_28_q ),
	.datab(!Xd_0__inst_mult_4_29_q ),
	.datac(!Xd_0__inst_mult_4_26_q ),
	.datad(!Xd_0__inst_mult_4_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_274 ),
	.cout(Xd_0__inst_mult_4_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_28_q ),
	.datab(!Xd_0__inst_mult_7_29_q ),
	.datac(!Xd_0__inst_mult_7_26_q ),
	.datad(!Xd_0__inst_mult_7_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_274 ),
	.cout(Xd_0__inst_mult_7_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_28_q ),
	.datab(!Xd_0__inst_mult_6_29_q ),
	.datac(!Xd_0__inst_mult_6_26_q ),
	.datad(!Xd_0__inst_mult_6_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_274 ),
	.cout(Xd_0__inst_mult_6_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_28_q ),
	.datab(!Xd_0__inst_mult_1_29_q ),
	.datac(!Xd_0__inst_mult_1_26_q ),
	.datad(!Xd_0__inst_mult_1_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_274 ),
	.cout(Xd_0__inst_mult_1_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_28_q ),
	.datab(!Xd_0__inst_mult_0_29_q ),
	.datac(!Xd_0__inst_mult_0_26_q ),
	.datad(!Xd_0__inst_mult_0_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_274 ),
	.cout(Xd_0__inst_mult_0_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_28_q ),
	.datab(!Xd_0__inst_mult_3_29_q ),
	.datac(!Xd_0__inst_mult_3_26_q ),
	.datad(!Xd_0__inst_mult_3_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_274 ),
	.cout(Xd_0__inst_mult_3_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_106 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_28_q ),
	.datab(!Xd_0__inst_mult_2_29_q ),
	.datac(!Xd_0__inst_mult_2_26_q ),
	.datad(!Xd_0__inst_mult_2_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_324 ),
	.cout(Xd_0__inst_mult_2_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_30_q ),
	.datab(!Xd_0__inst_mult_29_31_q ),
	.datac(!Xd_0__inst_mult_29_28_q ),
	.datad(!Xd_0__inst_mult_29_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_299 ),
	.cout(Xd_0__inst_mult_29_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_30_q ),
	.datab(!Xd_0__inst_mult_28_31_q ),
	.datac(!Xd_0__inst_mult_28_28_q ),
	.datad(!Xd_0__inst_mult_28_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_279 ),
	.cout(Xd_0__inst_mult_28_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_30_q ),
	.datab(!Xd_0__inst_mult_31_31_q ),
	.datac(!Xd_0__inst_mult_31_28_q ),
	.datad(!Xd_0__inst_mult_31_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_279 ),
	.cout(Xd_0__inst_mult_31_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_30_q ),
	.datab(!Xd_0__inst_mult_30_31_q ),
	.datac(!Xd_0__inst_mult_30_28_q ),
	.datad(!Xd_0__inst_mult_30_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_279 ),
	.cout(Xd_0__inst_mult_30_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_30_q ),
	.datab(!Xd_0__inst_mult_25_31_q ),
	.datac(!Xd_0__inst_mult_25_28_q ),
	.datad(!Xd_0__inst_mult_25_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_359 ),
	.cout(Xd_0__inst_mult_25_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_30_q ),
	.datab(!Xd_0__inst_mult_24_31_q ),
	.datac(!Xd_0__inst_mult_24_28_q ),
	.datad(!Xd_0__inst_mult_24_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_499 ),
	.cout(Xd_0__inst_mult_24_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_30_q ),
	.datab(!Xd_0__inst_mult_27_31_q ),
	.datac(!Xd_0__inst_mult_27_28_q ),
	.datad(!Xd_0__inst_mult_27_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_359 ),
	.cout(Xd_0__inst_mult_27_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_30_q ),
	.datab(!Xd_0__inst_mult_26_31_q ),
	.datac(!Xd_0__inst_mult_26_28_q ),
	.datad(!Xd_0__inst_mult_26_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_499 ),
	.cout(Xd_0__inst_mult_26_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_30_q ),
	.datab(!Xd_0__inst_mult_21_31_q ),
	.datac(!Xd_0__inst_mult_21_28_q ),
	.datad(!Xd_0__inst_mult_21_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_299 ),
	.cout(Xd_0__inst_mult_21_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_30_q ),
	.datab(!Xd_0__inst_mult_20_31_q ),
	.datac(!Xd_0__inst_mult_20_28_q ),
	.datad(!Xd_0__inst_mult_20_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_299 ),
	.cout(Xd_0__inst_mult_20_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_30_q ),
	.datab(!Xd_0__inst_mult_23_31_q ),
	.datac(!Xd_0__inst_mult_23_28_q ),
	.datad(!Xd_0__inst_mult_23_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_299 ),
	.cout(Xd_0__inst_mult_23_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_30_q ),
	.datab(!Xd_0__inst_mult_22_31_q ),
	.datac(!Xd_0__inst_mult_22_28_q ),
	.datad(!Xd_0__inst_mult_22_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_299 ),
	.cout(Xd_0__inst_mult_22_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_30_q ),
	.datab(!Xd_0__inst_mult_17_31_q ),
	.datac(!Xd_0__inst_mult_17_28_q ),
	.datad(!Xd_0__inst_mult_17_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_299 ),
	.cout(Xd_0__inst_mult_17_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_30_q ),
	.datab(!Xd_0__inst_mult_16_31_q ),
	.datac(!Xd_0__inst_mult_16_28_q ),
	.datad(!Xd_0__inst_mult_16_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_299 ),
	.cout(Xd_0__inst_mult_16_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_30_q ),
	.datab(!Xd_0__inst_mult_19_31_q ),
	.datac(!Xd_0__inst_mult_19_28_q ),
	.datad(!Xd_0__inst_mult_19_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_299 ),
	.cout(Xd_0__inst_mult_19_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_30_q ),
	.datab(!Xd_0__inst_mult_18_31_q ),
	.datac(!Xd_0__inst_mult_18_28_q ),
	.datad(!Xd_0__inst_mult_18_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_274 ),
	.cout(Xd_0__inst_mult_18_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_30_q ),
	.datab(!Xd_0__inst_mult_13_31_q ),
	.datac(!Xd_0__inst_mult_13_28_q ),
	.datad(!Xd_0__inst_mult_13_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_279 ),
	.cout(Xd_0__inst_mult_13_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_30_q ),
	.datab(!Xd_0__inst_mult_12_31_q ),
	.datac(!Xd_0__inst_mult_12_28_q ),
	.datad(!Xd_0__inst_mult_12_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_274 ),
	.cout(Xd_0__inst_mult_12_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_30_q ),
	.datab(!Xd_0__inst_mult_15_31_q ),
	.datac(!Xd_0__inst_mult_15_28_q ),
	.datad(!Xd_0__inst_mult_15_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_274 ),
	.cout(Xd_0__inst_mult_15_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_96 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_30_q ),
	.datab(!Xd_0__inst_mult_14_31_q ),
	.datac(!Xd_0__inst_mult_14_28_q ),
	.datad(!Xd_0__inst_mult_14_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_270 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_274 ),
	.cout(Xd_0__inst_mult_14_275 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_30_q ),
	.datab(!Xd_0__inst_mult_9_31_q ),
	.datac(!Xd_0__inst_mult_9_28_q ),
	.datad(!Xd_0__inst_mult_9_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_279 ),
	.cout(Xd_0__inst_mult_9_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_30_q ),
	.datab(!Xd_0__inst_mult_8_31_q ),
	.datac(!Xd_0__inst_mult_8_28_q ),
	.datad(!Xd_0__inst_mult_8_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_279 ),
	.cout(Xd_0__inst_mult_8_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_30_q ),
	.datab(!Xd_0__inst_mult_11_31_q ),
	.datac(!Xd_0__inst_mult_11_28_q ),
	.datad(!Xd_0__inst_mult_11_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_279 ),
	.cout(Xd_0__inst_mult_11_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_30_q ),
	.datab(!Xd_0__inst_mult_10_31_q ),
	.datac(!Xd_0__inst_mult_10_28_q ),
	.datad(!Xd_0__inst_mult_10_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_279 ),
	.cout(Xd_0__inst_mult_10_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_30_q ),
	.datab(!Xd_0__inst_mult_5_31_q ),
	.datac(!Xd_0__inst_mult_5_28_q ),
	.datad(!Xd_0__inst_mult_5_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_279 ),
	.cout(Xd_0__inst_mult_5_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_30_q ),
	.datab(!Xd_0__inst_mult_4_31_q ),
	.datac(!Xd_0__inst_mult_4_28_q ),
	.datad(!Xd_0__inst_mult_4_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_279 ),
	.cout(Xd_0__inst_mult_4_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_30_q ),
	.datab(!Xd_0__inst_mult_7_31_q ),
	.datac(!Xd_0__inst_mult_7_28_q ),
	.datad(!Xd_0__inst_mult_7_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_279 ),
	.cout(Xd_0__inst_mult_7_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_30_q ),
	.datab(!Xd_0__inst_mult_6_31_q ),
	.datac(!Xd_0__inst_mult_6_28_q ),
	.datad(!Xd_0__inst_mult_6_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_279 ),
	.cout(Xd_0__inst_mult_6_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_30_q ),
	.datab(!Xd_0__inst_mult_1_31_q ),
	.datac(!Xd_0__inst_mult_1_28_q ),
	.datad(!Xd_0__inst_mult_1_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_279 ),
	.cout(Xd_0__inst_mult_1_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_30_q ),
	.datab(!Xd_0__inst_mult_0_31_q ),
	.datac(!Xd_0__inst_mult_0_28_q ),
	.datad(!Xd_0__inst_mult_0_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_279 ),
	.cout(Xd_0__inst_mult_0_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_30_q ),
	.datab(!Xd_0__inst_mult_3_31_q ),
	.datac(!Xd_0__inst_mult_3_28_q ),
	.datad(!Xd_0__inst_mult_3_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_279 ),
	.cout(Xd_0__inst_mult_3_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_30_q ),
	.datab(!Xd_0__inst_mult_2_31_q ),
	.datac(!Xd_0__inst_mult_2_28_q ),
	.datad(!Xd_0__inst_mult_2_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_329 ),
	.cout(Xd_0__inst_mult_2_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_32_q ),
	.datab(!Xd_0__inst_mult_29_33_q ),
	.datac(!Xd_0__inst_mult_29_30_q ),
	.datad(!Xd_0__inst_mult_29_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_304 ),
	.cout(Xd_0__inst_mult_29_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_32_q ),
	.datab(!Xd_0__inst_mult_28_33_q ),
	.datac(!Xd_0__inst_mult_28_30_q ),
	.datad(!Xd_0__inst_mult_28_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_284 ),
	.cout(Xd_0__inst_mult_28_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_32_q ),
	.datab(!Xd_0__inst_mult_31_33_q ),
	.datac(!Xd_0__inst_mult_31_30_q ),
	.datad(!Xd_0__inst_mult_31_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_284 ),
	.cout(Xd_0__inst_mult_31_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_32_q ),
	.datab(!Xd_0__inst_mult_30_33_q ),
	.datac(!Xd_0__inst_mult_30_30_q ),
	.datad(!Xd_0__inst_mult_30_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_284 ),
	.cout(Xd_0__inst_mult_30_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_32_q ),
	.datab(!Xd_0__inst_mult_25_33_q ),
	.datac(!Xd_0__inst_mult_25_30_q ),
	.datad(!Xd_0__inst_mult_25_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_364 ),
	.cout(Xd_0__inst_mult_25_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_24_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_32_q ),
	.datab(!Xd_0__inst_mult_24_33_q ),
	.datac(!Xd_0__inst_mult_24_30_q ),
	.datad(!Xd_0__inst_mult_24_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_504 ),
	.cout(Xd_0__inst_mult_24_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_32_q ),
	.datab(!Xd_0__inst_mult_27_33_q ),
	.datac(!Xd_0__inst_mult_27_30_q ),
	.datad(!Xd_0__inst_mult_27_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_364 ),
	.cout(Xd_0__inst_mult_27_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_26_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_32_q ),
	.datab(!Xd_0__inst_mult_26_33_q ),
	.datac(!Xd_0__inst_mult_26_30_q ),
	.datad(!Xd_0__inst_mult_26_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_504 ),
	.cout(Xd_0__inst_mult_26_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_32_q ),
	.datab(!Xd_0__inst_mult_21_33_q ),
	.datac(!Xd_0__inst_mult_21_30_q ),
	.datad(!Xd_0__inst_mult_21_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_304 ),
	.cout(Xd_0__inst_mult_21_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_32_q ),
	.datab(!Xd_0__inst_mult_20_33_q ),
	.datac(!Xd_0__inst_mult_20_30_q ),
	.datad(!Xd_0__inst_mult_20_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_304 ),
	.cout(Xd_0__inst_mult_20_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_32_q ),
	.datab(!Xd_0__inst_mult_23_33_q ),
	.datac(!Xd_0__inst_mult_23_30_q ),
	.datad(!Xd_0__inst_mult_23_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_304 ),
	.cout(Xd_0__inst_mult_23_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_32_q ),
	.datab(!Xd_0__inst_mult_22_33_q ),
	.datac(!Xd_0__inst_mult_22_30_q ),
	.datad(!Xd_0__inst_mult_22_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_304 ),
	.cout(Xd_0__inst_mult_22_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_32_q ),
	.datab(!Xd_0__inst_mult_17_33_q ),
	.datac(!Xd_0__inst_mult_17_30_q ),
	.datad(!Xd_0__inst_mult_17_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_304 ),
	.cout(Xd_0__inst_mult_17_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_32_q ),
	.datab(!Xd_0__inst_mult_16_33_q ),
	.datac(!Xd_0__inst_mult_16_30_q ),
	.datad(!Xd_0__inst_mult_16_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_304 ),
	.cout(Xd_0__inst_mult_16_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_32_q ),
	.datab(!Xd_0__inst_mult_19_33_q ),
	.datac(!Xd_0__inst_mult_19_30_q ),
	.datad(!Xd_0__inst_mult_19_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_304 ),
	.cout(Xd_0__inst_mult_19_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_32_q ),
	.datab(!Xd_0__inst_mult_18_33_q ),
	.datac(!Xd_0__inst_mult_18_30_q ),
	.datad(!Xd_0__inst_mult_18_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_279 ),
	.cout(Xd_0__inst_mult_18_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_32_q ),
	.datab(!Xd_0__inst_mult_13_33_q ),
	.datac(!Xd_0__inst_mult_13_30_q ),
	.datad(!Xd_0__inst_mult_13_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_284 ),
	.cout(Xd_0__inst_mult_13_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_32_q ),
	.datab(!Xd_0__inst_mult_12_33_q ),
	.datac(!Xd_0__inst_mult_12_30_q ),
	.datad(!Xd_0__inst_mult_12_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_279 ),
	.cout(Xd_0__inst_mult_12_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_32_q ),
	.datab(!Xd_0__inst_mult_15_33_q ),
	.datac(!Xd_0__inst_mult_15_30_q ),
	.datad(!Xd_0__inst_mult_15_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_279 ),
	.cout(Xd_0__inst_mult_15_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_97 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_32_q ),
	.datab(!Xd_0__inst_mult_14_33_q ),
	.datac(!Xd_0__inst_mult_14_30_q ),
	.datad(!Xd_0__inst_mult_14_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_275 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_279 ),
	.cout(Xd_0__inst_mult_14_280 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_32_q ),
	.datab(!Xd_0__inst_mult_9_33_q ),
	.datac(!Xd_0__inst_mult_9_30_q ),
	.datad(!Xd_0__inst_mult_9_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_284 ),
	.cout(Xd_0__inst_mult_9_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_32_q ),
	.datab(!Xd_0__inst_mult_8_33_q ),
	.datac(!Xd_0__inst_mult_8_30_q ),
	.datad(!Xd_0__inst_mult_8_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_284 ),
	.cout(Xd_0__inst_mult_8_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_32_q ),
	.datab(!Xd_0__inst_mult_11_33_q ),
	.datac(!Xd_0__inst_mult_11_30_q ),
	.datad(!Xd_0__inst_mult_11_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_284 ),
	.cout(Xd_0__inst_mult_11_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_32_q ),
	.datab(!Xd_0__inst_mult_10_33_q ),
	.datac(!Xd_0__inst_mult_10_30_q ),
	.datad(!Xd_0__inst_mult_10_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_284 ),
	.cout(Xd_0__inst_mult_10_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(!Xd_0__inst_mult_5_30_q ),
	.datad(!Xd_0__inst_mult_5_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_284 ),
	.cout(Xd_0__inst_mult_5_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(!Xd_0__inst_mult_4_30_q ),
	.datad(!Xd_0__inst_mult_4_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_284 ),
	.cout(Xd_0__inst_mult_4_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(!Xd_0__inst_mult_7_30_q ),
	.datad(!Xd_0__inst_mult_7_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_284 ),
	.cout(Xd_0__inst_mult_7_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(!Xd_0__inst_mult_6_30_q ),
	.datad(!Xd_0__inst_mult_6_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_284 ),
	.cout(Xd_0__inst_mult_6_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(!Xd_0__inst_mult_1_30_q ),
	.datad(!Xd_0__inst_mult_1_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_284 ),
	.cout(Xd_0__inst_mult_1_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(!Xd_0__inst_mult_0_30_q ),
	.datad(!Xd_0__inst_mult_0_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_284 ),
	.cout(Xd_0__inst_mult_0_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(!Xd_0__inst_mult_3_30_q ),
	.datad(!Xd_0__inst_mult_3_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_284 ),
	.cout(Xd_0__inst_mult_3_285 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_108 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(!Xd_0__inst_mult_2_30_q ),
	.datad(!Xd_0__inst_mult_2_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_334 ),
	.cout(Xd_0__inst_mult_2_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_32_q ),
	.datab(!Xd_0__inst_mult_29_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_32_q ),
	.datab(!Xd_0__inst_mult_28_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_32_q ),
	.datab(!Xd_0__inst_mult_31_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_32_q ),
	.datab(!Xd_0__inst_mult_30_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_32_q ),
	.datab(!Xd_0__inst_mult_25_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_369 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_32_q ),
	.datab(!Xd_0__inst_mult_24_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_32_q ),
	.datab(!Xd_0__inst_mult_27_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_369 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_32_q ),
	.datab(!Xd_0__inst_mult_26_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_32_q ),
	.datab(!Xd_0__inst_mult_21_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_32_q ),
	.datab(!Xd_0__inst_mult_20_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_32_q ),
	.datab(!Xd_0__inst_mult_23_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_32_q ),
	.datab(!Xd_0__inst_mult_22_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_32_q ),
	.datab(!Xd_0__inst_mult_17_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_32_q ),
	.datab(!Xd_0__inst_mult_16_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_32_q ),
	.datab(!Xd_0__inst_mult_19_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_309 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_32_q ),
	.datab(!Xd_0__inst_mult_18_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_284 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_32_q ),
	.datab(!Xd_0__inst_mult_13_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_32_q ),
	.datab(!Xd_0__inst_mult_12_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_284 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_32_q ),
	.datab(!Xd_0__inst_mult_15_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_284 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_98 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_32_q ),
	.datab(!Xd_0__inst_mult_14_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_280 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_284 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_32_q ),
	.datab(!Xd_0__inst_mult_9_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_32_q ),
	.datab(!Xd_0__inst_mult_8_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_32_q ),
	.datab(!Xd_0__inst_mult_11_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_32_q ),
	.datab(!Xd_0__inst_mult_10_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_99 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_285 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_289 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_339 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_41 (
// Equation(s):

	.dataa(!din_a[371]),
	.datab(!din_b[371]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_41_sumout ),
	.cout(Xd_0__inst_i29_42 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_35 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[372]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_35_sumout ),
	.cout(Xd_0__inst_mult_31_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_40 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[360]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_40_sumout ),
	.cout(Xd_0__inst_mult_30_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_35 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[112]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_35_sumout ),
	.cout(Xd_0__inst_mult_9_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_294 ),
	.datab(!Xd_0__inst_mult_9_35_sumout ),
	.datac(!Xd_0__inst_mult_9_324 ),
	.datad(!Xd_0__inst_mult_9_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_299 ),
	.cout(Xd_0__inst_mult_9_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_46 (
// Equation(s):

	.dataa(!din_a[347]),
	.datab(!din_b[347]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_107 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_46_sumout ),
	.cout(Xd_0__inst_i29_47 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_51 (
// Equation(s):

	.dataa(!din_a[359]),
	.datab(!din_b[359]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_57 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_51_sumout ),
	.cout(Xd_0__inst_i29_52 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_45 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[348]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_45_sumout ),
	.cout(Xd_0__inst_mult_29_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_35 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[336]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_35_sumout ),
	.cout(Xd_0__inst_mult_28_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_35 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[100]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_35_sumout ),
	.cout(Xd_0__inst_mult_8_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_294 ),
	.datab(!Xd_0__inst_mult_8_35_sumout ),
	.datac(!Xd_0__inst_mult_8_324 ),
	.datad(!Xd_0__inst_mult_8_60_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_299 ),
	.cout(Xd_0__inst_mult_8_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_105 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[255]),
	.datac(!Xd_0__inst_mult_21_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_319 ),
	.cout(Xd_0__inst_mult_21_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_324 ),
	.datab(!Xd_0__inst_mult_21_319 ),
	.datac(!din_a[262]),
	.datad(!din_b[254]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_329 ),
	.cout(Xd_0__inst_mult_21_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_56 (
// Equation(s):

	.dataa(!din_a[323]),
	.datab(!din_b[323]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_62 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_56_sumout ),
	.cout(Xd_0__inst_i29_57 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_55 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[324]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_55_sumout ),
	.cout(Xd_0__inst_mult_27_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_55 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[312]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_55_sumout ),
	.cout(Xd_0__inst_mult_26_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_35 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[136]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_35_sumout ),
	.cout(Xd_0__inst_mult_11_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_294 ),
	.datab(!Xd_0__inst_mult_11_35_sumout ),
	.datac(!Xd_0__inst_mult_11_324 ),
	.datad(!Xd_0__inst_mult_11_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_299 ),
	.cout(Xd_0__inst_mult_11_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_61 (
// Equation(s):

	.dataa(!din_a[299]),
	.datab(!din_b[299]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_67 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_61_sumout ),
	.cout(Xd_0__inst_i29_62 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_66 (
// Equation(s):

	.dataa(!din_a[311]),
	.datab(!din_b[311]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_72 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_66_sumout ),
	.cout(Xd_0__inst_i29_67 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_50 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[300]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_50_sumout ),
	.cout(Xd_0__inst_mult_25_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_55 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[288]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_55_sumout ),
	.cout(Xd_0__inst_mult_24_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_35 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[124]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_35_sumout ),
	.cout(Xd_0__inst_mult_10_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_294 ),
	.datab(!Xd_0__inst_mult_10_35_sumout ),
	.datac(!Xd_0__inst_mult_10_324 ),
	.datad(!Xd_0__inst_mult_10_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_299 ),
	.cout(Xd_0__inst_mult_10_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_105 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[243]),
	.datac(!Xd_0__inst_mult_20_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_319 ),
	.cout(Xd_0__inst_mult_20_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_35 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[177]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_35_sumout ),
	.cout(Xd_0__inst_mult_14_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_324 ),
	.datab(!Xd_0__inst_mult_20_319 ),
	.datac(!din_a[250]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_329 ),
	.cout(Xd_0__inst_mult_20_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_116 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[303]),
	.datac(!din_a[306]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_374 ),
	.cout(Xd_0__inst_mult_25_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_117 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_414 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_379 ),
	.cout(Xd_0__inst_mult_25_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_118 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[301]),
	.datac(!din_a[309]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_384 ),
	.cout(Xd_0__inst_mult_25_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_384 ),
	.datab(!Xd_0__inst_mult_25_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_389 ),
	.cout(Xd_0__inst_mult_25_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_71 (
// Equation(s):

	.dataa(!din_a[275]),
	.datab(!din_b[275]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_77 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_71_sumout ),
	.cout(Xd_0__inst_i29_72 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_45 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[276]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_45_sumout ),
	.cout(Xd_0__inst_mult_23_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_45 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[264]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_45_sumout ),
	.cout(Xd_0__inst_mult_22_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_35 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[40]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_35_sumout ),
	.cout(Xd_0__inst_mult_3_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_294 ),
	.datab(!Xd_0__inst_mult_3_35_sumout ),
	.datac(!Xd_0__inst_mult_3_324 ),
	.datad(!Xd_0__inst_mult_3_55_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_299 ),
	.cout(Xd_0__inst_mult_3_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_76 (
// Equation(s):

	.dataa(!din_a[251]),
	.datab(!din_b[251]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_76_sumout ),
	.cout(Xd_0__inst_i29_77 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_81 (
// Equation(s):

	.dataa(!din_a[263]),
	.datab(!din_b[263]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_87 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_81_sumout ),
	.cout(Xd_0__inst_i29_82 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_45 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[252]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_45_sumout ),
	.cout(Xd_0__inst_mult_21_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_50 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[240]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_50_sumout ),
	.cout(Xd_0__inst_mult_20_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_35 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_35_sumout ),
	.cout(Xd_0__inst_mult_0_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_294 ),
	.datab(!Xd_0__inst_mult_0_35_sumout ),
	.datac(!Xd_0__inst_mult_0_324 ),
	.datad(!Xd_0__inst_mult_0_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_299 ),
	.cout(Xd_0__inst_mult_0_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_105 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[279]),
	.datac(!Xd_0__inst_mult_23_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_319 ),
	.cout(Xd_0__inst_mult_23_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_324 ),
	.datab(!Xd_0__inst_mult_23_319 ),
	.datac(!din_a[286]),
	.datad(!din_b[278]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_329 ),
	.cout(Xd_0__inst_mult_23_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_86 (
// Equation(s):

	.dataa(!din_a[227]),
	.datab(!din_b[227]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_92 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_86_sumout ),
	.cout(Xd_0__inst_i29_87 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_45 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[228]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_45_sumout ),
	.cout(Xd_0__inst_mult_19_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_35 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[216]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_35_sumout ),
	.cout(Xd_0__inst_mult_18_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_35 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_35_sumout ),
	.cout(Xd_0__inst_mult_6_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_294 ),
	.datab(!Xd_0__inst_mult_6_35_sumout ),
	.datac(!Xd_0__inst_mult_6_324 ),
	.datad(!Xd_0__inst_mult_6_55_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_299 ),
	.cout(Xd_0__inst_mult_6_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_91 (
// Equation(s):

	.dataa(!din_a[203]),
	.datab(!din_b[203]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_97 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_91_sumout ),
	.cout(Xd_0__inst_i29_92 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_96 (
// Equation(s):

	.dataa(!din_a[215]),
	.datab(!din_b[215]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_47 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_96_sumout ),
	.cout(Xd_0__inst_i29_97 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_45 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[204]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_45_sumout ),
	.cout(Xd_0__inst_mult_17_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_45 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[192]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_45_sumout ),
	.cout(Xd_0__inst_mult_16_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_35 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_35_sumout ),
	.cout(Xd_0__inst_mult_1_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_294 ),
	.datab(!Xd_0__inst_mult_1_35_sumout ),
	.datac(!Xd_0__inst_mult_1_324 ),
	.datad(!Xd_0__inst_mult_1_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_299 ),
	.cout(Xd_0__inst_mult_1_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_105 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[267]),
	.datac(!Xd_0__inst_mult_22_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_319 ),
	.cout(Xd_0__inst_mult_22_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_324 ),
	.datab(!Xd_0__inst_mult_22_319 ),
	.datac(!din_a[274]),
	.datad(!din_b[266]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_329 ),
	.cout(Xd_0__inst_mult_22_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_144 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[291]),
	.datac(!din_a[294]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_514 ),
	.cout(Xd_0__inst_mult_24_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_145 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_579 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_519 ),
	.cout(Xd_0__inst_mult_24_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_146 (
// Equation(s):

	.dataa(!din_a[296]),
	.datab(!din_b[289]),
	.datac(!din_a[297]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_524 ),
	.cout(Xd_0__inst_mult_24_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_147 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_524 ),
	.datab(!Xd_0__inst_mult_24_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_529 ),
	.cout(Xd_0__inst_mult_24_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_144 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[321]),
	.datac(!din_a[315]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_514 ),
	.cout(Xd_0__inst_mult_26_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_145 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_579 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_519 ),
	.cout(Xd_0__inst_mult_26_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_146 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[318]),
	.datac(!din_a[318]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_524 ),
	.cout(Xd_0__inst_mult_26_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_147 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_589 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_529 ),
	.cout(Xd_0__inst_mult_26_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_148 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_529 ),
	.datab(!Xd_0__inst_mult_26_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_534 ),
	.cout(Xd_0__inst_mult_26_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_101 (
// Equation(s):

	.dataa(!din_a[179]),
	.datab(!din_b[179]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_52 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_101_sumout ),
	.cout(Xd_0__inst_i29_102 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_35 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_35_sumout ),
	.cout(Xd_0__inst_mult_15_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_40 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_40_sumout ),
	.cout(Xd_0__inst_mult_14_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_35 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_35_sumout ),
	.cout(Xd_0__inst_mult_7_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_294 ),
	.datab(!Xd_0__inst_mult_7_35_sumout ),
	.datac(!Xd_0__inst_mult_7_324 ),
	.datad(!Xd_0__inst_mult_7_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_299 ),
	.cout(Xd_0__inst_mult_7_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_106 (
// Equation(s):

	.dataa(!din_a[155]),
	.datab(!din_b[155]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_112 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_106_sumout ),
	.cout(Xd_0__inst_i29_107 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_111 (
// Equation(s):

	.dataa(!din_a[167]),
	.datab(!din_b[167]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_111_sumout ),
	.cout(Xd_0__inst_i29_112 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_40 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_40_sumout ),
	.cout(Xd_0__inst_mult_13_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_35 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_35_sumout ),
	.cout(Xd_0__inst_mult_12_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_35 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[52]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_35_sumout ),
	.cout(Xd_0__inst_mult_4_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_294 ),
	.datab(!Xd_0__inst_mult_4_35_sumout ),
	.datac(!Xd_0__inst_mult_4_324 ),
	.datad(!Xd_0__inst_mult_4_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_299 ),
	.cout(Xd_0__inst_mult_4_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_105 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[231]),
	.datac(!Xd_0__inst_mult_19_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_319 ),
	.cout(Xd_0__inst_mult_19_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_324 ),
	.datab(!Xd_0__inst_mult_19_319 ),
	.datac(!din_a[238]),
	.datad(!din_b[230]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_329 ),
	.cout(Xd_0__inst_mult_19_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_116 (
// Equation(s):

	.dataa(!din_a[131]),
	.datab(!din_b[131]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_122 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_116_sumout ),
	.cout(Xd_0__inst_i29_117 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_40 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_40_sumout ),
	.cout(Xd_0__inst_mult_11_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_40 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_40_sumout ),
	.cout(Xd_0__inst_mult_10_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_294 ),
	.datab(!Xd_0__inst_mult_30_35_sumout ),
	.datac(!Xd_0__inst_mult_30_324 ),
	.datad(!Xd_0__inst_mult_30_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_299 ),
	.cout(Xd_0__inst_mult_30_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_121 (
// Equation(s):

	.dataa(!din_a[107]),
	.datab(!din_b[107]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_127 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_121_sumout ),
	.cout(Xd_0__inst_i29_122 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_126 (
// Equation(s):

	.dataa(!din_a[119]),
	.datab(!din_b[119]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_132 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_126_sumout ),
	.cout(Xd_0__inst_i29_127 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_40 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[108]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_40_sumout ),
	.cout(Xd_0__inst_mult_9_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_40 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_40_sumout ),
	.cout(Xd_0__inst_mult_8_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_35 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[64]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_35_sumout ),
	.cout(Xd_0__inst_mult_5_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_294 ),
	.datab(!Xd_0__inst_mult_5_35_sumout ),
	.datac(!Xd_0__inst_mult_5_324 ),
	.datad(!Xd_0__inst_mult_5_65_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_299 ),
	.cout(Xd_0__inst_mult_5_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_105 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[207]),
	.datac(!Xd_0__inst_mult_17_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_319 ),
	.cout(Xd_0__inst_mult_17_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_324 ),
	.datab(!Xd_0__inst_mult_17_319 ),
	.datac(!din_a[214]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_329 ),
	.cout(Xd_0__inst_mult_17_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_116 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[327]),
	.datac(!din_a[330]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_374 ),
	.cout(Xd_0__inst_mult_27_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_117 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_414 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_379 ),
	.cout(Xd_0__inst_mult_27_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_118 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[325]),
	.datac(!din_a[333]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_384 ),
	.cout(Xd_0__inst_mult_27_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_384 ),
	.datab(!Xd_0__inst_mult_27_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_389 ),
	.cout(Xd_0__inst_mult_27_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_131 (
// Equation(s):

	.dataa(!din_a[83]),
	.datab(!din_b[83]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_137 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_131_sumout ),
	.cout(Xd_0__inst_i29_132 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_40 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_40_sumout ),
	.cout(Xd_0__inst_mult_7_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_40 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_40_sumout ),
	.cout(Xd_0__inst_mult_6_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_45 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[160]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_45_sumout ),
	.cout(Xd_0__inst_mult_13_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_294 ),
	.datab(!Xd_0__inst_mult_13_45_sumout ),
	.datac(!Xd_0__inst_mult_13_324 ),
	.datad(!Xd_0__inst_mult_13_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_299 ),
	.cout(Xd_0__inst_mult_13_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_136 (
// Equation(s):

	.dataa(!din_a[59]),
	.datab(!din_b[59]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_142 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_136_sumout ),
	.cout(Xd_0__inst_i29_137 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_141 (
// Equation(s):

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_147 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_141_sumout ),
	.cout(Xd_0__inst_i29_142 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_40 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_40_sumout ),
	.cout(Xd_0__inst_mult_5_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_40 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_40_sumout ),
	.cout(Xd_0__inst_mult_4_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_110 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_344 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_35 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_35_sumout ),
	.cout(Xd_0__inst_mult_2_36 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_344 ),
	.datab(!Xd_0__inst_mult_2_35_sumout ),
	.datac(!Xd_0__inst_mult_2_379 ),
	.datad(!Xd_0__inst_mult_2_55_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_349 ),
	.cout(Xd_0__inst_mult_2_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_105 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[195]),
	.datac(!Xd_0__inst_mult_16_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_319 ),
	.cout(Xd_0__inst_mult_16_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_324 ),
	.datab(!Xd_0__inst_mult_16_319 ),
	.datac(!din_a[202]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_329 ),
	.cout(Xd_0__inst_mult_16_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_146 (
// Equation(s):

	.dataa(!din_a[35]),
	.datab(!din_b[35]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_146_sumout ),
	.cout(Xd_0__inst_i29_147 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_40 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_40_sumout ),
	.cout(Xd_0__inst_mult_3_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_40 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_40_sumout ),
	.cout(Xd_0__inst_mult_2_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_40 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[340]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_40_sumout ),
	.cout(Xd_0__inst_mult_28_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_294 ),
	.datab(!Xd_0__inst_mult_28_40_sumout ),
	.datac(!Xd_0__inst_mult_28_324 ),
	.datad(!Xd_0__inst_mult_28_60_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_299 ),
	.cout(Xd_0__inst_mult_28_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_151 (
// Equation(s):

	.dataa(!din_a[11]),
	.datab(!din_b[11]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_151_sumout ),
	.cout(Xd_0__inst_i29_152 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("off")
) Xd_0__inst_i29_156 (
// Equation(s):

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_i29_156_sumout ),
	.cout(Xd_0__inst_i29_157 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_40 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_40_sumout ),
	.cout(Xd_0__inst_mult_1_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_40 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_40_sumout ),
	.cout(Xd_0__inst_mult_0_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_100 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_294 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_40 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[376]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_40_sumout ),
	.cout(Xd_0__inst_mult_31_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_294 ),
	.datab(!Xd_0__inst_mult_31_40_sumout ),
	.datac(!Xd_0__inst_mult_31_324 ),
	.datad(!Xd_0__inst_mult_31_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_299 ),
	.cout(Xd_0__inst_mult_31_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_104 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_314 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_105 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[351]),
	.datac(!Xd_0__inst_mult_29_354 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_319 ),
	.cout(Xd_0__inst_mult_29_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_106 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_324 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_324 ),
	.datab(!Xd_0__inst_mult_29_319 ),
	.datac(!din_a[358]),
	.datad(!din_b[350]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_329 ),
	.cout(Xd_0__inst_mult_29_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_149 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[315]),
	.datac(!din_a[318]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_539 ),
	.cout(Xd_0__inst_mult_26_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_150 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_604 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_544 ),
	.cout(Xd_0__inst_mult_26_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_151 (
// Equation(s):

	.dataa(!din_a[320]),
	.datab(!din_b[313]),
	.datac(!din_a[321]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_549 ),
	.cout(Xd_0__inst_mult_26_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_152 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_549 ),
	.datab(!Xd_0__inst_mult_26_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_554 ),
	.cout(Xd_0__inst_mult_26_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_148 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[297]),
	.datac(!din_a[291]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_534 ),
	.cout(Xd_0__inst_mult_24_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_149 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_599 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_539 ),
	.cout(Xd_0__inst_mult_24_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_150 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[294]),
	.datac(!din_a[294]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_544 ),
	.cout(Xd_0__inst_mult_24_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_151 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_609 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_549 ),
	.cout(Xd_0__inst_mult_24_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_152 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_549 ),
	.datab(!Xd_0__inst_mult_24_539 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_554 ),
	.cout(Xd_0__inst_mult_24_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_2_112 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[29]),
	.datac(!din_a[25]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_354 ),
	.cout(Xd_0__inst_mult_2_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_108 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[349]),
	.datac(!din_a[349]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_334 ),
	.cout(Xd_0__inst_mult_29_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_102 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[337]),
	.datac(!din_a[337]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_304 ),
	.cout(Xd_0__inst_mult_28_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_102 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[373]),
	.datac(!din_a[373]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_304 ),
	.cout(Xd_0__inst_mult_31_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_102 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[361]),
	.datac(!din_a[361]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_304 ),
	.cout(Xd_0__inst_mult_30_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_120 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[301]),
	.datac(!din_a[301]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_394 ),
	.cout(Xd_0__inst_mult_25_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_153 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[289]),
	.datac(!din_a[289]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_559 ),
	.cout(Xd_0__inst_mult_24_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_120 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[325]),
	.datac(!din_a[325]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_394 ),
	.cout(Xd_0__inst_mult_27_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_153 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[313]),
	.datac(!din_a[313]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_559 ),
	.cout(Xd_0__inst_mult_26_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_108 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[253]),
	.datac(!din_a[253]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_334 ),
	.cout(Xd_0__inst_mult_21_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_108 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[241]),
	.datac(!din_a[241]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_334 ),
	.cout(Xd_0__inst_mult_20_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_108 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[277]),
	.datac(!din_a[277]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_334 ),
	.cout(Xd_0__inst_mult_23_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_108 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[265]),
	.datac(!din_a[265]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_334 ),
	.cout(Xd_0__inst_mult_22_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_108 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[205]),
	.datac(!din_a[205]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_334 ),
	.cout(Xd_0__inst_mult_17_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_108 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[193]),
	.datac(!din_a[193]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_334 ),
	.cout(Xd_0__inst_mult_16_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_108 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[229]),
	.datac(!din_a[229]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_334 ),
	.cout(Xd_0__inst_mult_19_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_99 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[217]),
	.datac(!din_a[217]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_289 ),
	.cout(Xd_0__inst_mult_18_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_102 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[157]),
	.datac(!din_a[157]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_304 ),
	.cout(Xd_0__inst_mult_13_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_99 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[145]),
	.datac(!din_a[145]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_289 ),
	.cout(Xd_0__inst_mult_12_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_99 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[181]),
	.datac(!din_a[181]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_289 ),
	.cout(Xd_0__inst_mult_15_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_99 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[169]),
	.datac(!din_a[169]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_289 ),
	.cout(Xd_0__inst_mult_14_290 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_102 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[109]),
	.datac(!din_a[109]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_304 ),
	.cout(Xd_0__inst_mult_9_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_102 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[97]),
	.datac(!din_a[97]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_304 ),
	.cout(Xd_0__inst_mult_8_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_102 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[133]),
	.datac(!din_a[133]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_304 ),
	.cout(Xd_0__inst_mult_11_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_102 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[121]),
	.datac(!din_a[121]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_304 ),
	.cout(Xd_0__inst_mult_10_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_102 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[61]),
	.datac(!din_a[61]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_304 ),
	.cout(Xd_0__inst_mult_5_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_102 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[49]),
	.datac(!din_a[49]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_304 ),
	.cout(Xd_0__inst_mult_4_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_102 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[85]),
	.datac(!din_a[85]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_304 ),
	.cout(Xd_0__inst_mult_7_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_102 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[73]),
	.datac(!din_a[73]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_304 ),
	.cout(Xd_0__inst_mult_6_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_102 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[13]),
	.datac(!din_a[13]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_304 ),
	.cout(Xd_0__inst_mult_1_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_102 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[1]),
	.datac(!din_a[1]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_304 ),
	.cout(Xd_0__inst_mult_0_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_102 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[37]),
	.datac(!din_a[37]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_304 ),
	.cout(Xd_0__inst_mult_3_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_113 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[25]),
	.datac(!din_a[25]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_359 ),
	.cout(Xd_0__inst_mult_2_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_374 ),
	.datab(!Xd_0__inst_mult_29_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_339 ),
	.cout(Xd_0__inst_mult_29_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_334 ),
	.datab(!Xd_0__inst_mult_28_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_309 ),
	.cout(Xd_0__inst_mult_28_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_334 ),
	.datab(!Xd_0__inst_mult_31_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_309 ),
	.cout(Xd_0__inst_mult_31_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_334 ),
	.datab(!Xd_0__inst_mult_30_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_309 ),
	.cout(Xd_0__inst_mult_30_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_434 ),
	.datab(!Xd_0__inst_mult_25_439 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_399 ),
	.cout(Xd_0__inst_mult_25_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_154 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_624 ),
	.datab(!Xd_0__inst_mult_24_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_564 ),
	.cout(Xd_0__inst_mult_24_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_434 ),
	.datab(!Xd_0__inst_mult_27_439 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_399 ),
	.cout(Xd_0__inst_mult_27_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_154 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_624 ),
	.datab(!Xd_0__inst_mult_26_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_564 ),
	.cout(Xd_0__inst_mult_26_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_374 ),
	.datab(!Xd_0__inst_mult_21_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_339 ),
	.cout(Xd_0__inst_mult_21_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_374 ),
	.datab(!Xd_0__inst_mult_20_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_339 ),
	.cout(Xd_0__inst_mult_20_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_374 ),
	.datab(!Xd_0__inst_mult_23_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_339 ),
	.cout(Xd_0__inst_mult_23_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_374 ),
	.datab(!Xd_0__inst_mult_22_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_339 ),
	.cout(Xd_0__inst_mult_22_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_374 ),
	.datab(!Xd_0__inst_mult_17_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_339 ),
	.cout(Xd_0__inst_mult_17_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_374 ),
	.datab(!Xd_0__inst_mult_16_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_339 ),
	.cout(Xd_0__inst_mult_16_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_374 ),
	.datab(!Xd_0__inst_mult_19_379 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_339 ),
	.cout(Xd_0__inst_mult_19_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_309 ),
	.datab(!Xd_0__inst_mult_18_314 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_294 ),
	.cout(Xd_0__inst_mult_18_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_334 ),
	.datab(!Xd_0__inst_mult_13_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_309 ),
	.cout(Xd_0__inst_mult_13_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_309 ),
	.datab(!Xd_0__inst_mult_12_314 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_294 ),
	.cout(Xd_0__inst_mult_12_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_309 ),
	.datab(!Xd_0__inst_mult_15_314 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_294 ),
	.cout(Xd_0__inst_mult_15_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_100 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_309 ),
	.datab(!Xd_0__inst_mult_14_314 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_294 ),
	.cout(Xd_0__inst_mult_14_295 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_334 ),
	.datab(!Xd_0__inst_mult_9_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_309 ),
	.cout(Xd_0__inst_mult_9_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_334 ),
	.datab(!Xd_0__inst_mult_8_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_309 ),
	.cout(Xd_0__inst_mult_8_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_334 ),
	.datab(!Xd_0__inst_mult_11_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_309 ),
	.cout(Xd_0__inst_mult_11_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_334 ),
	.datab(!Xd_0__inst_mult_10_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_309 ),
	.cout(Xd_0__inst_mult_10_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_334 ),
	.datab(!Xd_0__inst_mult_5_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_309 ),
	.cout(Xd_0__inst_mult_5_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_334 ),
	.datab(!Xd_0__inst_mult_4_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_309 ),
	.cout(Xd_0__inst_mult_4_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_334 ),
	.datab(!Xd_0__inst_mult_7_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_309 ),
	.cout(Xd_0__inst_mult_7_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_334 ),
	.datab(!Xd_0__inst_mult_6_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_309 ),
	.cout(Xd_0__inst_mult_6_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_334 ),
	.datab(!Xd_0__inst_mult_1_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_309 ),
	.cout(Xd_0__inst_mult_1_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_334 ),
	.datab(!Xd_0__inst_mult_0_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_309 ),
	.cout(Xd_0__inst_mult_0_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_103 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_334 ),
	.datab(!Xd_0__inst_mult_3_339 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_309 ),
	.cout(Xd_0__inst_mult_3_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_394 ),
	.datab(!Xd_0__inst_mult_2_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_364 ),
	.cout(Xd_0__inst_mult_2_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_384 ),
	.datab(!Xd_0__inst_mult_29_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_344 ),
	.cout(Xd_0__inst_mult_29_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_344 ),
	.datab(!Xd_0__inst_mult_28_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_314 ),
	.cout(Xd_0__inst_mult_28_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_344 ),
	.datab(!Xd_0__inst_mult_31_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_314 ),
	.cout(Xd_0__inst_mult_31_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_344 ),
	.datab(!Xd_0__inst_mult_30_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_314 ),
	.cout(Xd_0__inst_mult_30_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_444 ),
	.datab(!Xd_0__inst_mult_25_449 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_404 ),
	.cout(Xd_0__inst_mult_25_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_155 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_634 ),
	.datab(!Xd_0__inst_mult_24_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_569 ),
	.cout(Xd_0__inst_mult_24_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_444 ),
	.datab(!Xd_0__inst_mult_27_449 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_404 ),
	.cout(Xd_0__inst_mult_27_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_155 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_634 ),
	.datab(!Xd_0__inst_mult_26_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_569 ),
	.cout(Xd_0__inst_mult_26_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_384 ),
	.datab(!Xd_0__inst_mult_21_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_344 ),
	.cout(Xd_0__inst_mult_21_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_384 ),
	.datab(!Xd_0__inst_mult_20_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_344 ),
	.cout(Xd_0__inst_mult_20_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_384 ),
	.datab(!Xd_0__inst_mult_23_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_344 ),
	.cout(Xd_0__inst_mult_23_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_384 ),
	.datab(!Xd_0__inst_mult_22_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_344 ),
	.cout(Xd_0__inst_mult_22_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_384 ),
	.datab(!Xd_0__inst_mult_17_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_344 ),
	.cout(Xd_0__inst_mult_17_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_384 ),
	.datab(!Xd_0__inst_mult_16_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_344 ),
	.cout(Xd_0__inst_mult_16_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_110 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_384 ),
	.datab(!Xd_0__inst_mult_19_389 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_344 ),
	.cout(Xd_0__inst_mult_19_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_319 ),
	.datab(!Xd_0__inst_mult_18_324 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_299 ),
	.cout(Xd_0__inst_mult_18_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_344 ),
	.datab(!Xd_0__inst_mult_13_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_314 ),
	.cout(Xd_0__inst_mult_13_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_319 ),
	.datab(!Xd_0__inst_mult_12_324 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_299 ),
	.cout(Xd_0__inst_mult_12_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_319 ),
	.datab(!Xd_0__inst_mult_15_324 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_299 ),
	.cout(Xd_0__inst_mult_15_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_101 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_319 ),
	.datab(!Xd_0__inst_mult_14_324 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_295 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_299 ),
	.cout(Xd_0__inst_mult_14_300 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_344 ),
	.datab(!Xd_0__inst_mult_9_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_314 ),
	.cout(Xd_0__inst_mult_9_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_344 ),
	.datab(!Xd_0__inst_mult_8_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_314 ),
	.cout(Xd_0__inst_mult_8_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_344 ),
	.datab(!Xd_0__inst_mult_11_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_314 ),
	.cout(Xd_0__inst_mult_11_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_344 ),
	.datab(!Xd_0__inst_mult_10_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_314 ),
	.cout(Xd_0__inst_mult_10_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_344 ),
	.datab(!Xd_0__inst_mult_5_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_314 ),
	.cout(Xd_0__inst_mult_5_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_344 ),
	.datab(!Xd_0__inst_mult_4_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_314 ),
	.cout(Xd_0__inst_mult_4_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_344 ),
	.datab(!Xd_0__inst_mult_7_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_314 ),
	.cout(Xd_0__inst_mult_7_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_344 ),
	.datab(!Xd_0__inst_mult_6_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_314 ),
	.cout(Xd_0__inst_mult_6_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_344 ),
	.datab(!Xd_0__inst_mult_1_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_314 ),
	.cout(Xd_0__inst_mult_1_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_344 ),
	.datab(!Xd_0__inst_mult_0_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_314 ),
	.cout(Xd_0__inst_mult_0_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_104 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_344 ),
	.datab(!Xd_0__inst_mult_3_349 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_314 ),
	.cout(Xd_0__inst_mult_3_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_404 ),
	.datab(!Xd_0__inst_mult_2_409 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_369 ),
	.cout(Xd_0__inst_mult_2_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_394 ),
	.datab(!Xd_0__inst_mult_29_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_349 ),
	.cout(Xd_0__inst_mult_29_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_354 ),
	.datab(!Xd_0__inst_mult_28_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_319 ),
	.cout(Xd_0__inst_mult_28_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_354 ),
	.datab(!Xd_0__inst_mult_31_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_319 ),
	.cout(Xd_0__inst_mult_31_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_354 ),
	.datab(!Xd_0__inst_mult_30_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_319 ),
	.cout(Xd_0__inst_mult_30_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_454 ),
	.datab(!Xd_0__inst_mult_25_459 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_409 ),
	.cout(Xd_0__inst_mult_25_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_156 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_644 ),
	.datab(!Xd_0__inst_mult_24_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_574 ),
	.cout(Xd_0__inst_mult_24_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_454 ),
	.datab(!Xd_0__inst_mult_27_459 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_409 ),
	.cout(Xd_0__inst_mult_27_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_156 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_644 ),
	.datab(!Xd_0__inst_mult_26_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_574 ),
	.cout(Xd_0__inst_mult_26_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_394 ),
	.datab(!Xd_0__inst_mult_21_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_349 ),
	.cout(Xd_0__inst_mult_21_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_394 ),
	.datab(!Xd_0__inst_mult_20_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_349 ),
	.cout(Xd_0__inst_mult_20_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_394 ),
	.datab(!Xd_0__inst_mult_23_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_349 ),
	.cout(Xd_0__inst_mult_23_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_394 ),
	.datab(!Xd_0__inst_mult_22_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_349 ),
	.cout(Xd_0__inst_mult_22_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_394 ),
	.datab(!Xd_0__inst_mult_17_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_349 ),
	.cout(Xd_0__inst_mult_17_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_394 ),
	.datab(!Xd_0__inst_mult_16_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_349 ),
	.cout(Xd_0__inst_mult_16_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_394 ),
	.datab(!Xd_0__inst_mult_19_399 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_349 ),
	.cout(Xd_0__inst_mult_19_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_329 ),
	.datab(!Xd_0__inst_mult_18_334 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_304 ),
	.cout(Xd_0__inst_mult_18_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_354 ),
	.datab(!Xd_0__inst_mult_13_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_319 ),
	.cout(Xd_0__inst_mult_13_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_329 ),
	.datab(!Xd_0__inst_mult_12_334 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_304 ),
	.cout(Xd_0__inst_mult_12_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_329 ),
	.datab(!Xd_0__inst_mult_15_334 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_304 ),
	.cout(Xd_0__inst_mult_15_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_102 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_329 ),
	.datab(!Xd_0__inst_mult_14_334 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_300 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_304 ),
	.cout(Xd_0__inst_mult_14_305 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_354 ),
	.datab(!Xd_0__inst_mult_9_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_319 ),
	.cout(Xd_0__inst_mult_9_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_354 ),
	.datab(!Xd_0__inst_mult_8_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_319 ),
	.cout(Xd_0__inst_mult_8_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_354 ),
	.datab(!Xd_0__inst_mult_11_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_319 ),
	.cout(Xd_0__inst_mult_11_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_354 ),
	.datab(!Xd_0__inst_mult_10_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_319 ),
	.cout(Xd_0__inst_mult_10_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_354 ),
	.datab(!Xd_0__inst_mult_5_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_319 ),
	.cout(Xd_0__inst_mult_5_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_354 ),
	.datab(!Xd_0__inst_mult_4_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_319 ),
	.cout(Xd_0__inst_mult_4_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_354 ),
	.datab(!Xd_0__inst_mult_7_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_319 ),
	.cout(Xd_0__inst_mult_7_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_354 ),
	.datab(!Xd_0__inst_mult_6_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_319 ),
	.cout(Xd_0__inst_mult_6_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_354 ),
	.datab(!Xd_0__inst_mult_1_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_319 ),
	.cout(Xd_0__inst_mult_1_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_354 ),
	.datab(!Xd_0__inst_mult_0_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_319 ),
	.cout(Xd_0__inst_mult_0_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_105 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_354 ),
	.datab(!Xd_0__inst_mult_3_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_319 ),
	.cout(Xd_0__inst_mult_3_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_414 ),
	.datab(!Xd_0__inst_mult_2_419 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_374 ),
	.cout(Xd_0__inst_mult_2_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_40 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[226]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_40_sumout ),
	.cout(Xd_0__inst_mult_18_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_50 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[214]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_50_sumout ),
	.cout(Xd_0__inst_mult_17_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_55 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[250]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_55_sumout ),
	.cout(Xd_0__inst_mult_20_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_45 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_45_sumout ),
	.cout(Xd_0__inst_mult_2_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_55 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[310]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_55_sumout ),
	.cout(Xd_0__inst_mult_25_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_45 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[346]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_45_sumout ),
	.cout(Xd_0__inst_mult_28_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_45 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_45_sumout ),
	.cout(Xd_0__inst_mult_3_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_45 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_45_sumout ),
	.cout(Xd_0__inst_mult_6_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_45 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_45_sumout ),
	.cout(Xd_0__inst_mult_8_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_50 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[105]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_50_sumout ),
	.cout(Xd_0__inst_mult_8_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_40 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_40_sumout ),
	.cout(Xd_0__inst_mult_15_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_45 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_45_sumout ),
	.cout(Xd_0__inst_mult_5_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_50 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_50_sumout ),
	.cout(Xd_0__inst_mult_2_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_45 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[171]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_45_sumout ),
	.cout(Xd_0__inst_mult_14_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_45 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[135]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_45_sumout ),
	.cout(Xd_0__inst_mult_11_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_45 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[51]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_45_sumout ),
	.cout(Xd_0__inst_mult_4_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_45 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[15]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_45_sumout ),
	.cout(Xd_0__inst_mult_1_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_55 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[27]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_55_sumout ),
	.cout(Xd_0__inst_mult_2_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_45 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[3]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_45_sumout ),
	.cout(Xd_0__inst_mult_0_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_45 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[375]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_45_sumout ),
	.cout(Xd_0__inst_mult_31_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_60 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[310]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_60_sumout ),
	.cout(Xd_0__inst_mult_25_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_50 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[346]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_50_sumout ),
	.cout(Xd_0__inst_mult_28_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_50 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_50_sumout ),
	.cout(Xd_0__inst_mult_3_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_60 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[334]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_60_sumout ),
	.cout(Xd_0__inst_mult_27_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_50 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_50_sumout ),
	.cout(Xd_0__inst_mult_5_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_55 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[105]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_55_sumout ),
	.cout(Xd_0__inst_mult_8_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_45 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[189]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_45_sumout ),
	.cout(Xd_0__inst_mult_15_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_50 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_50_sumout ),
	.cout(Xd_0__inst_mult_6_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_55 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_55_sumout ),
	.cout(Xd_0__inst_mult_5_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_45 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[224]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_45_sumout ),
	.cout(Xd_0__inst_mult_18_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_106 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[112]),
	.datac(!Xd_0__inst_mult_9_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_324 ),
	.cout(Xd_0__inst_mult_9_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_45 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[111]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_45_sumout ),
	.cout(Xd_0__inst_mult_9_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_324 ),
	.datab(!Xd_0__inst_mult_9_45_sumout ),
	.datac(!Xd_0__inst_mult_9_494 ),
	.datad(!Xd_0__inst_mult_9_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_329 ),
	.cout(Xd_0__inst_mult_9_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_60 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_60_sumout ),
	.cout(Xd_0__inst_mult_5_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_106 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[100]),
	.datac(!Xd_0__inst_mult_8_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_324 ),
	.cout(Xd_0__inst_mult_8_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_60 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[99]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_60_sumout ),
	.cout(Xd_0__inst_mult_8_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_324 ),
	.datab(!Xd_0__inst_mult_8_60_sumout ),
	.datac(!Xd_0__inst_mult_8_494 ),
	.datad(!Xd_0__inst_mult_8_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_329 ),
	.cout(Xd_0__inst_mult_8_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_112 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[256]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_354 ),
	.cout(Xd_0__inst_mult_21_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_113 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_359 ),
	.cout(Xd_0__inst_mult_21_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_114 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[253]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_364 ),
	.cout(Xd_0__inst_mult_21_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_364 ),
	.datab(!Xd_0__inst_mult_21_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_369 ),
	.cout(Xd_0__inst_mult_21_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_106 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[136]),
	.datac(!Xd_0__inst_mult_11_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_324 ),
	.cout(Xd_0__inst_mult_11_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_324 ),
	.datab(!Xd_0__inst_mult_11_45_sumout ),
	.datac(!Xd_0__inst_mult_11_494 ),
	.datad(!Xd_0__inst_mult_11_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_329 ),
	.cout(Xd_0__inst_mult_11_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_106 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[124]),
	.datac(!Xd_0__inst_mult_10_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_324 ),
	.cout(Xd_0__inst_mult_10_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_45 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[123]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_45_sumout ),
	.cout(Xd_0__inst_mult_10_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_324 ),
	.datab(!Xd_0__inst_mult_10_45_sumout ),
	.datac(!Xd_0__inst_mult_10_494 ),
	.datad(!Xd_0__inst_mult_10_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_329 ),
	.cout(Xd_0__inst_mult_10_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_112 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[244]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_354 ),
	.cout(Xd_0__inst_mult_20_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_113 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_359 ),
	.cout(Xd_0__inst_mult_20_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_50 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[189]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_50_sumout ),
	.cout(Xd_0__inst_mult_15_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_114 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[241]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_364 ),
	.cout(Xd_0__inst_mult_20_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_364 ),
	.datab(!Xd_0__inst_mult_20_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_369 ),
	.cout(Xd_0__inst_mult_20_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_124 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[303]),
	.datac(!din_a[305]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_414 ),
	.cout(Xd_0__inst_mult_25_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_125 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_559 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_419 ),
	.cout(Xd_0__inst_mult_25_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_126 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[301]),
	.datac(!din_a[308]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_424 ),
	.cout(Xd_0__inst_mult_25_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_424 ),
	.datab(!Xd_0__inst_mult_25_419 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_429 ),
	.cout(Xd_0__inst_mult_25_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_106 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[40]),
	.datac(!Xd_0__inst_mult_3_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_324 ),
	.cout(Xd_0__inst_mult_3_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_55 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[184]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_55_sumout ),
	.cout(Xd_0__inst_mult_15_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_55 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[39]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_55_sumout ),
	.cout(Xd_0__inst_mult_3_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_324 ),
	.datab(!Xd_0__inst_mult_3_55_sumout ),
	.datac(!Xd_0__inst_mult_3_494 ),
	.datad(!Xd_0__inst_mult_3_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_329 ),
	.cout(Xd_0__inst_mult_3_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_106 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[4]),
	.datac(!Xd_0__inst_mult_0_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_324 ),
	.cout(Xd_0__inst_mult_0_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_324 ),
	.datab(!Xd_0__inst_mult_0_45_sumout ),
	.datac(!Xd_0__inst_mult_0_494 ),
	.datad(!Xd_0__inst_mult_0_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_329 ),
	.cout(Xd_0__inst_mult_0_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_112 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[280]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_354 ),
	.cout(Xd_0__inst_mult_23_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_113 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_359 ),
	.cout(Xd_0__inst_mult_23_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_114 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[277]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_364 ),
	.cout(Xd_0__inst_mult_23_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_364 ),
	.datab(!Xd_0__inst_mult_23_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_369 ),
	.cout(Xd_0__inst_mult_23_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_55 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[210]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_55_sumout ),
	.cout(Xd_0__inst_mult_17_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_50 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[198]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_50_sumout ),
	.cout(Xd_0__inst_mult_16_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_106 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[76]),
	.datac(!Xd_0__inst_mult_6_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_324 ),
	.cout(Xd_0__inst_mult_6_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_55 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[75]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_55_sumout ),
	.cout(Xd_0__inst_mult_6_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_324 ),
	.datab(!Xd_0__inst_mult_6_55_sumout ),
	.datac(!Xd_0__inst_mult_6_494 ),
	.datad(!Xd_0__inst_mult_6_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_329 ),
	.cout(Xd_0__inst_mult_6_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_106 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[16]),
	.datac(!Xd_0__inst_mult_1_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_324 ),
	.cout(Xd_0__inst_mult_1_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_324 ),
	.datab(!Xd_0__inst_mult_1_45_sumout ),
	.datac(!Xd_0__inst_mult_1_494 ),
	.datad(!Xd_0__inst_mult_1_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_329 ),
	.cout(Xd_0__inst_mult_1_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_112 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[268]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_354 ),
	.cout(Xd_0__inst_mult_22_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_113 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_359 ),
	.cout(Xd_0__inst_mult_22_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_114 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[265]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_364 ),
	.cout(Xd_0__inst_mult_22_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_364 ),
	.datab(!Xd_0__inst_mult_22_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_369 ),
	.cout(Xd_0__inst_mult_22_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_157 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[291]),
	.datac(!din_a[293]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_579 ),
	.cout(Xd_0__inst_mult_24_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_158 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_584 ),
	.cout(Xd_0__inst_mult_24_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_159 (
// Equation(s):

	.dataa(!din_a[295]),
	.datab(!din_b[289]),
	.datac(!din_a[296]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_589 ),
	.cout(Xd_0__inst_mult_24_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_160 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_589 ),
	.datab(!Xd_0__inst_mult_24_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_594 ),
	.cout(Xd_0__inst_mult_24_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_157 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[321]),
	.datac(!din_a[314]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_579 ),
	.cout(Xd_0__inst_mult_26_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_158 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[320]),
	.datac(!Xd_0__inst_mult_26_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_235 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_584 ),
	.cout(Xd_0__inst_mult_26_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_159 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[318]),
	.datac(!din_a[317]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_589 ),
	.cout(Xd_0__inst_mult_26_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_160 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_594 ),
	.cout(Xd_0__inst_mult_26_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_161 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_594 ),
	.datab(!Xd_0__inst_mult_26_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_599 ),
	.cout(Xd_0__inst_mult_26_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_106 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[88]),
	.datac(!Xd_0__inst_mult_7_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_324 ),
	.cout(Xd_0__inst_mult_7_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_45 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[87]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_45_sumout ),
	.cout(Xd_0__inst_mult_7_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_324 ),
	.datab(!Xd_0__inst_mult_7_45_sumout ),
	.datac(!Xd_0__inst_mult_7_494 ),
	.datad(!Xd_0__inst_mult_7_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_329 ),
	.cout(Xd_0__inst_mult_7_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_106 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[52]),
	.datac(!Xd_0__inst_mult_4_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_324 ),
	.cout(Xd_0__inst_mult_4_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_324 ),
	.datab(!Xd_0__inst_mult_4_45_sumout ),
	.datac(!Xd_0__inst_mult_4_494 ),
	.datad(!Xd_0__inst_mult_4_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_329 ),
	.cout(Xd_0__inst_mult_4_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_112 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[232]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_354 ),
	.cout(Xd_0__inst_mult_19_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_113 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_359 ),
	.cout(Xd_0__inst_mult_19_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_114 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[229]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_364 ),
	.cout(Xd_0__inst_mult_19_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_364 ),
	.datab(!Xd_0__inst_mult_19_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_369 ),
	.cout(Xd_0__inst_mult_19_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_106 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[364]),
	.datac(!Xd_0__inst_mult_30_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_324 ),
	.cout(Xd_0__inst_mult_30_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_45 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[363]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_45_sumout ),
	.cout(Xd_0__inst_mult_30_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_324 ),
	.datab(!Xd_0__inst_mult_30_45_sumout ),
	.datac(!Xd_0__inst_mult_30_494 ),
	.datad(!Xd_0__inst_mult_30_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_329 ),
	.cout(Xd_0__inst_mult_30_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_55 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[342]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_55_sumout ),
	.cout(Xd_0__inst_mult_28_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_106 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[64]),
	.datac(!Xd_0__inst_mult_5_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_324 ),
	.cout(Xd_0__inst_mult_5_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_65 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[63]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_65_sumout ),
	.cout(Xd_0__inst_mult_5_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_324 ),
	.datab(!Xd_0__inst_mult_5_65_sumout ),
	.datac(!Xd_0__inst_mult_5_494 ),
	.datad(!Xd_0__inst_mult_5_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_329 ),
	.cout(Xd_0__inst_mult_5_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_112 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[208]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_354 ),
	.cout(Xd_0__inst_mult_17_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_113 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_359 ),
	.cout(Xd_0__inst_mult_17_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_114 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[205]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_364 ),
	.cout(Xd_0__inst_mult_17_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_364 ),
	.datab(!Xd_0__inst_mult_17_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_369 ),
	.cout(Xd_0__inst_mult_17_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_124 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[327]),
	.datac(!din_a[329]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_414 ),
	.cout(Xd_0__inst_mult_27_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_125 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_559 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_419 ),
	.cout(Xd_0__inst_mult_27_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_126 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[325]),
	.datac(!din_a[332]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_424 ),
	.cout(Xd_0__inst_mult_27_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_424 ),
	.datab(!Xd_0__inst_mult_27_419 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_429 ),
	.cout(Xd_0__inst_mult_27_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_50 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[378]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_50_sumout ),
	.cout(Xd_0__inst_mult_31_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_106 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[160]),
	.datac(!Xd_0__inst_mult_13_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_324 ),
	.cout(Xd_0__inst_mult_13_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_50 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[220]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_50_sumout ),
	.cout(Xd_0__inst_mult_18_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_50 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[159]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_50_sumout ),
	.cout(Xd_0__inst_mult_13_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_324 ),
	.datab(!Xd_0__inst_mult_13_50_sumout ),
	.datac(!Xd_0__inst_mult_13_494 ),
	.datad(!Xd_0__inst_mult_13_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_329 ),
	.cout(Xd_0__inst_mult_13_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_117 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[28]),
	.datac(!Xd_0__inst_mult_2_529 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_379 ),
	.cout(Xd_0__inst_mult_2_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_379 ),
	.datab(!Xd_0__inst_mult_2_55_sumout ),
	.datac(!Xd_0__inst_mult_2_539 ),
	.datad(!Xd_0__inst_mult_2_534 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_384 ),
	.cout(Xd_0__inst_mult_2_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_112 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[196]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_354 ),
	.cout(Xd_0__inst_mult_16_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_113 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_359 ),
	.cout(Xd_0__inst_mult_16_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_114 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[193]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_364 ),
	.cout(Xd_0__inst_mult_16_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_364 ),
	.datab(!Xd_0__inst_mult_16_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_369 ),
	.cout(Xd_0__inst_mult_16_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_106 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[340]),
	.datac(!Xd_0__inst_mult_28_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_324 ),
	.cout(Xd_0__inst_mult_28_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_60 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[339]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_60_sumout ),
	.cout(Xd_0__inst_mult_28_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_324 ),
	.datab(!Xd_0__inst_mult_28_60_sumout ),
	.datac(!Xd_0__inst_mult_28_494 ),
	.datad(!Xd_0__inst_mult_28_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_329 ),
	.cout(Xd_0__inst_mult_28_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_70 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_70_sumout ),
	.cout(Xd_0__inst_mult_5_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_106 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[376]),
	.datac(!Xd_0__inst_mult_31_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_324 ),
	.cout(Xd_0__inst_mult_31_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_107 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_324 ),
	.datab(!Xd_0__inst_mult_31_45_sumout ),
	.datac(!Xd_0__inst_mult_31_494 ),
	.datad(!Xd_0__inst_mult_31_489 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_329 ),
	.cout(Xd_0__inst_mult_31_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_112 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[352]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_354 ),
	.cout(Xd_0__inst_mult_29_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_113 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_514 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_359 ),
	.cout(Xd_0__inst_mult_29_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_114 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[349]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_364 ),
	.cout(Xd_0__inst_mult_29_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_364 ),
	.datab(!Xd_0__inst_mult_29_359 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_369 ),
	.cout(Xd_0__inst_mult_29_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_162 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[315]),
	.datac(!din_a[317]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_604 ),
	.cout(Xd_0__inst_mult_26_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_163 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_609 ),
	.cout(Xd_0__inst_mult_26_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_164 (
// Equation(s):

	.dataa(!din_a[319]),
	.datab(!din_b[313]),
	.datac(!din_a[320]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_614 ),
	.cout(Xd_0__inst_mult_26_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_165 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_614 ),
	.datab(!Xd_0__inst_mult_26_609 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_619 ),
	.cout(Xd_0__inst_mult_26_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_161 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[297]),
	.datac(!din_a[290]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_599 ),
	.cout(Xd_0__inst_mult_24_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_162 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[296]),
	.datac(!Xd_0__inst_mult_24_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_245 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_604 ),
	.cout(Xd_0__inst_mult_24_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_163 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[294]),
	.datac(!din_a[293]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_609 ),
	.cout(Xd_0__inst_mult_24_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_164 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_614 ),
	.cout(Xd_0__inst_mult_24_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_165 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_614 ),
	.datab(!Xd_0__inst_mult_24_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_619 ),
	.cout(Xd_0__inst_mult_24_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_119 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[29]),
	.datac(!din_a[24]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_389 ),
	.cout(Xd_0__inst_mult_2_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_116 (
// Equation(s):

	.dataa(!din_a[349]),
	.datab(!din_b[349]),
	.datac(!din_a[350]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_374 ),
	.cout(Xd_0__inst_mult_29_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_29_117 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[350]),
	.datac(!din_a[349]),
	.datad(!din_b[351]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_379 ),
	.cout(Xd_0__inst_mult_29_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_108 (
// Equation(s):

	.dataa(!din_a[337]),
	.datab(!din_b[337]),
	.datac(!din_a[338]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_334 ),
	.cout(Xd_0__inst_mult_28_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_28_109 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[338]),
	.datac(!din_a[337]),
	.datad(!din_b[339]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_339 ),
	.cout(Xd_0__inst_mult_28_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_108 (
// Equation(s):

	.dataa(!din_a[373]),
	.datab(!din_b[373]),
	.datac(!din_a[374]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_334 ),
	.cout(Xd_0__inst_mult_31_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_31_109 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[374]),
	.datac(!din_a[373]),
	.datad(!din_b[375]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_339 ),
	.cout(Xd_0__inst_mult_31_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_40 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[147]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_40_sumout ),
	.cout(Xd_0__inst_mult_12_41 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_108 (
// Equation(s):

	.dataa(!din_a[361]),
	.datab(!din_b[361]),
	.datac(!din_a[362]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_334 ),
	.cout(Xd_0__inst_mult_30_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_30_109 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[362]),
	.datac(!din_a[361]),
	.datad(!din_b[363]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_339 ),
	.cout(Xd_0__inst_mult_30_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_128 (
// Equation(s):

	.dataa(!din_a[301]),
	.datab(!din_b[301]),
	.datac(!din_a[302]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_434 ),
	.cout(Xd_0__inst_mult_25_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_25_129 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[302]),
	.datac(!din_a[301]),
	.datad(!din_b[303]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_439 ),
	.cout(Xd_0__inst_mult_25_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_166 (
// Equation(s):

	.dataa(!din_a[289]),
	.datab(!din_b[289]),
	.datac(!din_a[290]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_624 ),
	.cout(Xd_0__inst_mult_24_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_24_167 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[290]),
	.datac(!din_a[289]),
	.datad(!din_b[291]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_629 ),
	.cout(Xd_0__inst_mult_24_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_128 (
// Equation(s):

	.dataa(!din_a[325]),
	.datab(!din_b[325]),
	.datac(!din_a[326]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_434 ),
	.cout(Xd_0__inst_mult_27_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_27_129 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[326]),
	.datac(!din_a[325]),
	.datad(!din_b[327]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_439 ),
	.cout(Xd_0__inst_mult_27_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_166 (
// Equation(s):

	.dataa(!din_a[313]),
	.datab(!din_b[313]),
	.datac(!din_a[314]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_624 ),
	.cout(Xd_0__inst_mult_26_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_26_167 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[314]),
	.datac(!din_a[313]),
	.datad(!din_b[315]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_629 ),
	.cout(Xd_0__inst_mult_26_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_116 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[253]),
	.datac(!din_a[254]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_374 ),
	.cout(Xd_0__inst_mult_21_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_21_117 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[254]),
	.datac(!din_a[253]),
	.datad(!din_b[255]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_379 ),
	.cout(Xd_0__inst_mult_21_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_116 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[241]),
	.datac(!din_a[242]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_374 ),
	.cout(Xd_0__inst_mult_20_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_20_117 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[242]),
	.datac(!din_a[241]),
	.datad(!din_b[243]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_379 ),
	.cout(Xd_0__inst_mult_20_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_116 (
// Equation(s):

	.dataa(!din_a[277]),
	.datab(!din_b[277]),
	.datac(!din_a[278]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_374 ),
	.cout(Xd_0__inst_mult_23_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_23_117 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[278]),
	.datac(!din_a[277]),
	.datad(!din_b[279]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_379 ),
	.cout(Xd_0__inst_mult_23_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_116 (
// Equation(s):

	.dataa(!din_a[265]),
	.datab(!din_b[265]),
	.datac(!din_a[266]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_374 ),
	.cout(Xd_0__inst_mult_22_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_22_117 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[266]),
	.datac(!din_a[265]),
	.datad(!din_b[267]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_379 ),
	.cout(Xd_0__inst_mult_22_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_116 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[205]),
	.datac(!din_a[206]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_374 ),
	.cout(Xd_0__inst_mult_17_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_17_117 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[206]),
	.datac(!din_a[205]),
	.datad(!din_b[207]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_379 ),
	.cout(Xd_0__inst_mult_17_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_116 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[193]),
	.datac(!din_a[194]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_374 ),
	.cout(Xd_0__inst_mult_16_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_16_117 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[194]),
	.datac(!din_a[193]),
	.datad(!din_b[195]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_379 ),
	.cout(Xd_0__inst_mult_16_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_116 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[229]),
	.datac(!din_a[230]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_374 ),
	.cout(Xd_0__inst_mult_19_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_19_117 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[230]),
	.datac(!din_a[229]),
	.datad(!din_b[231]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_379 ),
	.cout(Xd_0__inst_mult_19_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_103 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[217]),
	.datac(!din_a[218]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_309 ),
	.cout(Xd_0__inst_mult_18_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_18_104 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[218]),
	.datac(!din_a[217]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_314 ),
	.cout(Xd_0__inst_mult_18_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_60 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[214]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_60_sumout ),
	.cout(Xd_0__inst_mult_17_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_108 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[157]),
	.datac(!din_a[158]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_334 ),
	.cout(Xd_0__inst_mult_13_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_13_109 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[158]),
	.datac(!din_a[157]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_339 ),
	.cout(Xd_0__inst_mult_13_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_103 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[145]),
	.datac(!din_a[146]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_309 ),
	.cout(Xd_0__inst_mult_12_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_12_104 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[146]),
	.datac(!din_a[145]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_314 ),
	.cout(Xd_0__inst_mult_12_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_60 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_60_sumout ),
	.cout(Xd_0__inst_mult_15_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_103 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[181]),
	.datac(!din_a[182]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_309 ),
	.cout(Xd_0__inst_mult_15_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_15_104 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[182]),
	.datac(!din_a[181]),
	.datad(!din_b[183]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_314 ),
	.cout(Xd_0__inst_mult_15_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_75 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_75_sumout ),
	.cout(Xd_0__inst_mult_5_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_103 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[169]),
	.datac(!din_a[170]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_290 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_309 ),
	.cout(Xd_0__inst_mult_14_310 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_14_104 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[170]),
	.datac(!din_a[169]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_325 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_314 ),
	.cout(Xd_0__inst_mult_14_315 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_60 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_60_sumout ),
	.cout(Xd_0__inst_mult_3_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_108 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[109]),
	.datac(!din_a[110]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_334 ),
	.cout(Xd_0__inst_mult_9_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_9_109 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[110]),
	.datac(!din_a[109]),
	.datad(!din_b[111]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_339 ),
	.cout(Xd_0__inst_mult_9_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_108 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[97]),
	.datac(!din_a[98]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_334 ),
	.cout(Xd_0__inst_mult_8_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_8_109 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[98]),
	.datac(!din_a[97]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_339 ),
	.cout(Xd_0__inst_mult_8_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_108 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[133]),
	.datac(!din_a[134]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_334 ),
	.cout(Xd_0__inst_mult_11_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_11_109 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[134]),
	.datac(!din_a[133]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_339 ),
	.cout(Xd_0__inst_mult_11_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_108 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[121]),
	.datac(!din_a[122]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_334 ),
	.cout(Xd_0__inst_mult_10_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_10_109 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[122]),
	.datac(!din_a[121]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_339 ),
	.cout(Xd_0__inst_mult_10_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_108 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[61]),
	.datac(!din_a[62]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_334 ),
	.cout(Xd_0__inst_mult_5_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_5_109 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[62]),
	.datac(!din_a[61]),
	.datad(!din_b[63]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_339 ),
	.cout(Xd_0__inst_mult_5_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_108 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_334 ),
	.cout(Xd_0__inst_mult_4_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_4_109 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[50]),
	.datac(!din_a[49]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_339 ),
	.cout(Xd_0__inst_mult_4_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_108 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_334 ),
	.cout(Xd_0__inst_mult_7_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_7_109 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[86]),
	.datac(!din_a[85]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_339 ),
	.cout(Xd_0__inst_mult_7_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_108 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_334 ),
	.cout(Xd_0__inst_mult_6_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_6_109 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[74]),
	.datac(!din_a[73]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_339 ),
	.cout(Xd_0__inst_mult_6_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_108 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(!din_a[14]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_334 ),
	.cout(Xd_0__inst_mult_1_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_1_109 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[14]),
	.datac(!din_a[13]),
	.datad(!din_b[15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_339 ),
	.cout(Xd_0__inst_mult_1_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_108 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_334 ),
	.cout(Xd_0__inst_mult_0_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_0_109 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[2]),
	.datac(!din_a[1]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_339 ),
	.cout(Xd_0__inst_mult_0_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_108 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[38]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_334 ),
	.cout(Xd_0__inst_mult_3_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_3_109 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[38]),
	.datac(!din_a[37]),
	.datad(!din_b[39]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_339 ),
	.cout(Xd_0__inst_mult_3_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_65 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[183]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_65_sumout ),
	.cout(Xd_0__inst_mult_15_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_120 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_394 ),
	.cout(Xd_0__inst_mult_2_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_2_121 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[26]),
	.datac(!din_a[25]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_399 ),
	.cout(Xd_0__inst_mult_2_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_55 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[219]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_55_sumout ),
	.cout(Xd_0__inst_mult_18_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_118 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[349]),
	.datac(!din_a[351]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_384 ),
	.cout(Xd_0__inst_mult_29_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_119 (
// Equation(s):

	.dataa(!din_a[349]),
	.datab(!din_b[350]),
	.datac(!din_a[348]),
	.datad(!din_b[351]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_389 ),
	.cout(Xd_0__inst_mult_29_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_110 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[337]),
	.datac(!din_a[339]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_344 ),
	.cout(Xd_0__inst_mult_28_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_111 (
// Equation(s):

	.dataa(!din_a[337]),
	.datab(!din_b[338]),
	.datac(!din_a[336]),
	.datad(!din_b[339]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_349 ),
	.cout(Xd_0__inst_mult_28_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_110 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[373]),
	.datac(!din_a[375]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_344 ),
	.cout(Xd_0__inst_mult_31_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_111 (
// Equation(s):

	.dataa(!din_a[373]),
	.datab(!din_b[374]),
	.datac(!din_a[372]),
	.datad(!din_b[375]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_349 ),
	.cout(Xd_0__inst_mult_31_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_110 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[361]),
	.datac(!din_a[363]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_344 ),
	.cout(Xd_0__inst_mult_30_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_111 (
// Equation(s):

	.dataa(!din_a[361]),
	.datab(!din_b[362]),
	.datac(!din_a[360]),
	.datad(!din_b[363]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_349 ),
	.cout(Xd_0__inst_mult_30_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_130 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[301]),
	.datac(!din_a[303]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_444 ),
	.cout(Xd_0__inst_mult_25_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_131 (
// Equation(s):

	.dataa(!din_a[301]),
	.datab(!din_b[302]),
	.datac(!din_a[300]),
	.datad(!din_b[303]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_449 ),
	.cout(Xd_0__inst_mult_25_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_168 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[289]),
	.datac(!din_a[291]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_634 ),
	.cout(Xd_0__inst_mult_24_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_169 (
// Equation(s):

	.dataa(!din_a[289]),
	.datab(!din_b[290]),
	.datac(!din_a[288]),
	.datad(!din_b[291]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_639 ),
	.cout(Xd_0__inst_mult_24_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_130 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[325]),
	.datac(!din_a[327]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_444 ),
	.cout(Xd_0__inst_mult_27_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_131 (
// Equation(s):

	.dataa(!din_a[325]),
	.datab(!din_b[326]),
	.datac(!din_a[324]),
	.datad(!din_b[327]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_449 ),
	.cout(Xd_0__inst_mult_27_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_168 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[313]),
	.datac(!din_a[315]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_634 ),
	.cout(Xd_0__inst_mult_26_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_169 (
// Equation(s):

	.dataa(!din_a[313]),
	.datab(!din_b[314]),
	.datac(!din_a[312]),
	.datad(!din_b[315]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_639 ),
	.cout(Xd_0__inst_mult_26_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_118 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[253]),
	.datac(!din_a[255]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_384 ),
	.cout(Xd_0__inst_mult_21_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_119 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[254]),
	.datac(!din_a[252]),
	.datad(!din_b[255]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_389 ),
	.cout(Xd_0__inst_mult_21_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_118 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[241]),
	.datac(!din_a[243]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_384 ),
	.cout(Xd_0__inst_mult_20_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_119 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[242]),
	.datac(!din_a[240]),
	.datad(!din_b[243]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_389 ),
	.cout(Xd_0__inst_mult_20_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_118 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[277]),
	.datac(!din_a[279]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_384 ),
	.cout(Xd_0__inst_mult_23_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_119 (
// Equation(s):

	.dataa(!din_a[277]),
	.datab(!din_b[278]),
	.datac(!din_a[276]),
	.datad(!din_b[279]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_389 ),
	.cout(Xd_0__inst_mult_23_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_118 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[265]),
	.datac(!din_a[267]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_384 ),
	.cout(Xd_0__inst_mult_22_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_119 (
// Equation(s):

	.dataa(!din_a[265]),
	.datab(!din_b[266]),
	.datac(!din_a[264]),
	.datad(!din_b[267]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_389 ),
	.cout(Xd_0__inst_mult_22_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_118 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[205]),
	.datac(!din_a[207]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_384 ),
	.cout(Xd_0__inst_mult_17_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_119 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[206]),
	.datac(!din_a[204]),
	.datad(!din_b[207]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_389 ),
	.cout(Xd_0__inst_mult_17_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_118 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[193]),
	.datac(!din_a[195]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_384 ),
	.cout(Xd_0__inst_mult_16_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_119 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[194]),
	.datac(!din_a[192]),
	.datad(!din_b[195]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_389 ),
	.cout(Xd_0__inst_mult_16_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_118 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[229]),
	.datac(!din_a[231]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_384 ),
	.cout(Xd_0__inst_mult_19_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_119 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[230]),
	.datac(!din_a[228]),
	.datad(!din_b[231]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_389 ),
	.cout(Xd_0__inst_mult_19_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_105 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[217]),
	.datac(!din_a[219]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_319 ),
	.cout(Xd_0__inst_mult_18_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_106 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[218]),
	.datac(!din_a[216]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_324 ),
	.cout(Xd_0__inst_mult_18_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_110 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[157]),
	.datac(!din_a[159]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_344 ),
	.cout(Xd_0__inst_mult_13_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_111 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[158]),
	.datac(!din_a[156]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_349 ),
	.cout(Xd_0__inst_mult_13_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_105 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[145]),
	.datac(!din_a[147]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_319 ),
	.cout(Xd_0__inst_mult_12_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_106 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[146]),
	.datac(!din_a[144]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_324 ),
	.cout(Xd_0__inst_mult_12_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_105 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[181]),
	.datac(!din_a[183]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_319 ),
	.cout(Xd_0__inst_mult_15_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_106 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[182]),
	.datac(!din_a[180]),
	.datad(!din_b[183]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_324 ),
	.cout(Xd_0__inst_mult_15_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_105 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[169]),
	.datac(!din_a[171]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_310 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_319 ),
	.cout(Xd_0__inst_mult_14_320 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_106 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[170]),
	.datac(!din_a[168]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_324 ),
	.cout(Xd_0__inst_mult_14_325 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_110 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[109]),
	.datac(!din_a[111]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_344 ),
	.cout(Xd_0__inst_mult_9_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_111 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[110]),
	.datac(!din_a[108]),
	.datad(!din_b[111]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_349 ),
	.cout(Xd_0__inst_mult_9_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_110 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[97]),
	.datac(!din_a[99]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_344 ),
	.cout(Xd_0__inst_mult_8_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_111 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[98]),
	.datac(!din_a[96]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_349 ),
	.cout(Xd_0__inst_mult_8_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_110 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[133]),
	.datac(!din_a[135]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_344 ),
	.cout(Xd_0__inst_mult_11_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_111 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[134]),
	.datac(!din_a[132]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_349 ),
	.cout(Xd_0__inst_mult_11_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_110 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[121]),
	.datac(!din_a[123]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_344 ),
	.cout(Xd_0__inst_mult_10_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_111 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[122]),
	.datac(!din_a[120]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_349 ),
	.cout(Xd_0__inst_mult_10_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_110 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[61]),
	.datac(!din_a[63]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_344 ),
	.cout(Xd_0__inst_mult_5_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_111 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[62]),
	.datac(!din_a[60]),
	.datad(!din_b[63]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_349 ),
	.cout(Xd_0__inst_mult_5_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_110 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[49]),
	.datac(!din_a[51]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_344 ),
	.cout(Xd_0__inst_mult_4_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_111 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[50]),
	.datac(!din_a[48]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_349 ),
	.cout(Xd_0__inst_mult_4_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_110 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[85]),
	.datac(!din_a[87]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_344 ),
	.cout(Xd_0__inst_mult_7_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_111 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[86]),
	.datac(!din_a[84]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_349 ),
	.cout(Xd_0__inst_mult_7_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_110 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[73]),
	.datac(!din_a[75]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_344 ),
	.cout(Xd_0__inst_mult_6_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_111 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[74]),
	.datac(!din_a[72]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_349 ),
	.cout(Xd_0__inst_mult_6_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_110 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[13]),
	.datac(!din_a[15]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_344 ),
	.cout(Xd_0__inst_mult_1_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_111 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[14]),
	.datac(!din_a[12]),
	.datad(!din_b[15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_349 ),
	.cout(Xd_0__inst_mult_1_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_110 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[1]),
	.datac(!din_a[3]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_344 ),
	.cout(Xd_0__inst_mult_0_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_111 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[2]),
	.datac(!din_a[0]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_349 ),
	.cout(Xd_0__inst_mult_0_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_110 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[37]),
	.datac(!din_a[39]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_344 ),
	.cout(Xd_0__inst_mult_3_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_111 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[38]),
	.datac(!din_a[36]),
	.datad(!din_b[39]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_349 ),
	.cout(Xd_0__inst_mult_3_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_122 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[25]),
	.datac(!din_a[27]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_404 ),
	.cout(Xd_0__inst_mult_2_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_123 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[26]),
	.datac(!din_a[24]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_409 ),
	.cout(Xd_0__inst_mult_2_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_120 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[349]),
	.datac(!din_a[352]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_394 ),
	.cout(Xd_0__inst_mult_29_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_121 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[350]),
	.datac(!din_a[348]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_399 ),
	.cout(Xd_0__inst_mult_29_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_112 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[337]),
	.datac(!din_a[340]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_354 ),
	.cout(Xd_0__inst_mult_28_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_113 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[338]),
	.datac(!din_a[336]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_359 ),
	.cout(Xd_0__inst_mult_28_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_112 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[373]),
	.datac(!din_a[376]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_354 ),
	.cout(Xd_0__inst_mult_31_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_113 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[374]),
	.datac(!din_a[372]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_359 ),
	.cout(Xd_0__inst_mult_31_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_112 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[361]),
	.datac(!din_a[364]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_354 ),
	.cout(Xd_0__inst_mult_30_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_113 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[362]),
	.datac(!din_a[360]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_359 ),
	.cout(Xd_0__inst_mult_30_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_132 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[301]),
	.datac(!din_a[304]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_454 ),
	.cout(Xd_0__inst_mult_25_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_133 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[302]),
	.datac(!din_a[300]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_459 ),
	.cout(Xd_0__inst_mult_25_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_170 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[289]),
	.datac(!din_a[292]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_644 ),
	.cout(Xd_0__inst_mult_24_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_171 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[290]),
	.datac(!din_a[288]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_649 ),
	.cout(Xd_0__inst_mult_24_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_132 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[325]),
	.datac(!din_a[328]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_454 ),
	.cout(Xd_0__inst_mult_27_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_133 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[326]),
	.datac(!din_a[324]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_459 ),
	.cout(Xd_0__inst_mult_27_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_170 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[313]),
	.datac(!din_a[316]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_644 ),
	.cout(Xd_0__inst_mult_26_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_171 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[314]),
	.datac(!din_a[312]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_649 ),
	.cout(Xd_0__inst_mult_26_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_120 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[253]),
	.datac(!din_a[256]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_394 ),
	.cout(Xd_0__inst_mult_21_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_121 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[254]),
	.datac(!din_a[252]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_399 ),
	.cout(Xd_0__inst_mult_21_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_120 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[241]),
	.datac(!din_a[244]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_394 ),
	.cout(Xd_0__inst_mult_20_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_121 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[242]),
	.datac(!din_a[240]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_399 ),
	.cout(Xd_0__inst_mult_20_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_120 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[277]),
	.datac(!din_a[280]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_394 ),
	.cout(Xd_0__inst_mult_23_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_121 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[278]),
	.datac(!din_a[276]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_399 ),
	.cout(Xd_0__inst_mult_23_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_120 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[265]),
	.datac(!din_a[268]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_394 ),
	.cout(Xd_0__inst_mult_22_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_121 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[266]),
	.datac(!din_a[264]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_399 ),
	.cout(Xd_0__inst_mult_22_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_120 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[205]),
	.datac(!din_a[208]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_394 ),
	.cout(Xd_0__inst_mult_17_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_121 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[206]),
	.datac(!din_a[204]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_399 ),
	.cout(Xd_0__inst_mult_17_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_120 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[193]),
	.datac(!din_a[196]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_394 ),
	.cout(Xd_0__inst_mult_16_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_121 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[194]),
	.datac(!din_a[192]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_399 ),
	.cout(Xd_0__inst_mult_16_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_120 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[229]),
	.datac(!din_a[232]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_394 ),
	.cout(Xd_0__inst_mult_19_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_121 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[230]),
	.datac(!din_a[228]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_399 ),
	.cout(Xd_0__inst_mult_19_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_107 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[217]),
	.datac(!din_a[220]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_329 ),
	.cout(Xd_0__inst_mult_18_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_108 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[218]),
	.datac(!din_a[216]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_334 ),
	.cout(Xd_0__inst_mult_18_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_112 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[157]),
	.datac(!din_a[160]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_354 ),
	.cout(Xd_0__inst_mult_13_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_113 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[158]),
	.datac(!din_a[156]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_359 ),
	.cout(Xd_0__inst_mult_13_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_107 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[145]),
	.datac(!din_a[148]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_329 ),
	.cout(Xd_0__inst_mult_12_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_108 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[146]),
	.datac(!din_a[144]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_334 ),
	.cout(Xd_0__inst_mult_12_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_107 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[181]),
	.datac(!din_a[184]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_329 ),
	.cout(Xd_0__inst_mult_15_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_108 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[182]),
	.datac(!din_a[180]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_334 ),
	.cout(Xd_0__inst_mult_15_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_107 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[169]),
	.datac(!din_a[172]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_329 ),
	.cout(Xd_0__inst_mult_14_330 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_108 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[170]),
	.datac(!din_a[168]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_315 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_334 ),
	.cout(Xd_0__inst_mult_14_335 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_112 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[109]),
	.datac(!din_a[112]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_354 ),
	.cout(Xd_0__inst_mult_9_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_113 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[110]),
	.datac(!din_a[108]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_359 ),
	.cout(Xd_0__inst_mult_9_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_112 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[97]),
	.datac(!din_a[100]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_354 ),
	.cout(Xd_0__inst_mult_8_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_113 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[98]),
	.datac(!din_a[96]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_359 ),
	.cout(Xd_0__inst_mult_8_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_112 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[133]),
	.datac(!din_a[136]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_354 ),
	.cout(Xd_0__inst_mult_11_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_113 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[134]),
	.datac(!din_a[132]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_359 ),
	.cout(Xd_0__inst_mult_11_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_112 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[121]),
	.datac(!din_a[124]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_354 ),
	.cout(Xd_0__inst_mult_10_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_113 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[122]),
	.datac(!din_a[120]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_359 ),
	.cout(Xd_0__inst_mult_10_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_112 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[61]),
	.datac(!din_a[64]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_354 ),
	.cout(Xd_0__inst_mult_5_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_113 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[62]),
	.datac(!din_a[60]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_359 ),
	.cout(Xd_0__inst_mult_5_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_112 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(!din_a[52]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_354 ),
	.cout(Xd_0__inst_mult_4_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_113 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[50]),
	.datac(!din_a[48]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_359 ),
	.cout(Xd_0__inst_mult_4_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_112 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(!din_a[88]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_354 ),
	.cout(Xd_0__inst_mult_7_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_113 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[86]),
	.datac(!din_a[84]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_359 ),
	.cout(Xd_0__inst_mult_7_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_112 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(!din_a[76]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_354 ),
	.cout(Xd_0__inst_mult_6_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_113 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[74]),
	.datac(!din_a[72]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_359 ),
	.cout(Xd_0__inst_mult_6_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_112 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[13]),
	.datac(!din_a[16]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_354 ),
	.cout(Xd_0__inst_mult_1_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_113 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[14]),
	.datac(!din_a[12]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_359 ),
	.cout(Xd_0__inst_mult_1_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_112 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(!din_a[4]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_354 ),
	.cout(Xd_0__inst_mult_0_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_113 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[2]),
	.datac(!din_a[0]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_359 ),
	.cout(Xd_0__inst_mult_0_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_112 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[37]),
	.datac(!din_a[40]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_354 ),
	.cout(Xd_0__inst_mult_3_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_113 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[38]),
	.datac(!din_a[36]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_359 ),
	.cout(Xd_0__inst_mult_3_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_124 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(!din_a[28]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_414 ),
	.cout(Xd_0__inst_mult_2_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_125 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[26]),
	.datac(!din_a[24]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_419 ),
	.cout(Xd_0__inst_mult_2_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_529 ),
	.datab(!Xd_0__inst_mult_29_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_404 ),
	.cout(Xd_0__inst_mult_29_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_29_123 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[353]),
	.datac(!din_a[349]),
	.datad(!din_b[354]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_409 ),
	.cout(Xd_0__inst_mult_29_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_50 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[238]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_50_sumout ),
	.cout(Xd_0__inst_mult_19_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_499 ),
	.datab(!Xd_0__inst_mult_28_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_364 ),
	.cout(Xd_0__inst_mult_28_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_28_115 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[341]),
	.datac(!din_a[337]),
	.datad(!din_b[342]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_369 ),
	.cout(Xd_0__inst_mult_28_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_50 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[274]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_50_sumout ),
	.cout(Xd_0__inst_mult_22_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_499 ),
	.datab(!Xd_0__inst_mult_31_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_364 ),
	.cout(Xd_0__inst_mult_31_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_31_115 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[377]),
	.datac(!din_a[373]),
	.datad(!din_b[378]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_369 ),
	.cout(Xd_0__inst_mult_31_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_50 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[262]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_50_sumout ),
	.cout(Xd_0__inst_mult_21_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_499 ),
	.datab(!Xd_0__inst_mult_30_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_364 ),
	.cout(Xd_0__inst_mult_30_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_30_115 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[365]),
	.datac(!din_a[361]),
	.datad(!din_b[366]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_369 ),
	.cout(Xd_0__inst_mult_30_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_60 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[250]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_60_sumout ),
	.cout(Xd_0__inst_mult_20_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_574 ),
	.datab(!Xd_0__inst_mult_25_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_464 ),
	.cout(Xd_0__inst_mult_25_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_25_135 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[305]),
	.datac(!din_a[301]),
	.datad(!din_b[306]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_469 ),
	.cout(Xd_0__inst_mult_25_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_172 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_729 ),
	.datab(!Xd_0__inst_mult_24_734 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_654 ),
	.cout(Xd_0__inst_mult_24_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_24_173 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[293]),
	.datac(!din_a[289]),
	.datad(!din_b[294]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_659 ),
	.cout(Xd_0__inst_mult_24_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_50 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[370]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_50_sumout ),
	.cout(Xd_0__inst_mult_30_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_574 ),
	.datab(!Xd_0__inst_mult_27_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_464 ),
	.cout(Xd_0__inst_mult_27_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_27_135 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[329]),
	.datac(!din_a[325]),
	.datad(!din_b[330]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_469 ),
	.cout(Xd_0__inst_mult_27_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_50 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[358]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_50_sumout ),
	.cout(Xd_0__inst_mult_29_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_172 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_729 ),
	.datab(!Xd_0__inst_mult_26_734 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_654 ),
	.cout(Xd_0__inst_mult_26_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_26_173 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[317]),
	.datac(!din_a[313]),
	.datad(!din_b[318]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_659 ),
	.cout(Xd_0__inst_mult_26_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_50 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_50_sumout ),
	.cout(Xd_0__inst_mult_0_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_529 ),
	.datab(!Xd_0__inst_mult_21_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_404 ),
	.cout(Xd_0__inst_mult_21_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_21_123 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[257]),
	.datac(!din_a[253]),
	.datad(!din_b[258]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_409 ),
	.cout(Xd_0__inst_mult_21_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_50 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_50_sumout ),
	.cout(Xd_0__inst_mult_7_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_529 ),
	.datab(!Xd_0__inst_mult_20_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_404 ),
	.cout(Xd_0__inst_mult_20_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_20_123 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[245]),
	.datac(!din_a[241]),
	.datad(!din_b[246]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_409 ),
	.cout(Xd_0__inst_mult_20_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_50 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_50_sumout ),
	.cout(Xd_0__inst_mult_9_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_529 ),
	.datab(!Xd_0__inst_mult_23_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_404 ),
	.cout(Xd_0__inst_mult_23_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_23_123 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[281]),
	.datac(!din_a[277]),
	.datad(!din_b[282]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_409 ),
	.cout(Xd_0__inst_mult_23_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_65 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_65_sumout ),
	.cout(Xd_0__inst_mult_8_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_529 ),
	.datab(!Xd_0__inst_mult_22_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_404 ),
	.cout(Xd_0__inst_mult_22_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_22_123 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[269]),
	.datac(!din_a[265]),
	.datad(!din_b[270]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_409 ),
	.cout(Xd_0__inst_mult_22_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_529 ),
	.datab(!Xd_0__inst_mult_17_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_404 ),
	.cout(Xd_0__inst_mult_17_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_17_123 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[209]),
	.datac(!din_a[205]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_409 ),
	.cout(Xd_0__inst_mult_17_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_50 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[129]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_50_sumout ),
	.cout(Xd_0__inst_mult_10_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_529 ),
	.datab(!Xd_0__inst_mult_16_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_404 ),
	.cout(Xd_0__inst_mult_16_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_16_123 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[197]),
	.datac(!din_a[193]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_409 ),
	.cout(Xd_0__inst_mult_16_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_65 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_65_sumout ),
	.cout(Xd_0__inst_mult_3_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_529 ),
	.datab(!Xd_0__inst_mult_19_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_404 ),
	.cout(Xd_0__inst_mult_19_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_19_123 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[233]),
	.datac(!din_a[229]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_409 ),
	.cout(Xd_0__inst_mult_19_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_60 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_60_sumout ),
	.cout(Xd_0__inst_mult_6_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_474 ),
	.datab(!Xd_0__inst_mult_18_479 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_339 ),
	.cout(Xd_0__inst_mult_18_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_18_110 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[221]),
	.datac(!din_a[217]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_344 ),
	.cout(Xd_0__inst_mult_18_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_499 ),
	.datab(!Xd_0__inst_mult_13_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_364 ),
	.cout(Xd_0__inst_mult_13_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_13_115 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[161]),
	.datac(!din_a[157]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_369 ),
	.cout(Xd_0__inst_mult_13_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_474 ),
	.datab(!Xd_0__inst_mult_12_479 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_339 ),
	.cout(Xd_0__inst_mult_12_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_12_110 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[149]),
	.datac(!din_a[145]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_344 ),
	.cout(Xd_0__inst_mult_12_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_474 ),
	.datab(!Xd_0__inst_mult_15_479 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_339 ),
	.cout(Xd_0__inst_mult_15_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_15_110 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[185]),
	.datac(!din_a[181]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_344 ),
	.cout(Xd_0__inst_mult_15_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_109 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_474 ),
	.datab(!Xd_0__inst_mult_14_479 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_305 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_339 ),
	.cout(Xd_0__inst_mult_14_340 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_14_110 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[173]),
	.datac(!din_a[169]),
	.datad(!din_b[174]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_344 ),
	.cout(Xd_0__inst_mult_14_345 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_499 ),
	.datab(!Xd_0__inst_mult_9_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_364 ),
	.cout(Xd_0__inst_mult_9_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_9_115 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[113]),
	.datac(!din_a[109]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_369 ),
	.cout(Xd_0__inst_mult_9_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_499 ),
	.datab(!Xd_0__inst_mult_8_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_364 ),
	.cout(Xd_0__inst_mult_8_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_8_115 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[101]),
	.datac(!din_a[97]),
	.datad(!din_b[102]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_369 ),
	.cout(Xd_0__inst_mult_8_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_499 ),
	.datab(!Xd_0__inst_mult_11_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_364 ),
	.cout(Xd_0__inst_mult_11_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_11_115 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[137]),
	.datac(!din_a[133]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_369 ),
	.cout(Xd_0__inst_mult_11_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_499 ),
	.datab(!Xd_0__inst_mult_10_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_364 ),
	.cout(Xd_0__inst_mult_10_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_10_115 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[125]),
	.datac(!din_a[121]),
	.datad(!din_b[126]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_369 ),
	.cout(Xd_0__inst_mult_10_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_55 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[370]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_55_sumout ),
	.cout(Xd_0__inst_mult_30_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_499 ),
	.datab(!Xd_0__inst_mult_5_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_364 ),
	.cout(Xd_0__inst_mult_5_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_5_115 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[65]),
	.datac(!din_a[61]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_369 ),
	.cout(Xd_0__inst_mult_5_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_55 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[358]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_55_sumout ),
	.cout(Xd_0__inst_mult_29_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_499 ),
	.datab(!Xd_0__inst_mult_4_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_364 ),
	.cout(Xd_0__inst_mult_4_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_4_115 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[53]),
	.datac(!din_a[49]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_369 ),
	.cout(Xd_0__inst_mult_4_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_55 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_55_sumout ),
	.cout(Xd_0__inst_mult_0_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_499 ),
	.datab(!Xd_0__inst_mult_7_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_364 ),
	.cout(Xd_0__inst_mult_7_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_7_115 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[89]),
	.datac(!din_a[85]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_369 ),
	.cout(Xd_0__inst_mult_7_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_55 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_55_sumout ),
	.cout(Xd_0__inst_mult_7_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_499 ),
	.datab(!Xd_0__inst_mult_6_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_364 ),
	.cout(Xd_0__inst_mult_6_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_6_115 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[77]),
	.datac(!din_a[73]),
	.datad(!din_b[78]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_369 ),
	.cout(Xd_0__inst_mult_6_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_55 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[129]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_55_sumout ),
	.cout(Xd_0__inst_mult_10_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_499 ),
	.datab(!Xd_0__inst_mult_1_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_364 ),
	.cout(Xd_0__inst_mult_1_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_1_115 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[17]),
	.datac(!din_a[13]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_369 ),
	.cout(Xd_0__inst_mult_1_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_55 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_55_sumout ),
	.cout(Xd_0__inst_mult_9_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_499 ),
	.datab(!Xd_0__inst_mult_0_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_364 ),
	.cout(Xd_0__inst_mult_0_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_0_115 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[5]),
	.datac(!din_a[1]),
	.datad(!din_b[6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_369 ),
	.cout(Xd_0__inst_mult_0_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_45 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[153]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_45_sumout ),
	.cout(Xd_0__inst_mult_12_46 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_114 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_499 ),
	.datab(!Xd_0__inst_mult_3_504 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_320 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_364 ),
	.cout(Xd_0__inst_mult_3_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_3_115 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[41]),
	.datac(!din_a[37]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_369 ),
	.cout(Xd_0__inst_mult_3_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_60 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_60_sumout ),
	.cout(Xd_0__inst_mult_7_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_544 ),
	.datab(!Xd_0__inst_mult_2_549 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_424 ),
	.cout(Xd_0__inst_mult_2_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_60 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_60_sumout ),
	.cout(Xd_0__inst_mult_10_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_539 ),
	.datab(!Xd_0__inst_mult_29_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_414 ),
	.cout(Xd_0__inst_mult_29_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_125 (
// Equation(s):

	.dataa(!din_a[349]),
	.datab(!din_b[353]),
	.datac(!din_a[348]),
	.datad(!din_b[354]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_419 ),
	.cout(Xd_0__inst_mult_29_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_509 ),
	.datab(!Xd_0__inst_mult_28_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_374 ),
	.cout(Xd_0__inst_mult_28_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_117 (
// Equation(s):

	.dataa(!din_a[337]),
	.datab(!din_b[341]),
	.datac(!din_a[336]),
	.datad(!din_b[342]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_379 ),
	.cout(Xd_0__inst_mult_28_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_509 ),
	.datab(!Xd_0__inst_mult_31_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_374 ),
	.cout(Xd_0__inst_mult_31_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_117 (
// Equation(s):

	.dataa(!din_a[373]),
	.datab(!din_b[377]),
	.datac(!din_a[372]),
	.datad(!din_b[378]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_379 ),
	.cout(Xd_0__inst_mult_31_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_509 ),
	.datab(!Xd_0__inst_mult_30_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_374 ),
	.cout(Xd_0__inst_mult_30_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_117 (
// Equation(s):

	.dataa(!din_a[361]),
	.datab(!din_b[365]),
	.datac(!din_a[360]),
	.datad(!din_b[366]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_379 ),
	.cout(Xd_0__inst_mult_30_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_584 ),
	.datab(!Xd_0__inst_mult_25_589 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_474 ),
	.cout(Xd_0__inst_mult_25_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_137 (
// Equation(s):

	.dataa(!din_a[301]),
	.datab(!din_b[305]),
	.datac(!din_a[300]),
	.datad(!din_b[306]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_479 ),
	.cout(Xd_0__inst_mult_25_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_174 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_739 ),
	.datab(!Xd_0__inst_mult_24_744 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_664 ),
	.cout(Xd_0__inst_mult_24_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_175 (
// Equation(s):

	.dataa(!din_a[289]),
	.datab(!din_b[293]),
	.datac(!din_a[288]),
	.datad(!din_b[294]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_669 ),
	.cout(Xd_0__inst_mult_24_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_584 ),
	.datab(!Xd_0__inst_mult_27_589 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_474 ),
	.cout(Xd_0__inst_mult_27_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_137 (
// Equation(s):

	.dataa(!din_a[325]),
	.datab(!din_b[329]),
	.datac(!din_a[324]),
	.datad(!din_b[330]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_479 ),
	.cout(Xd_0__inst_mult_27_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_174 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_739 ),
	.datab(!Xd_0__inst_mult_26_744 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_664 ),
	.cout(Xd_0__inst_mult_26_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_175 (
// Equation(s):

	.dataa(!din_a[313]),
	.datab(!din_b[317]),
	.datac(!din_a[312]),
	.datad(!din_b[318]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_669 ),
	.cout(Xd_0__inst_mult_26_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_539 ),
	.datab(!Xd_0__inst_mult_21_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_414 ),
	.cout(Xd_0__inst_mult_21_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_125 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[257]),
	.datac(!din_a[252]),
	.datad(!din_b[258]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_419 ),
	.cout(Xd_0__inst_mult_21_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_539 ),
	.datab(!Xd_0__inst_mult_20_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_414 ),
	.cout(Xd_0__inst_mult_20_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_125 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[245]),
	.datac(!din_a[240]),
	.datad(!din_b[246]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_419 ),
	.cout(Xd_0__inst_mult_20_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_539 ),
	.datab(!Xd_0__inst_mult_23_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_414 ),
	.cout(Xd_0__inst_mult_23_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_125 (
// Equation(s):

	.dataa(!din_a[277]),
	.datab(!din_b[281]),
	.datac(!din_a[276]),
	.datad(!din_b[282]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_419 ),
	.cout(Xd_0__inst_mult_23_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_539 ),
	.datab(!Xd_0__inst_mult_22_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_414 ),
	.cout(Xd_0__inst_mult_22_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_125 (
// Equation(s):

	.dataa(!din_a[265]),
	.datab(!din_b[269]),
	.datac(!din_a[264]),
	.datad(!din_b[270]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_419 ),
	.cout(Xd_0__inst_mult_22_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_539 ),
	.datab(!Xd_0__inst_mult_17_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_414 ),
	.cout(Xd_0__inst_mult_17_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_125 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[209]),
	.datac(!din_a[204]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_419 ),
	.cout(Xd_0__inst_mult_17_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_539 ),
	.datab(!Xd_0__inst_mult_16_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_414 ),
	.cout(Xd_0__inst_mult_16_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_125 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[197]),
	.datac(!din_a[192]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_419 ),
	.cout(Xd_0__inst_mult_16_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_539 ),
	.datab(!Xd_0__inst_mult_19_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_414 ),
	.cout(Xd_0__inst_mult_19_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_125 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[233]),
	.datac(!din_a[228]),
	.datad(!din_b[234]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_419 ),
	.cout(Xd_0__inst_mult_19_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_484 ),
	.datab(!Xd_0__inst_mult_18_489 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_349 ),
	.cout(Xd_0__inst_mult_18_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_112 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[221]),
	.datac(!din_a[216]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_354 ),
	.cout(Xd_0__inst_mult_18_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_509 ),
	.datab(!Xd_0__inst_mult_13_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_374 ),
	.cout(Xd_0__inst_mult_13_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_117 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[161]),
	.datac(!din_a[156]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_379 ),
	.cout(Xd_0__inst_mult_13_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_484 ),
	.datab(!Xd_0__inst_mult_12_489 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_349 ),
	.cout(Xd_0__inst_mult_12_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_112 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[149]),
	.datac(!din_a[144]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_354 ),
	.cout(Xd_0__inst_mult_12_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_484 ),
	.datab(!Xd_0__inst_mult_15_489 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_349 ),
	.cout(Xd_0__inst_mult_15_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_112 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[185]),
	.datac(!din_a[180]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_354 ),
	.cout(Xd_0__inst_mult_15_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_111 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_484 ),
	.datab(!Xd_0__inst_mult_14_489 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_340 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_349 ),
	.cout(Xd_0__inst_mult_14_350 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_112 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[173]),
	.datac(!din_a[168]),
	.datad(!din_b[174]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_354 ),
	.cout(Xd_0__inst_mult_14_355 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_509 ),
	.datab(!Xd_0__inst_mult_9_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_374 ),
	.cout(Xd_0__inst_mult_9_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_117 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[113]),
	.datac(!din_a[108]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_379 ),
	.cout(Xd_0__inst_mult_9_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_509 ),
	.datab(!Xd_0__inst_mult_8_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_374 ),
	.cout(Xd_0__inst_mult_8_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_117 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[101]),
	.datac(!din_a[96]),
	.datad(!din_b[102]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_379 ),
	.cout(Xd_0__inst_mult_8_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_509 ),
	.datab(!Xd_0__inst_mult_11_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_374 ),
	.cout(Xd_0__inst_mult_11_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_117 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[137]),
	.datac(!din_a[132]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_379 ),
	.cout(Xd_0__inst_mult_11_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_509 ),
	.datab(!Xd_0__inst_mult_10_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_374 ),
	.cout(Xd_0__inst_mult_10_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_117 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[125]),
	.datac(!din_a[120]),
	.datad(!din_b[126]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_379 ),
	.cout(Xd_0__inst_mult_10_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_509 ),
	.datab(!Xd_0__inst_mult_5_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_374 ),
	.cout(Xd_0__inst_mult_5_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_117 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[65]),
	.datac(!din_a[60]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_379 ),
	.cout(Xd_0__inst_mult_5_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_509 ),
	.datab(!Xd_0__inst_mult_4_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_374 ),
	.cout(Xd_0__inst_mult_4_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_117 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[53]),
	.datac(!din_a[48]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_379 ),
	.cout(Xd_0__inst_mult_4_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_509 ),
	.datab(!Xd_0__inst_mult_7_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_374 ),
	.cout(Xd_0__inst_mult_7_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_117 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[89]),
	.datac(!din_a[84]),
	.datad(!din_b[90]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_379 ),
	.cout(Xd_0__inst_mult_7_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_509 ),
	.datab(!Xd_0__inst_mult_6_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_374 ),
	.cout(Xd_0__inst_mult_6_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_117 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[77]),
	.datac(!din_a[72]),
	.datad(!din_b[78]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_379 ),
	.cout(Xd_0__inst_mult_6_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_509 ),
	.datab(!Xd_0__inst_mult_1_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_374 ),
	.cout(Xd_0__inst_mult_1_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_117 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[17]),
	.datac(!din_a[12]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_379 ),
	.cout(Xd_0__inst_mult_1_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_509 ),
	.datab(!Xd_0__inst_mult_0_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_374 ),
	.cout(Xd_0__inst_mult_0_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_117 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[5]),
	.datac(!din_a[0]),
	.datad(!din_b[6]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_379 ),
	.cout(Xd_0__inst_mult_0_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_509 ),
	.datab(!Xd_0__inst_mult_3_514 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_374 ),
	.cout(Xd_0__inst_mult_3_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_117 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[41]),
	.datac(!din_a[36]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_379 ),
	.cout(Xd_0__inst_mult_3_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_554 ),
	.datab(!Xd_0__inst_mult_2_559 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_429 ),
	.cout(Xd_0__inst_mult_2_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_549 ),
	.datab(!Xd_0__inst_mult_29_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_424 ),
	.cout(Xd_0__inst_mult_29_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_127 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[353]),
	.datac(!din_a[348]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_429 ),
	.cout(Xd_0__inst_mult_29_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_519 ),
	.datab(!Xd_0__inst_mult_28_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_384 ),
	.cout(Xd_0__inst_mult_28_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_119 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[341]),
	.datac(!din_a[336]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_389 ),
	.cout(Xd_0__inst_mult_28_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_519 ),
	.datab(!Xd_0__inst_mult_31_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_384 ),
	.cout(Xd_0__inst_mult_31_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_119 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[377]),
	.datac(!din_a[372]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_389 ),
	.cout(Xd_0__inst_mult_31_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_519 ),
	.datab(!Xd_0__inst_mult_30_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_384 ),
	.cout(Xd_0__inst_mult_30_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_119 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[365]),
	.datac(!din_a[360]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_389 ),
	.cout(Xd_0__inst_mult_30_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_569 ),
	.datab(!Xd_0__inst_mult_25_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_484 ),
	.cout(Xd_0__inst_mult_25_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_139 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[305]),
	.datac(!din_a[300]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_489 ),
	.cout(Xd_0__inst_mult_25_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_176 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_709 ),
	.datab(!Xd_0__inst_mult_24_704 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_674 ),
	.cout(Xd_0__inst_mult_24_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_177 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[293]),
	.datac(!din_a[288]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_679 ),
	.cout(Xd_0__inst_mult_24_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_569 ),
	.datab(!Xd_0__inst_mult_27_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_484 ),
	.cout(Xd_0__inst_mult_27_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_139 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[329]),
	.datac(!din_a[324]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_489 ),
	.cout(Xd_0__inst_mult_27_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_176 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_724 ),
	.datab(!Xd_0__inst_mult_26_719 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_674 ),
	.cout(Xd_0__inst_mult_26_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_177 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[317]),
	.datac(!din_a[312]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_679 ),
	.cout(Xd_0__inst_mult_26_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_549 ),
	.datab(!Xd_0__inst_mult_21_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_424 ),
	.cout(Xd_0__inst_mult_21_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_127 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[257]),
	.datac(!din_a[252]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_429 ),
	.cout(Xd_0__inst_mult_21_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_549 ),
	.datab(!Xd_0__inst_mult_20_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_424 ),
	.cout(Xd_0__inst_mult_20_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_127 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[245]),
	.datac(!din_a[240]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_429 ),
	.cout(Xd_0__inst_mult_20_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_549 ),
	.datab(!Xd_0__inst_mult_23_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_424 ),
	.cout(Xd_0__inst_mult_23_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_127 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[281]),
	.datac(!din_a[276]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_429 ),
	.cout(Xd_0__inst_mult_23_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_549 ),
	.datab(!Xd_0__inst_mult_22_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_424 ),
	.cout(Xd_0__inst_mult_22_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_127 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[269]),
	.datac(!din_a[264]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_429 ),
	.cout(Xd_0__inst_mult_22_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_549 ),
	.datab(!Xd_0__inst_mult_17_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_424 ),
	.cout(Xd_0__inst_mult_17_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_127 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[209]),
	.datac(!din_a[204]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_429 ),
	.cout(Xd_0__inst_mult_17_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_549 ),
	.datab(!Xd_0__inst_mult_16_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_424 ),
	.cout(Xd_0__inst_mult_16_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_127 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[197]),
	.datac(!din_a[192]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_429 ),
	.cout(Xd_0__inst_mult_16_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_549 ),
	.datab(!Xd_0__inst_mult_19_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_424 ),
	.cout(Xd_0__inst_mult_19_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_127 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[233]),
	.datac(!din_a[228]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_429 ),
	.cout(Xd_0__inst_mult_19_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_494 ),
	.datab(!Xd_0__inst_mult_18_499 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_359 ),
	.cout(Xd_0__inst_mult_18_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_114 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[221]),
	.datac(!din_a[216]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_364 ),
	.cout(Xd_0__inst_mult_18_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_519 ),
	.datab(!Xd_0__inst_mult_13_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_384 ),
	.cout(Xd_0__inst_mult_13_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_119 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[161]),
	.datac(!din_a[156]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_389 ),
	.cout(Xd_0__inst_mult_13_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_494 ),
	.datab(!Xd_0__inst_mult_12_499 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_359 ),
	.cout(Xd_0__inst_mult_12_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_114 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[149]),
	.datac(!din_a[144]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_364 ),
	.cout(Xd_0__inst_mult_12_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_494 ),
	.datab(!Xd_0__inst_mult_15_499 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_359 ),
	.cout(Xd_0__inst_mult_15_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_114 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[185]),
	.datac(!din_a[180]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_364 ),
	.cout(Xd_0__inst_mult_15_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_113 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_494 ),
	.datab(!Xd_0__inst_mult_14_499 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_350 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_359 ),
	.cout(Xd_0__inst_mult_14_360 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_114 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[173]),
	.datac(!din_a[168]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_345 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_364 ),
	.cout(Xd_0__inst_mult_14_365 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_519 ),
	.datab(!Xd_0__inst_mult_9_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_384 ),
	.cout(Xd_0__inst_mult_9_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_119 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[113]),
	.datac(!din_a[108]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_389 ),
	.cout(Xd_0__inst_mult_9_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_519 ),
	.datab(!Xd_0__inst_mult_8_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_384 ),
	.cout(Xd_0__inst_mult_8_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_119 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[101]),
	.datac(!din_a[96]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_389 ),
	.cout(Xd_0__inst_mult_8_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_519 ),
	.datab(!Xd_0__inst_mult_11_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_384 ),
	.cout(Xd_0__inst_mult_11_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_119 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[137]),
	.datac(!din_a[132]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_389 ),
	.cout(Xd_0__inst_mult_11_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_519 ),
	.datab(!Xd_0__inst_mult_10_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_384 ),
	.cout(Xd_0__inst_mult_10_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_119 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[125]),
	.datac(!din_a[120]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_389 ),
	.cout(Xd_0__inst_mult_10_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_519 ),
	.datab(!Xd_0__inst_mult_5_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_384 ),
	.cout(Xd_0__inst_mult_5_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_119 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[65]),
	.datac(!din_a[60]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_389 ),
	.cout(Xd_0__inst_mult_5_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_519 ),
	.datab(!Xd_0__inst_mult_4_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_384 ),
	.cout(Xd_0__inst_mult_4_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_119 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[53]),
	.datac(!din_a[48]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_389 ),
	.cout(Xd_0__inst_mult_4_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_519 ),
	.datab(!Xd_0__inst_mult_7_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_384 ),
	.cout(Xd_0__inst_mult_7_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_119 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[89]),
	.datac(!din_a[84]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_389 ),
	.cout(Xd_0__inst_mult_7_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_519 ),
	.datab(!Xd_0__inst_mult_6_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_384 ),
	.cout(Xd_0__inst_mult_6_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_119 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[77]),
	.datac(!din_a[72]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_389 ),
	.cout(Xd_0__inst_mult_6_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_519 ),
	.datab(!Xd_0__inst_mult_1_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_384 ),
	.cout(Xd_0__inst_mult_1_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_119 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[17]),
	.datac(!din_a[12]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_389 ),
	.cout(Xd_0__inst_mult_1_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_519 ),
	.datab(!Xd_0__inst_mult_0_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_384 ),
	.cout(Xd_0__inst_mult_0_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_119 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[5]),
	.datac(!din_a[0]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_389 ),
	.cout(Xd_0__inst_mult_0_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_519 ),
	.datab(!Xd_0__inst_mult_3_524 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_384 ),
	.cout(Xd_0__inst_mult_3_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_119 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[41]),
	.datac(!din_a[36]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_389 ),
	.cout(Xd_0__inst_mult_3_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_564 ),
	.datab(!Xd_0__inst_mult_2_569 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_434 ),
	.cout(Xd_0__inst_mult_2_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_559 ),
	.datab(!Xd_0__inst_mult_29_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_434 ),
	.cout(Xd_0__inst_mult_29_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_569 ),
	.datab(!Xd_0__inst_mult_29_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_439 ),
	.cout(Xd_0__inst_mult_29_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_529 ),
	.datab(!Xd_0__inst_mult_28_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_394 ),
	.cout(Xd_0__inst_mult_28_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_539 ),
	.datab(!Xd_0__inst_mult_28_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_399 ),
	.cout(Xd_0__inst_mult_28_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_529 ),
	.datab(!Xd_0__inst_mult_31_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_394 ),
	.cout(Xd_0__inst_mult_31_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_539 ),
	.datab(!Xd_0__inst_mult_31_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_399 ),
	.cout(Xd_0__inst_mult_31_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_529 ),
	.datab(!Xd_0__inst_mult_30_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_394 ),
	.cout(Xd_0__inst_mult_30_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_539 ),
	.datab(!Xd_0__inst_mult_30_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_399 ),
	.cout(Xd_0__inst_mult_30_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_594 ),
	.datab(!Xd_0__inst_mult_25_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_494 ),
	.cout(Xd_0__inst_mult_25_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_178 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_749 ),
	.datab(!Xd_0__inst_mult_24_754 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_684 ),
	.cout(Xd_0__inst_mult_24_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_594 ),
	.datab(!Xd_0__inst_mult_27_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_102 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_494 ),
	.cout(Xd_0__inst_mult_27_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_178 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_749 ),
	.datab(!Xd_0__inst_mult_26_754 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_684 ),
	.cout(Xd_0__inst_mult_26_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_559 ),
	.datab(!Xd_0__inst_mult_21_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_434 ),
	.cout(Xd_0__inst_mult_21_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_569 ),
	.datab(!Xd_0__inst_mult_21_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_117 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_439 ),
	.cout(Xd_0__inst_mult_21_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_559 ),
	.datab(!Xd_0__inst_mult_20_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_434 ),
	.cout(Xd_0__inst_mult_20_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_569 ),
	.datab(!Xd_0__inst_mult_20_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_152 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_439 ),
	.cout(Xd_0__inst_mult_20_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_559 ),
	.datab(!Xd_0__inst_mult_23_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_434 ),
	.cout(Xd_0__inst_mult_23_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_569 ),
	.datab(!Xd_0__inst_mult_23_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_439 ),
	.cout(Xd_0__inst_mult_23_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_559 ),
	.datab(!Xd_0__inst_mult_22_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_434 ),
	.cout(Xd_0__inst_mult_22_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_569 ),
	.datab(!Xd_0__inst_mult_22_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_2 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_439 ),
	.cout(Xd_0__inst_mult_22_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_559 ),
	.datab(!Xd_0__inst_mult_17_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_434 ),
	.cout(Xd_0__inst_mult_17_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_569 ),
	.datab(!Xd_0__inst_mult_17_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_37 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_439 ),
	.cout(Xd_0__inst_mult_17_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_559 ),
	.datab(!Xd_0__inst_mult_16_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_434 ),
	.cout(Xd_0__inst_mult_16_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_569 ),
	.datab(!Xd_0__inst_mult_16_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_439 ),
	.cout(Xd_0__inst_mult_16_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_559 ),
	.datab(!Xd_0__inst_mult_19_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_434 ),
	.cout(Xd_0__inst_mult_19_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_569 ),
	.datab(!Xd_0__inst_mult_19_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_439 ),
	.cout(Xd_0__inst_mult_19_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_504 ),
	.datab(!Xd_0__inst_mult_18_509 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_369 ),
	.cout(Xd_0__inst_mult_18_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_514 ),
	.datab(!Xd_0__inst_mult_18_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_374 ),
	.cout(Xd_0__inst_mult_18_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_529 ),
	.datab(!Xd_0__inst_mult_13_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_394 ),
	.cout(Xd_0__inst_mult_13_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_539 ),
	.datab(!Xd_0__inst_mult_13_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_399 ),
	.cout(Xd_0__inst_mult_13_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_504 ),
	.datab(!Xd_0__inst_mult_12_509 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_369 ),
	.cout(Xd_0__inst_mult_12_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_514 ),
	.datab(!Xd_0__inst_mult_12_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_82 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_374 ),
	.cout(Xd_0__inst_mult_12_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_504 ),
	.datab(!Xd_0__inst_mult_15_509 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_369 ),
	.cout(Xd_0__inst_mult_15_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_514 ),
	.datab(!Xd_0__inst_mult_15_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_374 ),
	.cout(Xd_0__inst_mult_15_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_115 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_504 ),
	.datab(!Xd_0__inst_mult_14_509 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_369 ),
	.cout(Xd_0__inst_mult_14_370 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_116 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_514 ),
	.datab(!Xd_0__inst_mult_14_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_374 ),
	.cout(Xd_0__inst_mult_14_375 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_529 ),
	.datab(!Xd_0__inst_mult_9_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_394 ),
	.cout(Xd_0__inst_mult_9_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_539 ),
	.datab(!Xd_0__inst_mult_9_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_399 ),
	.cout(Xd_0__inst_mult_9_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_529 ),
	.datab(!Xd_0__inst_mult_8_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_394 ),
	.cout(Xd_0__inst_mult_8_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_539 ),
	.datab(!Xd_0__inst_mult_8_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_399 ),
	.cout(Xd_0__inst_mult_8_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_529 ),
	.datab(!Xd_0__inst_mult_11_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_394 ),
	.cout(Xd_0__inst_mult_11_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_539 ),
	.datab(!Xd_0__inst_mult_11_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_399 ),
	.cout(Xd_0__inst_mult_11_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_529 ),
	.datab(!Xd_0__inst_mult_10_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_394 ),
	.cout(Xd_0__inst_mult_10_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_539 ),
	.datab(!Xd_0__inst_mult_10_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_399 ),
	.cout(Xd_0__inst_mult_10_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_529 ),
	.datab(!Xd_0__inst_mult_5_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_394 ),
	.cout(Xd_0__inst_mult_5_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_539 ),
	.datab(!Xd_0__inst_mult_5_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_399 ),
	.cout(Xd_0__inst_mult_5_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_529 ),
	.datab(!Xd_0__inst_mult_4_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_394 ),
	.cout(Xd_0__inst_mult_4_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_539 ),
	.datab(!Xd_0__inst_mult_4_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_399 ),
	.cout(Xd_0__inst_mult_4_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_529 ),
	.datab(!Xd_0__inst_mult_7_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_394 ),
	.cout(Xd_0__inst_mult_7_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_539 ),
	.datab(!Xd_0__inst_mult_7_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_399 ),
	.cout(Xd_0__inst_mult_7_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_529 ),
	.datab(!Xd_0__inst_mult_6_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_394 ),
	.cout(Xd_0__inst_mult_6_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_539 ),
	.datab(!Xd_0__inst_mult_6_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_399 ),
	.cout(Xd_0__inst_mult_6_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_529 ),
	.datab(!Xd_0__inst_mult_1_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_394 ),
	.cout(Xd_0__inst_mult_1_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_539 ),
	.datab(!Xd_0__inst_mult_1_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_399 ),
	.cout(Xd_0__inst_mult_1_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_529 ),
	.datab(!Xd_0__inst_mult_0_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_394 ),
	.cout(Xd_0__inst_mult_0_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_539 ),
	.datab(!Xd_0__inst_mult_0_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_399 ),
	.cout(Xd_0__inst_mult_0_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_529 ),
	.datab(!Xd_0__inst_mult_3_534 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_394 ),
	.cout(Xd_0__inst_mult_3_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_539 ),
	.datab(!Xd_0__inst_mult_3_544 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_399 ),
	.cout(Xd_0__inst_mult_3_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_574 ),
	.datab(!Xd_0__inst_mult_2_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_439 ),
	.cout(Xd_0__inst_mult_2_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_584 ),
	.datab(!Xd_0__inst_mult_2_589 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_444 ),
	.cout(Xd_0__inst_mult_2_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_579 ),
	.datab(!Xd_0__inst_mult_29_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_444 ),
	.cout(Xd_0__inst_mult_29_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_589 ),
	.datab(!Xd_0__inst_mult_29_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_449 ),
	.cout(Xd_0__inst_mult_29_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_549 ),
	.datab(!Xd_0__inst_mult_28_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_404 ),
	.cout(Xd_0__inst_mult_28_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_559 ),
	.datab(!Xd_0__inst_mult_28_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_409 ),
	.cout(Xd_0__inst_mult_28_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_549 ),
	.datab(!Xd_0__inst_mult_31_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_404 ),
	.cout(Xd_0__inst_mult_31_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_559 ),
	.datab(!Xd_0__inst_mult_31_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_409 ),
	.cout(Xd_0__inst_mult_31_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_549 ),
	.datab(!Xd_0__inst_mult_30_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_404 ),
	.cout(Xd_0__inst_mult_30_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_559 ),
	.datab(!Xd_0__inst_mult_30_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_409 ),
	.cout(Xd_0__inst_mult_30_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_604 ),
	.datab(!Xd_0__inst_mult_25_609 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_499 ),
	.cout(Xd_0__inst_mult_25_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_179 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_759 ),
	.datab(!Xd_0__inst_mult_24_764 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_689 ),
	.cout(Xd_0__inst_mult_24_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_604 ),
	.datab(!Xd_0__inst_mult_27_609 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_499 ),
	.cout(Xd_0__inst_mult_27_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_179 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_759 ),
	.datab(!Xd_0__inst_mult_26_764 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_689 ),
	.cout(Xd_0__inst_mult_26_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_579 ),
	.datab(!Xd_0__inst_mult_21_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_444 ),
	.cout(Xd_0__inst_mult_21_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_589 ),
	.datab(!Xd_0__inst_mult_21_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_449 ),
	.cout(Xd_0__inst_mult_21_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_579 ),
	.datab(!Xd_0__inst_mult_20_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_444 ),
	.cout(Xd_0__inst_mult_20_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_589 ),
	.datab(!Xd_0__inst_mult_20_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_449 ),
	.cout(Xd_0__inst_mult_20_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_579 ),
	.datab(!Xd_0__inst_mult_23_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_444 ),
	.cout(Xd_0__inst_mult_23_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_589 ),
	.datab(!Xd_0__inst_mult_23_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_449 ),
	.cout(Xd_0__inst_mult_23_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_579 ),
	.datab(!Xd_0__inst_mult_22_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_444 ),
	.cout(Xd_0__inst_mult_22_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_589 ),
	.datab(!Xd_0__inst_mult_22_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_449 ),
	.cout(Xd_0__inst_mult_22_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_579 ),
	.datab(!Xd_0__inst_mult_17_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_444 ),
	.cout(Xd_0__inst_mult_17_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_589 ),
	.datab(!Xd_0__inst_mult_17_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_449 ),
	.cout(Xd_0__inst_mult_17_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_579 ),
	.datab(!Xd_0__inst_mult_16_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_444 ),
	.cout(Xd_0__inst_mult_16_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_589 ),
	.datab(!Xd_0__inst_mult_16_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_449 ),
	.cout(Xd_0__inst_mult_16_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_579 ),
	.datab(!Xd_0__inst_mult_19_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_444 ),
	.cout(Xd_0__inst_mult_19_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_589 ),
	.datab(!Xd_0__inst_mult_19_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_449 ),
	.cout(Xd_0__inst_mult_19_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_524 ),
	.datab(!Xd_0__inst_mult_18_529 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_379 ),
	.cout(Xd_0__inst_mult_18_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_534 ),
	.datab(!Xd_0__inst_mult_18_539 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_384 ),
	.cout(Xd_0__inst_mult_18_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_549 ),
	.datab(!Xd_0__inst_mult_13_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_404 ),
	.cout(Xd_0__inst_mult_13_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_559 ),
	.datab(!Xd_0__inst_mult_13_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_409 ),
	.cout(Xd_0__inst_mult_13_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_524 ),
	.datab(!Xd_0__inst_mult_12_529 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_379 ),
	.cout(Xd_0__inst_mult_12_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_534 ),
	.datab(!Xd_0__inst_mult_12_539 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_384 ),
	.cout(Xd_0__inst_mult_12_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_524 ),
	.datab(!Xd_0__inst_mult_15_529 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_379 ),
	.cout(Xd_0__inst_mult_15_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_534 ),
	.datab(!Xd_0__inst_mult_15_539 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_384 ),
	.cout(Xd_0__inst_mult_15_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_117 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_524 ),
	.datab(!Xd_0__inst_mult_14_529 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_370 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_379 ),
	.cout(Xd_0__inst_mult_14_380 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_118 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_534 ),
	.datab(!Xd_0__inst_mult_14_539 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_375 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_384 ),
	.cout(Xd_0__inst_mult_14_385 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_549 ),
	.datab(!Xd_0__inst_mult_9_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_404 ),
	.cout(Xd_0__inst_mult_9_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_559 ),
	.datab(!Xd_0__inst_mult_9_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_409 ),
	.cout(Xd_0__inst_mult_9_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_549 ),
	.datab(!Xd_0__inst_mult_8_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_404 ),
	.cout(Xd_0__inst_mult_8_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_559 ),
	.datab(!Xd_0__inst_mult_8_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_409 ),
	.cout(Xd_0__inst_mult_8_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_549 ),
	.datab(!Xd_0__inst_mult_11_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_404 ),
	.cout(Xd_0__inst_mult_11_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_559 ),
	.datab(!Xd_0__inst_mult_11_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_409 ),
	.cout(Xd_0__inst_mult_11_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_549 ),
	.datab(!Xd_0__inst_mult_10_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_404 ),
	.cout(Xd_0__inst_mult_10_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_559 ),
	.datab(!Xd_0__inst_mult_10_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_409 ),
	.cout(Xd_0__inst_mult_10_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_549 ),
	.datab(!Xd_0__inst_mult_5_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_404 ),
	.cout(Xd_0__inst_mult_5_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_559 ),
	.datab(!Xd_0__inst_mult_5_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_409 ),
	.cout(Xd_0__inst_mult_5_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_549 ),
	.datab(!Xd_0__inst_mult_4_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_404 ),
	.cout(Xd_0__inst_mult_4_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_559 ),
	.datab(!Xd_0__inst_mult_4_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_409 ),
	.cout(Xd_0__inst_mult_4_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_549 ),
	.datab(!Xd_0__inst_mult_7_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_404 ),
	.cout(Xd_0__inst_mult_7_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_559 ),
	.datab(!Xd_0__inst_mult_7_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_409 ),
	.cout(Xd_0__inst_mult_7_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_549 ),
	.datab(!Xd_0__inst_mult_6_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_404 ),
	.cout(Xd_0__inst_mult_6_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_559 ),
	.datab(!Xd_0__inst_mult_6_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_409 ),
	.cout(Xd_0__inst_mult_6_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_549 ),
	.datab(!Xd_0__inst_mult_1_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_404 ),
	.cout(Xd_0__inst_mult_1_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_559 ),
	.datab(!Xd_0__inst_mult_1_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_409 ),
	.cout(Xd_0__inst_mult_1_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_549 ),
	.datab(!Xd_0__inst_mult_0_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_404 ),
	.cout(Xd_0__inst_mult_0_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_559 ),
	.datab(!Xd_0__inst_mult_0_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_409 ),
	.cout(Xd_0__inst_mult_0_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_549 ),
	.datab(!Xd_0__inst_mult_3_554 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_404 ),
	.cout(Xd_0__inst_mult_3_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_559 ),
	.datab(!Xd_0__inst_mult_3_564 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_409 ),
	.cout(Xd_0__inst_mult_3_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_594 ),
	.datab(!Xd_0__inst_mult_2_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_449 ),
	.cout(Xd_0__inst_mult_2_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_604 ),
	.datab(!Xd_0__inst_mult_2_609 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_454 ),
	.cout(Xd_0__inst_mult_2_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_524 ),
	.datab(!Xd_0__inst_mult_29_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_454 ),
	.cout(Xd_0__inst_mult_29_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_599 ),
	.datab(!Xd_0__inst_mult_29_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_459 ),
	.cout(Xd_0__inst_mult_29_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_569 ),
	.datab(!Xd_0__inst_mult_28_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_414 ),
	.cout(Xd_0__inst_mult_28_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_579 ),
	.datab(!Xd_0__inst_mult_28_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_419 ),
	.cout(Xd_0__inst_mult_28_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_569 ),
	.datab(!Xd_0__inst_mult_31_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_414 ),
	.cout(Xd_0__inst_mult_31_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_579 ),
	.datab(!Xd_0__inst_mult_31_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_419 ),
	.cout(Xd_0__inst_mult_31_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_569 ),
	.datab(!Xd_0__inst_mult_30_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_414 ),
	.cout(Xd_0__inst_mult_30_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_579 ),
	.datab(!Xd_0__inst_mult_30_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_419 ),
	.cout(Xd_0__inst_mult_30_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_614 ),
	.datab(!Xd_0__inst_mult_25_619 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_504 ),
	.cout(Xd_0__inst_mult_25_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_24_180 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_24_724 ),
	.datab(!Xd_0__inst_mult_24_769 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_694 ),
	.cout(Xd_0__inst_mult_24_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_614 ),
	.datab(!Xd_0__inst_mult_27_619 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_504 ),
	.cout(Xd_0__inst_mult_27_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_26_180 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_26_709 ),
	.datab(!Xd_0__inst_mult_26_769 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_694 ),
	.cout(Xd_0__inst_mult_26_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_524 ),
	.datab(!Xd_0__inst_mult_21_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_454 ),
	.cout(Xd_0__inst_mult_21_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_599 ),
	.datab(!Xd_0__inst_mult_21_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_459 ),
	.cout(Xd_0__inst_mult_21_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_524 ),
	.datab(!Xd_0__inst_mult_20_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_454 ),
	.cout(Xd_0__inst_mult_20_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_599 ),
	.datab(!Xd_0__inst_mult_20_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_459 ),
	.cout(Xd_0__inst_mult_20_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_524 ),
	.datab(!Xd_0__inst_mult_23_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_454 ),
	.cout(Xd_0__inst_mult_23_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_599 ),
	.datab(!Xd_0__inst_mult_23_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_459 ),
	.cout(Xd_0__inst_mult_23_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_524 ),
	.datab(!Xd_0__inst_mult_22_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_454 ),
	.cout(Xd_0__inst_mult_22_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_599 ),
	.datab(!Xd_0__inst_mult_22_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_459 ),
	.cout(Xd_0__inst_mult_22_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_524 ),
	.datab(!Xd_0__inst_mult_17_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_454 ),
	.cout(Xd_0__inst_mult_17_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_599 ),
	.datab(!Xd_0__inst_mult_17_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_459 ),
	.cout(Xd_0__inst_mult_17_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_524 ),
	.datab(!Xd_0__inst_mult_16_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_454 ),
	.cout(Xd_0__inst_mult_16_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_599 ),
	.datab(!Xd_0__inst_mult_16_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_459 ),
	.cout(Xd_0__inst_mult_16_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_524 ),
	.datab(!Xd_0__inst_mult_19_519 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_454 ),
	.cout(Xd_0__inst_mult_19_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_599 ),
	.datab(!Xd_0__inst_mult_19_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_459 ),
	.cout(Xd_0__inst_mult_19_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_544 ),
	.datab(!Xd_0__inst_mult_18_549 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_389 ),
	.cout(Xd_0__inst_mult_18_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_554 ),
	.datab(!Xd_0__inst_mult_18_559 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_394 ),
	.cout(Xd_0__inst_mult_18_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_569 ),
	.datab(!Xd_0__inst_mult_13_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_414 ),
	.cout(Xd_0__inst_mult_13_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_579 ),
	.datab(!Xd_0__inst_mult_13_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_419 ),
	.cout(Xd_0__inst_mult_13_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_544 ),
	.datab(!Xd_0__inst_mult_12_549 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_389 ),
	.cout(Xd_0__inst_mult_12_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_554 ),
	.datab(!Xd_0__inst_mult_12_559 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_394 ),
	.cout(Xd_0__inst_mult_12_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_544 ),
	.datab(!Xd_0__inst_mult_15_549 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_389 ),
	.cout(Xd_0__inst_mult_15_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_554 ),
	.datab(!Xd_0__inst_mult_15_559 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_394 ),
	.cout(Xd_0__inst_mult_15_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_119 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_544 ),
	.datab(!Xd_0__inst_mult_14_549 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_380 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_389 ),
	.cout(Xd_0__inst_mult_14_390 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_120 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_554 ),
	.datab(!Xd_0__inst_mult_14_559 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_385 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_394 ),
	.cout(Xd_0__inst_mult_14_395 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_569 ),
	.datab(!Xd_0__inst_mult_9_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_414 ),
	.cout(Xd_0__inst_mult_9_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_579 ),
	.datab(!Xd_0__inst_mult_9_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_419 ),
	.cout(Xd_0__inst_mult_9_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_569 ),
	.datab(!Xd_0__inst_mult_8_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_414 ),
	.cout(Xd_0__inst_mult_8_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_579 ),
	.datab(!Xd_0__inst_mult_8_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_419 ),
	.cout(Xd_0__inst_mult_8_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_569 ),
	.datab(!Xd_0__inst_mult_11_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_414 ),
	.cout(Xd_0__inst_mult_11_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_579 ),
	.datab(!Xd_0__inst_mult_11_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_419 ),
	.cout(Xd_0__inst_mult_11_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_569 ),
	.datab(!Xd_0__inst_mult_10_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_414 ),
	.cout(Xd_0__inst_mult_10_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_579 ),
	.datab(!Xd_0__inst_mult_10_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_419 ),
	.cout(Xd_0__inst_mult_10_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_569 ),
	.datab(!Xd_0__inst_mult_5_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_414 ),
	.cout(Xd_0__inst_mult_5_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_579 ),
	.datab(!Xd_0__inst_mult_5_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_419 ),
	.cout(Xd_0__inst_mult_5_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_569 ),
	.datab(!Xd_0__inst_mult_4_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_414 ),
	.cout(Xd_0__inst_mult_4_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_579 ),
	.datab(!Xd_0__inst_mult_4_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_419 ),
	.cout(Xd_0__inst_mult_4_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_569 ),
	.datab(!Xd_0__inst_mult_7_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_414 ),
	.cout(Xd_0__inst_mult_7_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_579 ),
	.datab(!Xd_0__inst_mult_7_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_419 ),
	.cout(Xd_0__inst_mult_7_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_569 ),
	.datab(!Xd_0__inst_mult_6_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_414 ),
	.cout(Xd_0__inst_mult_6_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_579 ),
	.datab(!Xd_0__inst_mult_6_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_419 ),
	.cout(Xd_0__inst_mult_6_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_569 ),
	.datab(!Xd_0__inst_mult_1_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_414 ),
	.cout(Xd_0__inst_mult_1_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_579 ),
	.datab(!Xd_0__inst_mult_1_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_419 ),
	.cout(Xd_0__inst_mult_1_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_569 ),
	.datab(!Xd_0__inst_mult_0_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_414 ),
	.cout(Xd_0__inst_mult_0_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_579 ),
	.datab(!Xd_0__inst_mult_0_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_419 ),
	.cout(Xd_0__inst_mult_0_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_569 ),
	.datab(!Xd_0__inst_mult_3_574 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_414 ),
	.cout(Xd_0__inst_mult_3_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_579 ),
	.datab(!Xd_0__inst_mult_3_584 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_419 ),
	.cout(Xd_0__inst_mult_3_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_614 ),
	.datab(!Xd_0__inst_mult_2_619 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_459 ),
	.cout(Xd_0__inst_mult_2_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_624 ),
	.datab(!Xd_0__inst_mult_2_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_464 ),
	.cout(Xd_0__inst_mult_2_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_609 ),
	.datab(!Xd_0__inst_mult_29_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_464 ),
	.cout(Xd_0__inst_mult_29_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_589 ),
	.datab(!Xd_0__inst_mult_28_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_424 ),
	.cout(Xd_0__inst_mult_28_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_599 ),
	.datab(!Xd_0__inst_mult_28_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_429 ),
	.cout(Xd_0__inst_mult_28_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_589 ),
	.datab(!Xd_0__inst_mult_31_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_424 ),
	.cout(Xd_0__inst_mult_31_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_599 ),
	.datab(!Xd_0__inst_mult_31_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_429 ),
	.cout(Xd_0__inst_mult_31_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_589 ),
	.datab(!Xd_0__inst_mult_30_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_424 ),
	.cout(Xd_0__inst_mult_30_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_599 ),
	.datab(!Xd_0__inst_mult_30_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_429 ),
	.cout(Xd_0__inst_mult_30_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_624 ),
	.datab(!Xd_0__inst_mult_25_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_509 ),
	.cout(Xd_0__inst_mult_25_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_624 ),
	.datab(!Xd_0__inst_mult_27_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_509 ),
	.cout(Xd_0__inst_mult_27_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_609 ),
	.datab(!Xd_0__inst_mult_21_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_464 ),
	.cout(Xd_0__inst_mult_21_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_609 ),
	.datab(!Xd_0__inst_mult_20_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_464 ),
	.cout(Xd_0__inst_mult_20_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_609 ),
	.datab(!Xd_0__inst_mult_23_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_464 ),
	.cout(Xd_0__inst_mult_23_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_609 ),
	.datab(!Xd_0__inst_mult_22_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_464 ),
	.cout(Xd_0__inst_mult_22_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_609 ),
	.datab(!Xd_0__inst_mult_17_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_464 ),
	.cout(Xd_0__inst_mult_17_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_609 ),
	.datab(!Xd_0__inst_mult_16_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_464 ),
	.cout(Xd_0__inst_mult_16_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_609 ),
	.datab(!Xd_0__inst_mult_19_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_464 ),
	.cout(Xd_0__inst_mult_19_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_564 ),
	.datab(!Xd_0__inst_mult_18_569 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_399 ),
	.cout(Xd_0__inst_mult_18_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_574 ),
	.datab(!Xd_0__inst_mult_18_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_404 ),
	.cout(Xd_0__inst_mult_18_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_589 ),
	.datab(!Xd_0__inst_mult_13_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_424 ),
	.cout(Xd_0__inst_mult_13_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_599 ),
	.datab(!Xd_0__inst_mult_13_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_429 ),
	.cout(Xd_0__inst_mult_13_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_564 ),
	.datab(!Xd_0__inst_mult_12_569 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_399 ),
	.cout(Xd_0__inst_mult_12_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_574 ),
	.datab(!Xd_0__inst_mult_12_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_404 ),
	.cout(Xd_0__inst_mult_12_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_564 ),
	.datab(!Xd_0__inst_mult_15_569 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_399 ),
	.cout(Xd_0__inst_mult_15_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_574 ),
	.datab(!Xd_0__inst_mult_15_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_404 ),
	.cout(Xd_0__inst_mult_15_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_121 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_564 ),
	.datab(!Xd_0__inst_mult_14_569 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_399 ),
	.cout(Xd_0__inst_mult_14_400 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_122 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_574 ),
	.datab(!Xd_0__inst_mult_14_579 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_404 ),
	.cout(Xd_0__inst_mult_14_405 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_589 ),
	.datab(!Xd_0__inst_mult_9_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_424 ),
	.cout(Xd_0__inst_mult_9_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_599 ),
	.datab(!Xd_0__inst_mult_9_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_429 ),
	.cout(Xd_0__inst_mult_9_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_589 ),
	.datab(!Xd_0__inst_mult_8_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_424 ),
	.cout(Xd_0__inst_mult_8_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_599 ),
	.datab(!Xd_0__inst_mult_8_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_429 ),
	.cout(Xd_0__inst_mult_8_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_589 ),
	.datab(!Xd_0__inst_mult_11_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_424 ),
	.cout(Xd_0__inst_mult_11_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_599 ),
	.datab(!Xd_0__inst_mult_11_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_429 ),
	.cout(Xd_0__inst_mult_11_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_589 ),
	.datab(!Xd_0__inst_mult_10_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_424 ),
	.cout(Xd_0__inst_mult_10_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_599 ),
	.datab(!Xd_0__inst_mult_10_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_429 ),
	.cout(Xd_0__inst_mult_10_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_589 ),
	.datab(!Xd_0__inst_mult_5_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_424 ),
	.cout(Xd_0__inst_mult_5_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_599 ),
	.datab(!Xd_0__inst_mult_5_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_429 ),
	.cout(Xd_0__inst_mult_5_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_589 ),
	.datab(!Xd_0__inst_mult_4_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_424 ),
	.cout(Xd_0__inst_mult_4_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_599 ),
	.datab(!Xd_0__inst_mult_4_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_429 ),
	.cout(Xd_0__inst_mult_4_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_589 ),
	.datab(!Xd_0__inst_mult_7_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_424 ),
	.cout(Xd_0__inst_mult_7_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_599 ),
	.datab(!Xd_0__inst_mult_7_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_429 ),
	.cout(Xd_0__inst_mult_7_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_589 ),
	.datab(!Xd_0__inst_mult_6_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_424 ),
	.cout(Xd_0__inst_mult_6_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_599 ),
	.datab(!Xd_0__inst_mult_6_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_429 ),
	.cout(Xd_0__inst_mult_6_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_589 ),
	.datab(!Xd_0__inst_mult_1_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_424 ),
	.cout(Xd_0__inst_mult_1_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_599 ),
	.datab(!Xd_0__inst_mult_1_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_429 ),
	.cout(Xd_0__inst_mult_1_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_589 ),
	.datab(!Xd_0__inst_mult_0_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_424 ),
	.cout(Xd_0__inst_mult_0_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_599 ),
	.datab(!Xd_0__inst_mult_0_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_429 ),
	.cout(Xd_0__inst_mult_0_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_589 ),
	.datab(!Xd_0__inst_mult_3_594 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_424 ),
	.cout(Xd_0__inst_mult_3_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_599 ),
	.datab(!Xd_0__inst_mult_3_604 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_429 ),
	.cout(Xd_0__inst_mult_3_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_634 ),
	.datab(!Xd_0__inst_mult_2_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_469 ),
	.cout(Xd_0__inst_mult_2_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_644 ),
	.datab(!Xd_0__inst_mult_2_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_474 ),
	.cout(Xd_0__inst_mult_2_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_619 ),
	.datab(!Xd_0__inst_mult_29_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_469 ),
	.cout(Xd_0__inst_mult_29_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_494 ),
	.datab(!Xd_0__inst_mult_28_489 ),
	.datac(!din_a[346]),
	.datad(!din_b[338]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_434 ),
	.cout(Xd_0__inst_mult_28_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_609 ),
	.datab(!Xd_0__inst_mult_28_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_439 ),
	.cout(Xd_0__inst_mult_28_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_494 ),
	.datab(!Xd_0__inst_mult_31_489 ),
	.datac(!din_a[382]),
	.datad(!din_b[374]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_434 ),
	.cout(Xd_0__inst_mult_31_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_609 ),
	.datab(!Xd_0__inst_mult_31_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_439 ),
	.cout(Xd_0__inst_mult_31_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_494 ),
	.datab(!Xd_0__inst_mult_30_489 ),
	.datac(!din_a[370]),
	.datad(!din_b[362]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_434 ),
	.cout(Xd_0__inst_mult_30_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_609 ),
	.datab(!Xd_0__inst_mult_30_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_439 ),
	.cout(Xd_0__inst_mult_30_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_144 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_634 ),
	.datab(!Xd_0__inst_mult_25_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_514 ),
	.cout(Xd_0__inst_mult_25_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_144 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_634 ),
	.datab(!Xd_0__inst_mult_27_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_514 ),
	.cout(Xd_0__inst_mult_27_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_619 ),
	.datab(!Xd_0__inst_mult_21_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_469 ),
	.cout(Xd_0__inst_mult_21_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_619 ),
	.datab(!Xd_0__inst_mult_20_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_469 ),
	.cout(Xd_0__inst_mult_20_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_619 ),
	.datab(!Xd_0__inst_mult_23_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_469 ),
	.cout(Xd_0__inst_mult_23_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_619 ),
	.datab(!Xd_0__inst_mult_22_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_469 ),
	.cout(Xd_0__inst_mult_22_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_619 ),
	.datab(!Xd_0__inst_mult_17_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_469 ),
	.cout(Xd_0__inst_mult_17_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_619 ),
	.datab(!Xd_0__inst_mult_16_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_469 ),
	.cout(Xd_0__inst_mult_16_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_619 ),
	.datab(!Xd_0__inst_mult_19_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_469 ),
	.cout(Xd_0__inst_mult_19_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_584 ),
	.datab(!Xd_0__inst_mult_18_589 ),
	.datac(!din_a[226]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_409 ),
	.cout(Xd_0__inst_mult_18_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_594 ),
	.datab(!Xd_0__inst_mult_18_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_414 ),
	.cout(Xd_0__inst_mult_18_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_494 ),
	.datab(!Xd_0__inst_mult_13_489 ),
	.datac(!din_a[166]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_434 ),
	.cout(Xd_0__inst_mult_13_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_609 ),
	.datab(!Xd_0__inst_mult_13_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_439 ),
	.cout(Xd_0__inst_mult_13_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_584 ),
	.datab(!Xd_0__inst_mult_12_589 ),
	.datac(!din_a[154]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_409 ),
	.cout(Xd_0__inst_mult_12_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_594 ),
	.datab(!Xd_0__inst_mult_12_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_414 ),
	.cout(Xd_0__inst_mult_12_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_584 ),
	.datab(!Xd_0__inst_mult_15_589 ),
	.datac(!din_a[190]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_409 ),
	.cout(Xd_0__inst_mult_15_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_594 ),
	.datab(!Xd_0__inst_mult_15_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_414 ),
	.cout(Xd_0__inst_mult_15_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_123 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_584 ),
	.datab(!Xd_0__inst_mult_14_589 ),
	.datac(!din_a[178]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_409 ),
	.cout(Xd_0__inst_mult_14_410 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_124 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_594 ),
	.datab(!Xd_0__inst_mult_14_599 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_405 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_414 ),
	.cout(Xd_0__inst_mult_14_415 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_494 ),
	.datab(!Xd_0__inst_mult_9_489 ),
	.datac(!din_a[118]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_434 ),
	.cout(Xd_0__inst_mult_9_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_609 ),
	.datab(!Xd_0__inst_mult_9_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_439 ),
	.cout(Xd_0__inst_mult_9_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_494 ),
	.datab(!Xd_0__inst_mult_8_489 ),
	.datac(!din_a[106]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_434 ),
	.cout(Xd_0__inst_mult_8_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_609 ),
	.datab(!Xd_0__inst_mult_8_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_439 ),
	.cout(Xd_0__inst_mult_8_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_494 ),
	.datab(!Xd_0__inst_mult_11_489 ),
	.datac(!din_a[142]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_434 ),
	.cout(Xd_0__inst_mult_11_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_609 ),
	.datab(!Xd_0__inst_mult_11_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_439 ),
	.cout(Xd_0__inst_mult_11_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_494 ),
	.datab(!Xd_0__inst_mult_10_489 ),
	.datac(!din_a[130]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_434 ),
	.cout(Xd_0__inst_mult_10_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_609 ),
	.datab(!Xd_0__inst_mult_10_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_439 ),
	.cout(Xd_0__inst_mult_10_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_494 ),
	.datab(!Xd_0__inst_mult_5_489 ),
	.datac(!din_a[70]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_434 ),
	.cout(Xd_0__inst_mult_5_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_609 ),
	.datab(!Xd_0__inst_mult_5_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_439 ),
	.cout(Xd_0__inst_mult_5_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_494 ),
	.datab(!Xd_0__inst_mult_4_489 ),
	.datac(!din_a[58]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_434 ),
	.cout(Xd_0__inst_mult_4_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_609 ),
	.datab(!Xd_0__inst_mult_4_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_439 ),
	.cout(Xd_0__inst_mult_4_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_494 ),
	.datab(!Xd_0__inst_mult_7_489 ),
	.datac(!din_a[94]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_434 ),
	.cout(Xd_0__inst_mult_7_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_609 ),
	.datab(!Xd_0__inst_mult_7_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_439 ),
	.cout(Xd_0__inst_mult_7_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_494 ),
	.datab(!Xd_0__inst_mult_6_489 ),
	.datac(!din_a[82]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_434 ),
	.cout(Xd_0__inst_mult_6_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_609 ),
	.datab(!Xd_0__inst_mult_6_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_439 ),
	.cout(Xd_0__inst_mult_6_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_494 ),
	.datab(!Xd_0__inst_mult_1_489 ),
	.datac(!din_a[22]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_434 ),
	.cout(Xd_0__inst_mult_1_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_609 ),
	.datab(!Xd_0__inst_mult_1_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_439 ),
	.cout(Xd_0__inst_mult_1_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_494 ),
	.datab(!Xd_0__inst_mult_0_489 ),
	.datac(!din_a[10]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_434 ),
	.cout(Xd_0__inst_mult_0_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_609 ),
	.datab(!Xd_0__inst_mult_0_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_439 ),
	.cout(Xd_0__inst_mult_0_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_494 ),
	.datab(!Xd_0__inst_mult_3_489 ),
	.datac(!din_a[46]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_434 ),
	.cout(Xd_0__inst_mult_3_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_609 ),
	.datab(!Xd_0__inst_mult_3_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_439 ),
	.cout(Xd_0__inst_mult_3_440 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_539 ),
	.datab(!Xd_0__inst_mult_2_534 ),
	.datac(!din_a[34]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_479 ),
	.cout(Xd_0__inst_mult_2_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_654 ),
	.datab(!Xd_0__inst_mult_2_659 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_484 ),
	.cout(Xd_0__inst_mult_2_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_629 ),
	.datab(!Xd_0__inst_mult_29_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_474 ),
	.cout(Xd_0__inst_mult_29_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_619 ),
	.datab(!Xd_0__inst_mult_28_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_444 ),
	.cout(Xd_0__inst_mult_28_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_619 ),
	.datab(!Xd_0__inst_mult_31_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_444 ),
	.cout(Xd_0__inst_mult_31_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_619 ),
	.datab(!Xd_0__inst_mult_30_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_444 ),
	.cout(Xd_0__inst_mult_30_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_145 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_644 ),
	.datab(!Xd_0__inst_mult_25_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_519 ),
	.cout(Xd_0__inst_mult_25_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_145 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_644 ),
	.datab(!Xd_0__inst_mult_27_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_519 ),
	.cout(Xd_0__inst_mult_27_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_629 ),
	.datab(!Xd_0__inst_mult_21_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_474 ),
	.cout(Xd_0__inst_mult_21_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_629 ),
	.datab(!Xd_0__inst_mult_20_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_474 ),
	.cout(Xd_0__inst_mult_20_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_629 ),
	.datab(!Xd_0__inst_mult_23_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_474 ),
	.cout(Xd_0__inst_mult_23_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_629 ),
	.datab(!Xd_0__inst_mult_22_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_474 ),
	.cout(Xd_0__inst_mult_22_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_629 ),
	.datab(!Xd_0__inst_mult_17_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_474 ),
	.cout(Xd_0__inst_mult_17_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_629 ),
	.datab(!Xd_0__inst_mult_16_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_474 ),
	.cout(Xd_0__inst_mult_16_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_629 ),
	.datab(!Xd_0__inst_mult_19_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_474 ),
	.cout(Xd_0__inst_mult_19_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_604 ),
	.datab(!Xd_0__inst_mult_18_55_sumout ),
	.datac(!Xd_0__inst_mult_18_584 ),
	.datad(!Xd_0__inst_mult_18_589 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_419 ),
	.cout(Xd_0__inst_mult_18_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_609 ),
	.datab(!Xd_0__inst_mult_18_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_424 ),
	.cout(Xd_0__inst_mult_18_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_619 ),
	.datab(!Xd_0__inst_mult_13_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_444 ),
	.cout(Xd_0__inst_mult_13_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_604 ),
	.datab(!Xd_0__inst_mult_12_40_sumout ),
	.datac(!Xd_0__inst_mult_12_584 ),
	.datad(!Xd_0__inst_mult_12_589 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_419 ),
	.cout(Xd_0__inst_mult_12_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_609 ),
	.datab(!Xd_0__inst_mult_12_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_424 ),
	.cout(Xd_0__inst_mult_12_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_604 ),
	.datab(!Xd_0__inst_mult_15_65_sumout ),
	.datac(!Xd_0__inst_mult_15_584 ),
	.datad(!Xd_0__inst_mult_15_589 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_419 ),
	.cout(Xd_0__inst_mult_15_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_609 ),
	.datab(!Xd_0__inst_mult_15_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_424 ),
	.cout(Xd_0__inst_mult_15_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_125 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_604 ),
	.datab(!Xd_0__inst_mult_14_45_sumout ),
	.datac(!Xd_0__inst_mult_14_584 ),
	.datad(!Xd_0__inst_mult_14_589 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_410 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_419 ),
	.cout(Xd_0__inst_mult_14_420 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_126 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_609 ),
	.datab(!Xd_0__inst_mult_14_614 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_424 ),
	.cout(Xd_0__inst_mult_14_425 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_619 ),
	.datab(!Xd_0__inst_mult_9_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_444 ),
	.cout(Xd_0__inst_mult_9_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_619 ),
	.datab(!Xd_0__inst_mult_8_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_444 ),
	.cout(Xd_0__inst_mult_8_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_619 ),
	.datab(!Xd_0__inst_mult_11_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_444 ),
	.cout(Xd_0__inst_mult_11_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_619 ),
	.datab(!Xd_0__inst_mult_10_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_444 ),
	.cout(Xd_0__inst_mult_10_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_619 ),
	.datab(!Xd_0__inst_mult_5_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_444 ),
	.cout(Xd_0__inst_mult_5_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_619 ),
	.datab(!Xd_0__inst_mult_4_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_444 ),
	.cout(Xd_0__inst_mult_4_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_619 ),
	.datab(!Xd_0__inst_mult_7_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_444 ),
	.cout(Xd_0__inst_mult_7_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_619 ),
	.datab(!Xd_0__inst_mult_6_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_444 ),
	.cout(Xd_0__inst_mult_6_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_619 ),
	.datab(!Xd_0__inst_mult_1_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_444 ),
	.cout(Xd_0__inst_mult_1_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_619 ),
	.datab(!Xd_0__inst_mult_0_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_444 ),
	.cout(Xd_0__inst_mult_0_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_619 ),
	.datab(!Xd_0__inst_mult_3_624 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_440 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_444 ),
	.cout(Xd_0__inst_mult_3_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_664 ),
	.datab(!Xd_0__inst_mult_2_669 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_489 ),
	.cout(Xd_0__inst_mult_2_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_639 ),
	.datab(!Xd_0__inst_mult_29_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_479 ),
	.cout(Xd_0__inst_mult_29_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_629 ),
	.datab(!Xd_0__inst_mult_28_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_449 ),
	.cout(Xd_0__inst_mult_28_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_629 ),
	.datab(!Xd_0__inst_mult_31_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_449 ),
	.cout(Xd_0__inst_mult_31_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_629 ),
	.datab(!Xd_0__inst_mult_30_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_449 ),
	.cout(Xd_0__inst_mult_30_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_146 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_654 ),
	.datab(!Xd_0__inst_mult_25_659 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_524 ),
	.cout(Xd_0__inst_mult_25_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_146 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_654 ),
	.datab(!Xd_0__inst_mult_27_659 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_524 ),
	.cout(Xd_0__inst_mult_27_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_639 ),
	.datab(!Xd_0__inst_mult_21_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_479 ),
	.cout(Xd_0__inst_mult_21_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_639 ),
	.datab(!Xd_0__inst_mult_20_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_479 ),
	.cout(Xd_0__inst_mult_20_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_639 ),
	.datab(!Xd_0__inst_mult_23_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_479 ),
	.cout(Xd_0__inst_mult_23_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_639 ),
	.datab(!Xd_0__inst_mult_22_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_479 ),
	.cout(Xd_0__inst_mult_22_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_639 ),
	.datab(!Xd_0__inst_mult_17_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_479 ),
	.cout(Xd_0__inst_mult_17_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_639 ),
	.datab(!Xd_0__inst_mult_16_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_479 ),
	.cout(Xd_0__inst_mult_16_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_639 ),
	.datab(!Xd_0__inst_mult_19_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_479 ),
	.cout(Xd_0__inst_mult_19_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_619 ),
	.datab(!Xd_0__inst_mult_18_50_sumout ),
	.datac(!Xd_0__inst_mult_18_604 ),
	.datad(!Xd_0__inst_mult_18_55_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_429 ),
	.cout(Xd_0__inst_mult_18_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_624 ),
	.datab(!Xd_0__inst_mult_18_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_434 ),
	.cout(Xd_0__inst_mult_18_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_629 ),
	.datab(!Xd_0__inst_mult_13_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_449 ),
	.cout(Xd_0__inst_mult_13_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_619 ),
	.datab(!Xd_0__inst_mult_12_70_sumout ),
	.datac(!Xd_0__inst_mult_12_604 ),
	.datad(!Xd_0__inst_mult_12_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_429 ),
	.cout(Xd_0__inst_mult_12_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_624 ),
	.datab(!Xd_0__inst_mult_12_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_434 ),
	.cout(Xd_0__inst_mult_12_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_619 ),
	.datab(!Xd_0__inst_mult_15_55_sumout ),
	.datac(!Xd_0__inst_mult_15_604 ),
	.datad(!Xd_0__inst_mult_15_65_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_429 ),
	.cout(Xd_0__inst_mult_15_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_624 ),
	.datab(!Xd_0__inst_mult_15_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_434 ),
	.cout(Xd_0__inst_mult_15_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_127 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_619 ),
	.datab(!Xd_0__inst_mult_14_75_sumout ),
	.datac(!Xd_0__inst_mult_14_604 ),
	.datad(!Xd_0__inst_mult_14_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_429 ),
	.cout(Xd_0__inst_mult_14_430 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_128 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_624 ),
	.datab(!Xd_0__inst_mult_14_629 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_425 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_434 ),
	.cout(Xd_0__inst_mult_14_435 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_629 ),
	.datab(!Xd_0__inst_mult_9_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_449 ),
	.cout(Xd_0__inst_mult_9_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_629 ),
	.datab(!Xd_0__inst_mult_8_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_449 ),
	.cout(Xd_0__inst_mult_8_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_629 ),
	.datab(!Xd_0__inst_mult_11_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_449 ),
	.cout(Xd_0__inst_mult_11_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_629 ),
	.datab(!Xd_0__inst_mult_10_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_449 ),
	.cout(Xd_0__inst_mult_10_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_629 ),
	.datab(!Xd_0__inst_mult_5_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_449 ),
	.cout(Xd_0__inst_mult_5_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_629 ),
	.datab(!Xd_0__inst_mult_4_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_449 ),
	.cout(Xd_0__inst_mult_4_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_629 ),
	.datab(!Xd_0__inst_mult_7_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_449 ),
	.cout(Xd_0__inst_mult_7_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_629 ),
	.datab(!Xd_0__inst_mult_6_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_449 ),
	.cout(Xd_0__inst_mult_6_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_629 ),
	.datab(!Xd_0__inst_mult_1_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_449 ),
	.cout(Xd_0__inst_mult_1_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_629 ),
	.datab(!Xd_0__inst_mult_0_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_449 ),
	.cout(Xd_0__inst_mult_0_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_629 ),
	.datab(!Xd_0__inst_mult_3_634 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_449 ),
	.cout(Xd_0__inst_mult_3_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_674 ),
	.datab(!Xd_0__inst_mult_2_679 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_494 ),
	.cout(Xd_0__inst_mult_2_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_649 ),
	.datab(!Xd_0__inst_mult_29_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_484 ),
	.cout(Xd_0__inst_mult_29_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_639 ),
	.datab(!Xd_0__inst_mult_28_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_454 ),
	.cout(Xd_0__inst_mult_28_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_639 ),
	.datab(!Xd_0__inst_mult_31_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_454 ),
	.cout(Xd_0__inst_mult_31_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_639 ),
	.datab(!Xd_0__inst_mult_30_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_454 ),
	.cout(Xd_0__inst_mult_30_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_147 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_664 ),
	.datab(!Xd_0__inst_mult_25_669 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_529 ),
	.cout(Xd_0__inst_mult_25_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_147 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_664 ),
	.datab(!Xd_0__inst_mult_27_669 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_529 ),
	.cout(Xd_0__inst_mult_27_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_649 ),
	.datab(!Xd_0__inst_mult_21_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_484 ),
	.cout(Xd_0__inst_mult_21_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_649 ),
	.datab(!Xd_0__inst_mult_20_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_484 ),
	.cout(Xd_0__inst_mult_20_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_649 ),
	.datab(!Xd_0__inst_mult_23_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_484 ),
	.cout(Xd_0__inst_mult_23_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_649 ),
	.datab(!Xd_0__inst_mult_22_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_484 ),
	.cout(Xd_0__inst_mult_22_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_649 ),
	.datab(!Xd_0__inst_mult_17_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_484 ),
	.cout(Xd_0__inst_mult_17_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_649 ),
	.datab(!Xd_0__inst_mult_16_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_484 ),
	.cout(Xd_0__inst_mult_16_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_138 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_649 ),
	.datab(!Xd_0__inst_mult_19_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_484 ),
	.cout(Xd_0__inst_mult_19_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_619 ),
	.datab(!Xd_0__inst_mult_18_50_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_439 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_634 ),
	.datab(!Xd_0__inst_mult_18_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_444 ),
	.cout(Xd_0__inst_mult_18_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_639 ),
	.datab(!Xd_0__inst_mult_13_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_454 ),
	.cout(Xd_0__inst_mult_13_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_619 ),
	.datab(!Xd_0__inst_mult_12_70_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_439 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_634 ),
	.datab(!Xd_0__inst_mult_12_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_444 ),
	.cout(Xd_0__inst_mult_12_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_619 ),
	.datab(!Xd_0__inst_mult_15_55_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_439 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_634 ),
	.datab(!Xd_0__inst_mult_15_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_444 ),
	.cout(Xd_0__inst_mult_15_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_129 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_619 ),
	.datab(!Xd_0__inst_mult_14_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_439 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_130 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_634 ),
	.datab(!Xd_0__inst_mult_14_639 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_435 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_444 ),
	.cout(Xd_0__inst_mult_14_445 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_639 ),
	.datab(!Xd_0__inst_mult_9_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_454 ),
	.cout(Xd_0__inst_mult_9_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_639 ),
	.datab(!Xd_0__inst_mult_8_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_454 ),
	.cout(Xd_0__inst_mult_8_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_639 ),
	.datab(!Xd_0__inst_mult_11_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_454 ),
	.cout(Xd_0__inst_mult_11_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_639 ),
	.datab(!Xd_0__inst_mult_10_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_454 ),
	.cout(Xd_0__inst_mult_10_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_639 ),
	.datab(!Xd_0__inst_mult_5_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_454 ),
	.cout(Xd_0__inst_mult_5_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_639 ),
	.datab(!Xd_0__inst_mult_4_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_454 ),
	.cout(Xd_0__inst_mult_4_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_639 ),
	.datab(!Xd_0__inst_mult_7_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_454 ),
	.cout(Xd_0__inst_mult_7_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_639 ),
	.datab(!Xd_0__inst_mult_6_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_454 ),
	.cout(Xd_0__inst_mult_6_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_639 ),
	.datab(!Xd_0__inst_mult_1_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_454 ),
	.cout(Xd_0__inst_mult_1_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_639 ),
	.datab(!Xd_0__inst_mult_0_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_454 ),
	.cout(Xd_0__inst_mult_0_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_639 ),
	.datab(!Xd_0__inst_mult_3_644 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_454 ),
	.cout(Xd_0__inst_mult_3_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_684 ),
	.datab(!Xd_0__inst_mult_2_689 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_499 ),
	.cout(Xd_0__inst_mult_2_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_29_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_659 ),
	.datab(!Xd_0__inst_mult_29_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_489 ),
	.cout(Xd_0__inst_mult_29_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_60 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[354]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_60_sumout ),
	.cout(Xd_0__inst_mult_29_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_28_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_649 ),
	.datab(!Xd_0__inst_mult_28_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_459 ),
	.cout(Xd_0__inst_mult_28_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_31_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_649 ),
	.datab(!Xd_0__inst_mult_31_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_459 ),
	.cout(Xd_0__inst_mult_31_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_30_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_649 ),
	.datab(!Xd_0__inst_mult_30_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_459 ),
	.cout(Xd_0__inst_mult_30_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_60 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[366]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_60_sumout ),
	.cout(Xd_0__inst_mult_30_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_25_148 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_674 ),
	.datab(!Xd_0__inst_mult_25_679 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_534 ),
	.cout(Xd_0__inst_mult_25_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_65 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[306]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_65_sumout ),
	.cout(Xd_0__inst_mult_25_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_60 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[294]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_60_sumout ),
	.cout(Xd_0__inst_mult_24_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_27_148 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_674 ),
	.datab(!Xd_0__inst_mult_27_679 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_534 ),
	.cout(Xd_0__inst_mult_27_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_65 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[330]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_65_sumout ),
	.cout(Xd_0__inst_mult_27_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_60 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[318]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_60_sumout ),
	.cout(Xd_0__inst_mult_26_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_21_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_659 ),
	.datab(!Xd_0__inst_mult_21_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_489 ),
	.cout(Xd_0__inst_mult_21_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_55 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[258]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_55_sumout ),
	.cout(Xd_0__inst_mult_21_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_20_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_659 ),
	.datab(!Xd_0__inst_mult_20_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_489 ),
	.cout(Xd_0__inst_mult_20_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_65 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[246]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_65_sumout ),
	.cout(Xd_0__inst_mult_20_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_23_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_659 ),
	.datab(!Xd_0__inst_mult_23_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_489 ),
	.cout(Xd_0__inst_mult_23_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_50 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[282]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_50_sumout ),
	.cout(Xd_0__inst_mult_23_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_22_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_659 ),
	.datab(!Xd_0__inst_mult_22_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_489 ),
	.cout(Xd_0__inst_mult_22_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_55 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[270]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_55_sumout ),
	.cout(Xd_0__inst_mult_22_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_17_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_659 ),
	.datab(!Xd_0__inst_mult_17_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_489 ),
	.cout(Xd_0__inst_mult_17_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_16_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_659 ),
	.datab(!Xd_0__inst_mult_16_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_489 ),
	.cout(Xd_0__inst_mult_16_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_19_139 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_659 ),
	.datab(!Xd_0__inst_mult_19_664 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_489 ),
	.cout(Xd_0__inst_mult_19_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_55 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[234]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_55_sumout ),
	.cout(Xd_0__inst_mult_19_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_18_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_644 ),
	.datab(!Xd_0__inst_mult_18_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_449 ),
	.cout(Xd_0__inst_mult_18_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_60 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[222]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_60_sumout ),
	.cout(Xd_0__inst_mult_18_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_13_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_649 ),
	.datab(!Xd_0__inst_mult_13_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_459 ),
	.cout(Xd_0__inst_mult_13_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_55 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[162]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_55_sumout ),
	.cout(Xd_0__inst_mult_13_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_12_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_644 ),
	.datab(!Xd_0__inst_mult_12_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_449 ),
	.cout(Xd_0__inst_mult_12_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_50 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[150]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_50_sumout ),
	.cout(Xd_0__inst_mult_12_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_15_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_644 ),
	.datab(!Xd_0__inst_mult_15_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_449 ),
	.cout(Xd_0__inst_mult_15_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_70 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[186]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_70_sumout ),
	.cout(Xd_0__inst_mult_15_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_14_131 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_644 ),
	.datab(!Xd_0__inst_mult_14_649 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_445 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_449 ),
	.cout(Xd_0__inst_mult_14_450 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_50 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[174]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_50_sumout ),
	.cout(Xd_0__inst_mult_14_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_9_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_649 ),
	.datab(!Xd_0__inst_mult_9_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_459 ),
	.cout(Xd_0__inst_mult_9_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_60 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[114]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_60_sumout ),
	.cout(Xd_0__inst_mult_9_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_8_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_649 ),
	.datab(!Xd_0__inst_mult_8_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_459 ),
	.cout(Xd_0__inst_mult_8_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_70 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_70_sumout ),
	.cout(Xd_0__inst_mult_8_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_11_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_649 ),
	.datab(!Xd_0__inst_mult_11_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_459 ),
	.cout(Xd_0__inst_mult_11_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_50 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[138]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_50_sumout ),
	.cout(Xd_0__inst_mult_11_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_10_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_649 ),
	.datab(!Xd_0__inst_mult_10_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_459 ),
	.cout(Xd_0__inst_mult_10_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_65 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[126]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_65_sumout ),
	.cout(Xd_0__inst_mult_10_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_5_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_649 ),
	.datab(!Xd_0__inst_mult_5_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_459 ),
	.cout(Xd_0__inst_mult_5_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_4_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_649 ),
	.datab(!Xd_0__inst_mult_4_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_459 ),
	.cout(Xd_0__inst_mult_4_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_50 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_50_sumout ),
	.cout(Xd_0__inst_mult_4_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_7_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_649 ),
	.datab(!Xd_0__inst_mult_7_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_459 ),
	.cout(Xd_0__inst_mult_7_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_65 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_65_sumout ),
	.cout(Xd_0__inst_mult_7_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_6_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_649 ),
	.datab(!Xd_0__inst_mult_6_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_459 ),
	.cout(Xd_0__inst_mult_6_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_65 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_65_sumout ),
	.cout(Xd_0__inst_mult_6_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_1_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_649 ),
	.datab(!Xd_0__inst_mult_1_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_459 ),
	.cout(Xd_0__inst_mult_1_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_50 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_50_sumout ),
	.cout(Xd_0__inst_mult_1_51 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_0_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_649 ),
	.datab(!Xd_0__inst_mult_0_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_459 ),
	.cout(Xd_0__inst_mult_0_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_60 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_51 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_60_sumout ),
	.cout(Xd_0__inst_mult_0_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_3_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_649 ),
	.datab(!Xd_0__inst_mult_3_654 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_459 ),
	.cout(Xd_0__inst_mult_3_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_70 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_70_sumout ),
	.cout(Xd_0__inst_mult_3_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000011116666),
	.shared_arith("off")
) Xd_0__inst_mult_2_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_694 ),
	.datab(!Xd_0__inst_mult_2_699 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_504 ),
	.cout(Xd_0__inst_mult_2_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_60 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_60_sumout ),
	.cout(Xd_0__inst_mult_2_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_669 ),
	.datab(!Xd_0__inst_mult_29_674 ),
	.datac(!din_a[357]),
	.datad(!din_b[356]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_494 ),
	.cout(Xd_0__inst_mult_29_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_65 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[355]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_65_sumout ),
	.cout(Xd_0__inst_mult_29_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_659 ),
	.datab(!Xd_0__inst_mult_28_664 ),
	.datac(!din_a[345]),
	.datad(!din_b[344]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_464 ),
	.cout(Xd_0__inst_mult_28_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_65 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[343]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_65_sumout ),
	.cout(Xd_0__inst_mult_28_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_659 ),
	.datab(!Xd_0__inst_mult_31_664 ),
	.datac(!din_a[381]),
	.datad(!din_b[380]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_464 ),
	.cout(Xd_0__inst_mult_31_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_55 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[379]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_55_sumout ),
	.cout(Xd_0__inst_mult_31_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_659 ),
	.datab(!Xd_0__inst_mult_30_664 ),
	.datac(!din_a[369]),
	.datad(!din_b[368]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_464 ),
	.cout(Xd_0__inst_mult_30_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_65 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[367]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_65_sumout ),
	.cout(Xd_0__inst_mult_30_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_149 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_684 ),
	.datab(!Xd_0__inst_mult_25_689 ),
	.datac(!din_a[309]),
	.datad(!din_b[308]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_539 ),
	.cout(Xd_0__inst_mult_25_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_70 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[307]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_70_sumout ),
	.cout(Xd_0__inst_mult_25_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_65 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[295]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_65_sumout ),
	.cout(Xd_0__inst_mult_24_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_149 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_684 ),
	.datab(!Xd_0__inst_mult_27_689 ),
	.datac(!din_a[333]),
	.datad(!din_b[332]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_539 ),
	.cout(Xd_0__inst_mult_27_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_70 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[331]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_70_sumout ),
	.cout(Xd_0__inst_mult_27_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_65 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[319]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_65_sumout ),
	.cout(Xd_0__inst_mult_26_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_669 ),
	.datab(!Xd_0__inst_mult_21_674 ),
	.datac(!din_a[261]),
	.datad(!din_b[260]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_494 ),
	.cout(Xd_0__inst_mult_21_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_60 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[259]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_60_sumout ),
	.cout(Xd_0__inst_mult_21_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_669 ),
	.datab(!Xd_0__inst_mult_20_674 ),
	.datac(!din_a[249]),
	.datad(!din_b[248]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_494 ),
	.cout(Xd_0__inst_mult_20_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_70 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[247]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_70_sumout ),
	.cout(Xd_0__inst_mult_20_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_669 ),
	.datab(!Xd_0__inst_mult_23_674 ),
	.datac(!din_a[285]),
	.datad(!din_b[284]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_494 ),
	.cout(Xd_0__inst_mult_23_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_55 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[283]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_55_sumout ),
	.cout(Xd_0__inst_mult_23_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_669 ),
	.datab(!Xd_0__inst_mult_22_674 ),
	.datac(!din_a[273]),
	.datad(!din_b[272]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_494 ),
	.cout(Xd_0__inst_mult_22_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_60 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[271]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_60_sumout ),
	.cout(Xd_0__inst_mult_22_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_669 ),
	.datab(!Xd_0__inst_mult_17_674 ),
	.datac(!din_a[213]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_494 ),
	.cout(Xd_0__inst_mult_17_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_65 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[211]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_65_sumout ),
	.cout(Xd_0__inst_mult_17_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_669 ),
	.datab(!Xd_0__inst_mult_16_674 ),
	.datac(!din_a[201]),
	.datad(!din_b[200]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_494 ),
	.cout(Xd_0__inst_mult_16_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_55 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[199]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_55_sumout ),
	.cout(Xd_0__inst_mult_16_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_140 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_669 ),
	.datab(!Xd_0__inst_mult_19_674 ),
	.datac(!din_a[237]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_494 ),
	.cout(Xd_0__inst_mult_19_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_60 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[235]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_60_sumout ),
	.cout(Xd_0__inst_mult_19_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_654 ),
	.datab(!Xd_0__inst_mult_18_659 ),
	.datac(!din_a[225]),
	.datad(!din_b[224]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_454 ),
	.cout(Xd_0__inst_mult_18_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_65 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[223]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_65_sumout ),
	.cout(Xd_0__inst_mult_18_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_659 ),
	.datab(!Xd_0__inst_mult_13_664 ),
	.datac(!din_a[165]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_464 ),
	.cout(Xd_0__inst_mult_13_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_60 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_60_sumout ),
	.cout(Xd_0__inst_mult_13_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_654 ),
	.datab(!Xd_0__inst_mult_12_659 ),
	.datac(!din_a[153]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_454 ),
	.cout(Xd_0__inst_mult_12_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_55 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_55_sumout ),
	.cout(Xd_0__inst_mult_12_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_654 ),
	.datab(!Xd_0__inst_mult_15_659 ),
	.datac(!din_a[189]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_454 ),
	.cout(Xd_0__inst_mult_15_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_75 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_75_sumout ),
	.cout(Xd_0__inst_mult_15_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_132 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_654 ),
	.datab(!Xd_0__inst_mult_14_659 ),
	.datac(!din_a[177]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_450 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_454 ),
	.cout(Xd_0__inst_mult_14_455 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_55 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_55_sumout ),
	.cout(Xd_0__inst_mult_14_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_659 ),
	.datab(!Xd_0__inst_mult_9_664 ),
	.datac(!din_a[117]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_464 ),
	.cout(Xd_0__inst_mult_9_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_65 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[115]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_65_sumout ),
	.cout(Xd_0__inst_mult_9_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_659 ),
	.datab(!Xd_0__inst_mult_8_664 ),
	.datac(!din_a[105]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_464 ),
	.cout(Xd_0__inst_mult_8_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_75 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_75_sumout ),
	.cout(Xd_0__inst_mult_8_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_659 ),
	.datab(!Xd_0__inst_mult_11_664 ),
	.datac(!din_a[141]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_464 ),
	.cout(Xd_0__inst_mult_11_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_55 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_55_sumout ),
	.cout(Xd_0__inst_mult_11_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_659 ),
	.datab(!Xd_0__inst_mult_10_664 ),
	.datac(!din_a[129]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_464 ),
	.cout(Xd_0__inst_mult_10_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_70 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_70_sumout ),
	.cout(Xd_0__inst_mult_10_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_659 ),
	.datab(!Xd_0__inst_mult_5_664 ),
	.datac(!din_a[69]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_464 ),
	.cout(Xd_0__inst_mult_5_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_659 ),
	.datab(!Xd_0__inst_mult_4_664 ),
	.datac(!din_a[57]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_464 ),
	.cout(Xd_0__inst_mult_4_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_55 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_55_sumout ),
	.cout(Xd_0__inst_mult_4_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_659 ),
	.datab(!Xd_0__inst_mult_7_664 ),
	.datac(!din_a[93]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_464 ),
	.cout(Xd_0__inst_mult_7_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_70 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_i29_157 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_70_sumout ),
	.cout(Xd_0__inst_mult_7_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_659 ),
	.datab(!Xd_0__inst_mult_6_664 ),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_464 ),
	.cout(Xd_0__inst_mult_6_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_70 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_70_sumout ),
	.cout(Xd_0__inst_mult_6_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_659 ),
	.datab(!Xd_0__inst_mult_1_664 ),
	.datac(!din_a[21]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_464 ),
	.cout(Xd_0__inst_mult_1_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_55 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_55_sumout ),
	.cout(Xd_0__inst_mult_1_56 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_659 ),
	.datab(!Xd_0__inst_mult_0_664 ),
	.datac(!din_a[9]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_464 ),
	.cout(Xd_0__inst_mult_0_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_65 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_56 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_65_sumout ),
	.cout(Xd_0__inst_mult_0_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_659 ),
	.datab(!Xd_0__inst_mult_3_664 ),
	.datac(!din_a[45]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_464 ),
	.cout(Xd_0__inst_mult_3_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_75 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_75_sumout ),
	.cout(Xd_0__inst_mult_3_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_704 ),
	.datab(!Xd_0__inst_mult_2_709 ),
	.datac(!din_a[33]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_509 ),
	.cout(Xd_0__inst_mult_2_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_65 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_65_sumout ),
	.cout(Xd_0__inst_mult_2_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_679 ),
	.datab(!Xd_0__inst_mult_29_80_sumout ),
	.datac(!Xd_0__inst_mult_29_669 ),
	.datad(!Xd_0__inst_mult_29_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_499 ),
	.cout(Xd_0__inst_mult_29_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_70 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[356]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_70_sumout ),
	.cout(Xd_0__inst_mult_29_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_669 ),
	.datab(!Xd_0__inst_mult_28_80_sumout ),
	.datac(!Xd_0__inst_mult_28_659 ),
	.datad(!Xd_0__inst_mult_28_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_469 ),
	.cout(Xd_0__inst_mult_28_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_70 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[344]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_70_sumout ),
	.cout(Xd_0__inst_mult_28_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_669 ),
	.datab(!Xd_0__inst_mult_31_80_sumout ),
	.datac(!Xd_0__inst_mult_31_659 ),
	.datad(!Xd_0__inst_mult_31_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_469 ),
	.cout(Xd_0__inst_mult_31_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_60 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[380]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_60_sumout ),
	.cout(Xd_0__inst_mult_31_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_669 ),
	.datab(!Xd_0__inst_mult_30_80_sumout ),
	.datac(!Xd_0__inst_mult_30_659 ),
	.datad(!Xd_0__inst_mult_30_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_469 ),
	.cout(Xd_0__inst_mult_30_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_70 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[368]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_70_sumout ),
	.cout(Xd_0__inst_mult_30_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_150 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_694 ),
	.datab(!Xd_0__inst_mult_25_40_sumout ),
	.datac(!Xd_0__inst_mult_25_684 ),
	.datad(!Xd_0__inst_mult_25_689 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_544 ),
	.cout(Xd_0__inst_mult_25_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_75 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[308]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_75_sumout ),
	.cout(Xd_0__inst_mult_25_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_70 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[296]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_70_sumout ),
	.cout(Xd_0__inst_mult_24_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_150 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_694 ),
	.datab(!Xd_0__inst_mult_27_40_sumout ),
	.datac(!Xd_0__inst_mult_27_684 ),
	.datad(!Xd_0__inst_mult_27_689 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_544 ),
	.cout(Xd_0__inst_mult_27_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_75 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[332]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_75_sumout ),
	.cout(Xd_0__inst_mult_27_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_70 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[320]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_70_sumout ),
	.cout(Xd_0__inst_mult_26_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_679 ),
	.datab(!Xd_0__inst_mult_21_80_sumout ),
	.datac(!Xd_0__inst_mult_21_669 ),
	.datad(!Xd_0__inst_mult_21_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_499 ),
	.cout(Xd_0__inst_mult_21_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_65 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[260]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_65_sumout ),
	.cout(Xd_0__inst_mult_21_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_679 ),
	.datab(!Xd_0__inst_mult_20_40_sumout ),
	.datac(!Xd_0__inst_mult_20_669 ),
	.datad(!Xd_0__inst_mult_20_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_499 ),
	.cout(Xd_0__inst_mult_20_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_75 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[248]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_75_sumout ),
	.cout(Xd_0__inst_mult_20_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_679 ),
	.datab(!Xd_0__inst_mult_23_80_sumout ),
	.datac(!Xd_0__inst_mult_23_669 ),
	.datad(!Xd_0__inst_mult_23_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_499 ),
	.cout(Xd_0__inst_mult_23_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_60 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[284]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_60_sumout ),
	.cout(Xd_0__inst_mult_23_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_679 ),
	.datab(!Xd_0__inst_mult_22_80_sumout ),
	.datac(!Xd_0__inst_mult_22_669 ),
	.datad(!Xd_0__inst_mult_22_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_499 ),
	.cout(Xd_0__inst_mult_22_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_65 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[272]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_65_sumout ),
	.cout(Xd_0__inst_mult_22_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_679 ),
	.datab(!Xd_0__inst_mult_17_80_sumout ),
	.datac(!Xd_0__inst_mult_17_669 ),
	.datad(!Xd_0__inst_mult_17_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_499 ),
	.cout(Xd_0__inst_mult_17_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_70 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[212]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_70_sumout ),
	.cout(Xd_0__inst_mult_17_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_679 ),
	.datab(!Xd_0__inst_mult_16_75_sumout ),
	.datac(!Xd_0__inst_mult_16_669 ),
	.datad(!Xd_0__inst_mult_16_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_499 ),
	.cout(Xd_0__inst_mult_16_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_60 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[200]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_60_sumout ),
	.cout(Xd_0__inst_mult_16_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_141 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_679 ),
	.datab(!Xd_0__inst_mult_19_75_sumout ),
	.datac(!Xd_0__inst_mult_19_669 ),
	.datad(!Xd_0__inst_mult_19_674 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_499 ),
	.cout(Xd_0__inst_mult_19_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_65 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[236]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_65_sumout ),
	.cout(Xd_0__inst_mult_19_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_664 ),
	.datab(!Xd_0__inst_mult_18_75_sumout ),
	.datac(!Xd_0__inst_mult_18_654 ),
	.datad(!Xd_0__inst_mult_18_659 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_459 ),
	.cout(Xd_0__inst_mult_18_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_669 ),
	.datab(!Xd_0__inst_mult_13_75_sumout ),
	.datac(!Xd_0__inst_mult_13_659 ),
	.datad(!Xd_0__inst_mult_13_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_469 ),
	.cout(Xd_0__inst_mult_13_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_65 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[164]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_65_sumout ),
	.cout(Xd_0__inst_mult_13_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_664 ),
	.datab(!Xd_0__inst_mult_12_80_sumout ),
	.datac(!Xd_0__inst_mult_12_654 ),
	.datad(!Xd_0__inst_mult_12_659 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_459 ),
	.cout(Xd_0__inst_mult_12_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_60 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[152]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_60_sumout ),
	.cout(Xd_0__inst_mult_12_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_664 ),
	.datab(!Xd_0__inst_mult_15_50_sumout ),
	.datac(!Xd_0__inst_mult_15_654 ),
	.datad(!Xd_0__inst_mult_15_659 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_459 ),
	.cout(Xd_0__inst_mult_15_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_80 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_80_sumout ),
	.cout(Xd_0__inst_mult_15_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_133 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_664 ),
	.datab(!Xd_0__inst_mult_14_35_sumout ),
	.datac(!Xd_0__inst_mult_14_654 ),
	.datad(!Xd_0__inst_mult_14_659 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_459 ),
	.cout(Xd_0__inst_mult_14_460 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_60 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[176]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_60_sumout ),
	.cout(Xd_0__inst_mult_14_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_669 ),
	.datab(!Xd_0__inst_mult_9_75_sumout ),
	.datac(!Xd_0__inst_mult_9_659 ),
	.datad(!Xd_0__inst_mult_9_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_469 ),
	.cout(Xd_0__inst_mult_9_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_70 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_70_sumout ),
	.cout(Xd_0__inst_mult_9_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_669 ),
	.datab(!Xd_0__inst_mult_8_50_sumout ),
	.datac(!Xd_0__inst_mult_8_659 ),
	.datad(!Xd_0__inst_mult_8_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_469 ),
	.cout(Xd_0__inst_mult_8_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_80 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[104]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_80_sumout ),
	.cout(Xd_0__inst_mult_8_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_669 ),
	.datab(!Xd_0__inst_mult_11_75_sumout ),
	.datac(!Xd_0__inst_mult_11_659 ),
	.datad(!Xd_0__inst_mult_11_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_469 ),
	.cout(Xd_0__inst_mult_11_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_60 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[140]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_60_sumout ),
	.cout(Xd_0__inst_mult_11_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_669 ),
	.datab(!Xd_0__inst_mult_10_50_sumout ),
	.datac(!Xd_0__inst_mult_10_659 ),
	.datad(!Xd_0__inst_mult_10_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_469 ),
	.cout(Xd_0__inst_mult_10_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_75 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[128]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_75_sumout ),
	.cout(Xd_0__inst_mult_10_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_669 ),
	.datab(!Xd_0__inst_mult_5_45_sumout ),
	.datac(!Xd_0__inst_mult_5_659 ),
	.datad(!Xd_0__inst_mult_5_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_469 ),
	.cout(Xd_0__inst_mult_5_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_80 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_80_sumout ),
	.cout(Xd_0__inst_mult_5_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_669 ),
	.datab(!Xd_0__inst_mult_4_75_sumout ),
	.datac(!Xd_0__inst_mult_4_659 ),
	.datad(!Xd_0__inst_mult_4_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_469 ),
	.cout(Xd_0__inst_mult_4_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_60 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_60_sumout ),
	.cout(Xd_0__inst_mult_4_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_669 ),
	.datab(!Xd_0__inst_mult_7_50_sumout ),
	.datac(!Xd_0__inst_mult_7_659 ),
	.datad(!Xd_0__inst_mult_7_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_469 ),
	.cout(Xd_0__inst_mult_7_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_75 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_75_sumout ),
	.cout(Xd_0__inst_mult_7_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_669 ),
	.datab(!Xd_0__inst_mult_6_45_sumout ),
	.datac(!Xd_0__inst_mult_6_659 ),
	.datad(!Xd_0__inst_mult_6_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_469 ),
	.cout(Xd_0__inst_mult_6_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_75 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_75_sumout ),
	.cout(Xd_0__inst_mult_6_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_669 ),
	.datab(!Xd_0__inst_mult_1_75_sumout ),
	.datac(!Xd_0__inst_mult_1_659 ),
	.datad(!Xd_0__inst_mult_1_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_469 ),
	.cout(Xd_0__inst_mult_1_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_60 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_60_sumout ),
	.cout(Xd_0__inst_mult_1_61 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_669 ),
	.datab(!Xd_0__inst_mult_0_50_sumout ),
	.datac(!Xd_0__inst_mult_0_659 ),
	.datad(!Xd_0__inst_mult_0_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_469 ),
	.cout(Xd_0__inst_mult_0_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_70 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_61 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_70_sumout ),
	.cout(Xd_0__inst_mult_0_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_669 ),
	.datab(!Xd_0__inst_mult_3_45_sumout ),
	.datac(!Xd_0__inst_mult_3_659 ),
	.datad(!Xd_0__inst_mult_3_664 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_469 ),
	.cout(Xd_0__inst_mult_3_470 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_80 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_80_sumout ),
	.cout(Xd_0__inst_mult_3_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_144 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_714 ),
	.datab(!Xd_0__inst_mult_2_45_sumout ),
	.datac(!Xd_0__inst_mult_2_704 ),
	.datad(!Xd_0__inst_mult_2_709 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_514 ),
	.cout(Xd_0__inst_mult_2_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_70 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_70_sumout ),
	.cout(Xd_0__inst_mult_2_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_29_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_684 ),
	.datab(!Xd_0__inst_mult_29_50_sumout ),
	.datac(!Xd_0__inst_mult_29_679 ),
	.datad(!Xd_0__inst_mult_29_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_504 ),
	.cout(Xd_0__inst_mult_29_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_75 (
// Equation(s):

	.dataa(!din_a[358]),
	.datab(!din_b[357]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_75_sumout ),
	.cout(Xd_0__inst_mult_29_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_28_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_674 ),
	.datab(!Xd_0__inst_mult_28_45_sumout ),
	.datac(!Xd_0__inst_mult_28_669 ),
	.datad(!Xd_0__inst_mult_28_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_474 ),
	.cout(Xd_0__inst_mult_28_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_75 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[345]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_75_sumout ),
	.cout(Xd_0__inst_mult_28_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_31_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_674 ),
	.datab(!Xd_0__inst_mult_31_75_sumout ),
	.datac(!Xd_0__inst_mult_31_669 ),
	.datad(!Xd_0__inst_mult_31_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_474 ),
	.cout(Xd_0__inst_mult_31_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_65 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[381]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_65_sumout ),
	.cout(Xd_0__inst_mult_31_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_30_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_674 ),
	.datab(!Xd_0__inst_mult_30_50_sumout ),
	.datac(!Xd_0__inst_mult_30_669 ),
	.datad(!Xd_0__inst_mult_30_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_474 ),
	.cout(Xd_0__inst_mult_30_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_75 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[369]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_75_sumout ),
	.cout(Xd_0__inst_mult_30_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_25_151 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_699 ),
	.datab(!Xd_0__inst_mult_25_55_sumout ),
	.datac(!Xd_0__inst_mult_25_694 ),
	.datad(!Xd_0__inst_mult_25_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_549 ),
	.cout(Xd_0__inst_mult_25_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_80 (
// Equation(s):

	.dataa(!din_a[310]),
	.datab(!din_b[309]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_80_sumout ),
	.cout(Xd_0__inst_mult_25_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_75 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[297]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_75_sumout ),
	.cout(Xd_0__inst_mult_24_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_27_151 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_699 ),
	.datab(!Xd_0__inst_mult_27_35_sumout ),
	.datac(!Xd_0__inst_mult_27_694 ),
	.datad(!Xd_0__inst_mult_27_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_549 ),
	.cout(Xd_0__inst_mult_27_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_80 (
// Equation(s):

	.dataa(!din_a[334]),
	.datab(!din_b[333]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_80_sumout ),
	.cout(Xd_0__inst_mult_27_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_75 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[321]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_75_sumout ),
	.cout(Xd_0__inst_mult_26_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_21_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_684 ),
	.datab(!Xd_0__inst_mult_21_75_sumout ),
	.datac(!Xd_0__inst_mult_21_679 ),
	.datad(!Xd_0__inst_mult_21_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_504 ),
	.cout(Xd_0__inst_mult_21_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_70 (
// Equation(s):

	.dataa(!din_a[262]),
	.datab(!din_b[261]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_70_sumout ),
	.cout(Xd_0__inst_mult_21_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_20_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_684 ),
	.datab(!Xd_0__inst_mult_20_60_sumout ),
	.datac(!Xd_0__inst_mult_20_679 ),
	.datad(!Xd_0__inst_mult_20_40_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_504 ),
	.cout(Xd_0__inst_mult_20_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_80 (
// Equation(s):

	.dataa(!din_a[250]),
	.datab(!din_b[249]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_80_sumout ),
	.cout(Xd_0__inst_mult_20_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_23_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_684 ),
	.datab(!Xd_0__inst_mult_23_75_sumout ),
	.datac(!Xd_0__inst_mult_23_679 ),
	.datad(!Xd_0__inst_mult_23_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_504 ),
	.cout(Xd_0__inst_mult_23_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_65 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[285]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_65_sumout ),
	.cout(Xd_0__inst_mult_23_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_22_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_684 ),
	.datab(!Xd_0__inst_mult_22_75_sumout ),
	.datac(!Xd_0__inst_mult_22_679 ),
	.datad(!Xd_0__inst_mult_22_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_504 ),
	.cout(Xd_0__inst_mult_22_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_70 (
// Equation(s):

	.dataa(!din_a[274]),
	.datab(!din_b[273]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_70_sumout ),
	.cout(Xd_0__inst_mult_22_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_17_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_684 ),
	.datab(!Xd_0__inst_mult_17_60_sumout ),
	.datac(!Xd_0__inst_mult_17_679 ),
	.datad(!Xd_0__inst_mult_17_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_504 ),
	.cout(Xd_0__inst_mult_17_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_75 (
// Equation(s):

	.dataa(!din_a[214]),
	.datab(!din_b[213]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_75_sumout ),
	.cout(Xd_0__inst_mult_17_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_16_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_684 ),
	.datab(!Xd_0__inst_mult_16_80_sumout ),
	.datac(!Xd_0__inst_mult_16_679 ),
	.datad(!Xd_0__inst_mult_16_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_504 ),
	.cout(Xd_0__inst_mult_16_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_65 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[201]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_65_sumout ),
	.cout(Xd_0__inst_mult_16_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_19_142 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_684 ),
	.datab(!Xd_0__inst_mult_19_80_sumout ),
	.datac(!Xd_0__inst_mult_19_679 ),
	.datad(!Xd_0__inst_mult_19_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_504 ),
	.cout(Xd_0__inst_mult_19_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_70 (
// Equation(s):

	.dataa(!din_a[238]),
	.datab(!din_b[237]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_66 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_70_sumout ),
	.cout(Xd_0__inst_mult_19_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_18_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_669 ),
	.datab(!Xd_0__inst_mult_18_80_sumout ),
	.datac(!Xd_0__inst_mult_18_664 ),
	.datad(!Xd_0__inst_mult_18_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_464 ),
	.cout(Xd_0__inst_mult_18_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_70 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[225]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_70_sumout ),
	.cout(Xd_0__inst_mult_18_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_13_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_674 ),
	.datab(!Xd_0__inst_mult_13_80_sumout ),
	.datac(!Xd_0__inst_mult_13_669 ),
	.datad(!Xd_0__inst_mult_13_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_474 ),
	.cout(Xd_0__inst_mult_13_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_70 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_70_sumout ),
	.cout(Xd_0__inst_mult_13_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_12_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_669 ),
	.datab(!Xd_0__inst_mult_12_75_sumout ),
	.datac(!Xd_0__inst_mult_12_664 ),
	.datad(!Xd_0__inst_mult_12_80_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_464 ),
	.cout(Xd_0__inst_mult_12_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_15_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_669 ),
	.datab(!Xd_0__inst_mult_15_60_sumout ),
	.datac(!Xd_0__inst_mult_15_664 ),
	.datad(!Xd_0__inst_mult_15_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_464 ),
	.cout(Xd_0__inst_mult_15_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_14_134 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_669 ),
	.datab(!Xd_0__inst_mult_14_80_sumout ),
	.datac(!Xd_0__inst_mult_14_664 ),
	.datad(!Xd_0__inst_mult_14_35_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_464 ),
	.cout(Xd_0__inst_mult_14_465 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_65 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[177]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_65_sumout ),
	.cout(Xd_0__inst_mult_14_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_9_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_674 ),
	.datab(!Xd_0__inst_mult_9_80_sumout ),
	.datac(!Xd_0__inst_mult_9_669 ),
	.datad(!Xd_0__inst_mult_9_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_474 ),
	.cout(Xd_0__inst_mult_9_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_8_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_674 ),
	.datab(!Xd_0__inst_mult_8_65_sumout ),
	.datac(!Xd_0__inst_mult_8_669 ),
	.datad(!Xd_0__inst_mult_8_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_474 ),
	.cout(Xd_0__inst_mult_8_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_11_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_674 ),
	.datab(!Xd_0__inst_mult_11_80_sumout ),
	.datac(!Xd_0__inst_mult_11_669 ),
	.datad(!Xd_0__inst_mult_11_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_474 ),
	.cout(Xd_0__inst_mult_11_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_65 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[141]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_65_sumout ),
	.cout(Xd_0__inst_mult_11_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_10_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_674 ),
	.datab(!Xd_0__inst_mult_10_80_sumout ),
	.datac(!Xd_0__inst_mult_10_669 ),
	.datad(!Xd_0__inst_mult_10_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_474 ),
	.cout(Xd_0__inst_mult_10_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_5_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_674 ),
	.datab(!Xd_0__inst_mult_5_75_sumout ),
	.datac(!Xd_0__inst_mult_5_669 ),
	.datad(!Xd_0__inst_mult_5_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_474 ),
	.cout(Xd_0__inst_mult_5_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_4_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_674 ),
	.datab(!Xd_0__inst_mult_4_80_sumout ),
	.datac(!Xd_0__inst_mult_4_669 ),
	.datad(!Xd_0__inst_mult_4_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_474 ),
	.cout(Xd_0__inst_mult_4_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_65 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_65_sumout ),
	.cout(Xd_0__inst_mult_4_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_7_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_674 ),
	.datab(!Xd_0__inst_mult_7_80_sumout ),
	.datac(!Xd_0__inst_mult_7_669 ),
	.datad(!Xd_0__inst_mult_7_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_474 ),
	.cout(Xd_0__inst_mult_7_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_6_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_674 ),
	.datab(!Xd_0__inst_mult_6_80_sumout ),
	.datac(!Xd_0__inst_mult_6_669 ),
	.datad(!Xd_0__inst_mult_6_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_474 ),
	.cout(Xd_0__inst_mult_6_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_1_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_674 ),
	.datab(!Xd_0__inst_mult_1_80_sumout ),
	.datac(!Xd_0__inst_mult_1_669 ),
	.datad(!Xd_0__inst_mult_1_75_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_474 ),
	.cout(Xd_0__inst_mult_1_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_65 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_65_sumout ),
	.cout(Xd_0__inst_mult_1_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_0_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_674 ),
	.datab(!Xd_0__inst_mult_0_80_sumout ),
	.datac(!Xd_0__inst_mult_0_669 ),
	.datad(!Xd_0__inst_mult_0_50_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_474 ),
	.cout(Xd_0__inst_mult_0_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_3_136 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_674 ),
	.datab(!Xd_0__inst_mult_3_60_sumout ),
	.datac(!Xd_0__inst_mult_3_669 ),
	.datad(!Xd_0__inst_mult_3_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_470 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_474 ),
	.cout(Xd_0__inst_mult_3_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000066669),
	.shared_arith("off")
) Xd_0__inst_mult_2_145 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_719 ),
	.datab(!Xd_0__inst_mult_2_80_sumout ),
	.datac(!Xd_0__inst_mult_2_714 ),
	.datad(!Xd_0__inst_mult_2_45_sumout ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_519 ),
	.cout(Xd_0__inst_mult_2_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_75 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_75_sumout ),
	.cout(Xd_0__inst_mult_2_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_29_684 ),
	.datab(!Xd_0__inst_mult_29_50_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_28_674 ),
	.datab(!Xd_0__inst_mult_28_45_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_31_674 ),
	.datab(!Xd_0__inst_mult_31_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_70 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[382]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_70_sumout ),
	.cout(Xd_0__inst_mult_31_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_30_674 ),
	.datab(!Xd_0__inst_mult_30_50_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_152 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_25_699 ),
	.datab(!Xd_0__inst_mult_25_55_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_554 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_24_80 (
// Equation(s):

	.dataa(!din_a[298]),
	.datab(!din_b[298]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_80_sumout ),
	.cout(Xd_0__inst_mult_24_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_152 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_27_699 ),
	.datab(!Xd_0__inst_mult_27_35_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_554 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_26_80 (
// Equation(s):

	.dataa(!din_a[322]),
	.datab(!din_b[322]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_80_sumout ),
	.cout(Xd_0__inst_mult_26_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_21_684 ),
	.datab(!Xd_0__inst_mult_21_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_20_684 ),
	.datab(!Xd_0__inst_mult_20_60_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_23_684 ),
	.datab(!Xd_0__inst_mult_23_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_70 (
// Equation(s):

	.dataa(!din_a[286]),
	.datab(!din_b[286]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_70_sumout ),
	.cout(Xd_0__inst_mult_23_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_22_684 ),
	.datab(!Xd_0__inst_mult_22_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_17_684 ),
	.datab(!Xd_0__inst_mult_17_60_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_16_684 ),
	.datab(!Xd_0__inst_mult_16_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_70 (
// Equation(s):

	.dataa(!din_a[202]),
	.datab(!din_b[202]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_70_sumout ),
	.cout(Xd_0__inst_mult_16_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_143 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_19_684 ),
	.datab(!Xd_0__inst_mult_19_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_509 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_18_669 ),
	.datab(!Xd_0__inst_mult_18_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_469 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_13_674 ),
	.datab(!Xd_0__inst_mult_13_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_12_669 ),
	.datab(!Xd_0__inst_mult_12_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_469 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_65 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_65_sumout ),
	.cout(Xd_0__inst_mult_12_66 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_15_669 ),
	.datab(!Xd_0__inst_mult_15_60_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_469 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_135 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_14_669 ),
	.datab(!Xd_0__inst_mult_14_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_465 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_469 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_70 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_70_sumout ),
	.cout(Xd_0__inst_mult_14_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_9_674 ),
	.datab(!Xd_0__inst_mult_9_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_8_674 ),
	.datab(!Xd_0__inst_mult_8_65_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_11_674 ),
	.datab(!Xd_0__inst_mult_11_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_70 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_70_sumout ),
	.cout(Xd_0__inst_mult_11_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_10_674 ),
	.datab(!Xd_0__inst_mult_10_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_5_674 ),
	.datab(!Xd_0__inst_mult_5_75_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_4_674 ),
	.datab(!Xd_0__inst_mult_4_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_70 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_70_sumout ),
	.cout(Xd_0__inst_mult_4_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_7_674 ),
	.datab(!Xd_0__inst_mult_7_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_6_674 ),
	.datab(!Xd_0__inst_mult_6_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_1_674 ),
	.datab(!Xd_0__inst_mult_1_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_70 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_70_sumout ),
	.cout(Xd_0__inst_mult_1_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_0_674 ),
	.datab(!Xd_0__inst_mult_0_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_75 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_75_sumout ),
	.cout(Xd_0__inst_mult_0_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_137 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_3_674 ),
	.datab(!Xd_0__inst_mult_3_60_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_479 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_146 (
// Equation(s):

	.dataa(!Xd_0__inst_mult_2_719 ),
	.datab(!Xd_0__inst_mult_2_80_sumout ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_524 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_139 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[111]),
	.datac(!Xd_0__inst_mult_9_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_489 ),
	.cout(Xd_0__inst_mult_9_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_139 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[99]),
	.datac(!Xd_0__inst_mult_8_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_489 ),
	.cout(Xd_0__inst_mult_8_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_144 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[255]),
	.datac(!din_a[259]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_514 ),
	.cout(Xd_0__inst_mult_21_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_145 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_519 ),
	.cout(Xd_0__inst_mult_21_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_146 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[253]),
	.datac(!din_a[262]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_524 ),
	.cout(Xd_0__inst_mult_21_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_139 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[135]),
	.datac(!Xd_0__inst_mult_11_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_489 ),
	.cout(Xd_0__inst_mult_11_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_139 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[123]),
	.datac(!Xd_0__inst_mult_10_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_489 ),
	.cout(Xd_0__inst_mult_10_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_144 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[243]),
	.datac(!din_a[247]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_514 ),
	.cout(Xd_0__inst_mult_20_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_145 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_519 ),
	.cout(Xd_0__inst_mult_20_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_146 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[241]),
	.datac(!din_a[250]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_524 ),
	.cout(Xd_0__inst_mult_20_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_153 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[303]),
	.datac(!din_a[304]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_559 ),
	.cout(Xd_0__inst_mult_25_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_154 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_564 ),
	.cout(Xd_0__inst_mult_25_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_155 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[301]),
	.datac(!din_a[307]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_569 ),
	.cout(Xd_0__inst_mult_25_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_139 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[39]),
	.datac(!Xd_0__inst_mult_3_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_489 ),
	.cout(Xd_0__inst_mult_3_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_70 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[148]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_46 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_70_sumout ),
	.cout(Xd_0__inst_mult_12_71 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_139 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[3]),
	.datac(!Xd_0__inst_mult_0_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_489 ),
	.cout(Xd_0__inst_mult_0_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_144 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[279]),
	.datac(!din_a[283]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_514 ),
	.cout(Xd_0__inst_mult_23_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_145 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_519 ),
	.cout(Xd_0__inst_mult_23_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_146 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[277]),
	.datac(!din_a[286]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_524 ),
	.cout(Xd_0__inst_mult_23_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_139 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[75]),
	.datac(!Xd_0__inst_mult_6_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_489 ),
	.cout(Xd_0__inst_mult_6_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_139 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[15]),
	.datac(!Xd_0__inst_mult_1_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_489 ),
	.cout(Xd_0__inst_mult_1_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_144 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[267]),
	.datac(!din_a[271]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_514 ),
	.cout(Xd_0__inst_mult_22_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_145 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_519 ),
	.cout(Xd_0__inst_mult_22_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_146 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[265]),
	.datac(!din_a[274]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_524 ),
	.cout(Xd_0__inst_mult_22_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_181 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[291]),
	.datac(!din_a[292]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_699 ),
	.cout(Xd_0__inst_mult_24_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_182 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_704 ),
	.cout(Xd_0__inst_mult_24_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_183 (
// Equation(s):

	.dataa(!din_a[294]),
	.datab(!din_b[289]),
	.datac(!din_a[295]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_709 ),
	.cout(Xd_0__inst_mult_24_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_181 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[321]),
	.datac(!din_a[313]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_699 ),
	.cout(Xd_0__inst_mult_26_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_182 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[318]),
	.datac(!din_a[316]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_704 ),
	.cout(Xd_0__inst_mult_26_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_183 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_709 ),
	.cout(Xd_0__inst_mult_26_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_139 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[87]),
	.datac(!Xd_0__inst_mult_7_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_489 ),
	.cout(Xd_0__inst_mult_7_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_139 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[51]),
	.datac(!Xd_0__inst_mult_4_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_489 ),
	.cout(Xd_0__inst_mult_4_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_144 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[231]),
	.datac(!din_a[235]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_514 ),
	.cout(Xd_0__inst_mult_19_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_145 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_519 ),
	.cout(Xd_0__inst_mult_19_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_146 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[229]),
	.datac(!din_a[238]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_524 ),
	.cout(Xd_0__inst_mult_19_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_139 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[363]),
	.datac(!Xd_0__inst_mult_30_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_489 ),
	.cout(Xd_0__inst_mult_30_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_139 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[63]),
	.datac(!Xd_0__inst_mult_5_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_489 ),
	.cout(Xd_0__inst_mult_5_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_144 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[207]),
	.datac(!din_a[211]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_514 ),
	.cout(Xd_0__inst_mult_17_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_145 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_519 ),
	.cout(Xd_0__inst_mult_17_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_146 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[205]),
	.datac(!din_a[214]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_524 ),
	.cout(Xd_0__inst_mult_17_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_153 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[327]),
	.datac(!din_a[328]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_559 ),
	.cout(Xd_0__inst_mult_27_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_154 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_564 ),
	.cout(Xd_0__inst_mult_27_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_155 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[325]),
	.datac(!din_a[331]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_569 ),
	.cout(Xd_0__inst_mult_27_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_139 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[159]),
	.datac(!Xd_0__inst_mult_13_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_489 ),
	.cout(Xd_0__inst_mult_13_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_147 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_529 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_148 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[27]),
	.datac(!Xd_0__inst_mult_2_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_534 ),
	.cout(Xd_0__inst_mult_2_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_149 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_539 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_144 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[195]),
	.datac(!din_a[199]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_514 ),
	.cout(Xd_0__inst_mult_16_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_145 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_519 ),
	.cout(Xd_0__inst_mult_16_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_146 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[193]),
	.datac(!din_a[202]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_524 ),
	.cout(Xd_0__inst_mult_16_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_139 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[339]),
	.datac(!Xd_0__inst_mult_28_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_489 ),
	.cout(Xd_0__inst_mult_28_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_138 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_484 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_139 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[375]),
	.datac(!Xd_0__inst_mult_31_679 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_489 ),
	.cout(Xd_0__inst_mult_31_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_140 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_494 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_144 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[351]),
	.datac(!din_a[355]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_514 ),
	.cout(Xd_0__inst_mult_29_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_145 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_519 ),
	.cout(Xd_0__inst_mult_29_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_146 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[349]),
	.datac(!din_a[358]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_524 ),
	.cout(Xd_0__inst_mult_29_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_184 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[315]),
	.datac(!din_a[316]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_714 ),
	.cout(Xd_0__inst_mult_26_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_185 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_719 ),
	.cout(Xd_0__inst_mult_26_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_186 (
// Equation(s):

	.dataa(!din_a[318]),
	.datab(!din_b[313]),
	.datac(!din_a[319]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_724 ),
	.cout(Xd_0__inst_mult_26_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_184 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[297]),
	.datac(!din_a[289]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_714 ),
	.cout(Xd_0__inst_mult_24_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_185 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[294]),
	.datac(!din_a[292]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_719 ),
	.cout(Xd_0__inst_mult_24_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_186 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_724 ),
	.cout(Xd_0__inst_mult_24_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_75 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[274]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_75_sumout ),
	.cout(Xd_0__inst_mult_22_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_75 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_75_sumout ),
	.cout(Xd_0__inst_mult_12_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_80 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_80_sumout ),
	.cout(Xd_0__inst_mult_10_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_80 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_80_sumout ),
	.cout(Xd_0__inst_mult_0_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_147 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[349]),
	.datac(!din_a[353]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_529 ),
	.cout(Xd_0__inst_mult_29_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_148 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_534 ),
	.cout(Xd_0__inst_mult_29_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_141 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[337]),
	.datac(!din_a[341]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_499 ),
	.cout(Xd_0__inst_mult_28_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_142 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_504 ),
	.cout(Xd_0__inst_mult_28_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_141 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[373]),
	.datac(!din_a[377]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_499 ),
	.cout(Xd_0__inst_mult_31_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_142 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_504 ),
	.cout(Xd_0__inst_mult_31_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_141 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[361]),
	.datac(!din_a[365]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_499 ),
	.cout(Xd_0__inst_mult_30_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_142 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_504 ),
	.cout(Xd_0__inst_mult_30_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_75 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[262]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_75_sumout ),
	.cout(Xd_0__inst_mult_21_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_156 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[301]),
	.datac(!din_a[305]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_574 ),
	.cout(Xd_0__inst_mult_25_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_157 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_579 ),
	.cout(Xd_0__inst_mult_25_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_187 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[289]),
	.datac(!din_a[293]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_729 ),
	.cout(Xd_0__inst_mult_24_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_188 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_734 ),
	.cout(Xd_0__inst_mult_24_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_75 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[382]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_75_sumout ),
	.cout(Xd_0__inst_mult_31_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_156 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[325]),
	.datac(!din_a[329]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_455 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_574 ),
	.cout(Xd_0__inst_mult_27_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_157 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_579 ),
	.cout(Xd_0__inst_mult_27_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_75 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[286]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_75_sumout ),
	.cout(Xd_0__inst_mult_23_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_187 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[313]),
	.datac(!din_a[317]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_729 ),
	.cout(Xd_0__inst_mult_26_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_188 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_734 ),
	.cout(Xd_0__inst_mult_26_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_75 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_75_sumout ),
	.cout(Xd_0__inst_mult_1_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_147 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[253]),
	.datac(!din_a[257]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_529 ),
	.cout(Xd_0__inst_mult_21_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_148 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_534 ),
	.cout(Xd_0__inst_mult_21_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_75 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[57]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_75_sumout ),
	.cout(Xd_0__inst_mult_4_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_147 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[241]),
	.datac(!din_a[245]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_529 ),
	.cout(Xd_0__inst_mult_20_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_148 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_534 ),
	.cout(Xd_0__inst_mult_20_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_147 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[277]),
	.datac(!din_a[281]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_529 ),
	.cout(Xd_0__inst_mult_23_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_148 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_534 ),
	.cout(Xd_0__inst_mult_23_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_80 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_80_sumout ),
	.cout(Xd_0__inst_mult_2_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_147 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[265]),
	.datac(!din_a[269]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_529 ),
	.cout(Xd_0__inst_mult_22_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_148 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_534 ),
	.cout(Xd_0__inst_mult_22_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_147 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[205]),
	.datac(!din_a[209]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_529 ),
	.cout(Xd_0__inst_mult_17_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_148 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_534 ),
	.cout(Xd_0__inst_mult_17_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_75 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[141]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_75_sumout ),
	.cout(Xd_0__inst_mult_11_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_147 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[193]),
	.datac(!din_a[197]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_529 ),
	.cout(Xd_0__inst_mult_16_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_148 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_534 ),
	.cout(Xd_0__inst_mult_16_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_147 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[229]),
	.datac(!din_a[233]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_395 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_529 ),
	.cout(Xd_0__inst_mult_19_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_148 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_534 ),
	.cout(Xd_0__inst_mult_19_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_136 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[217]),
	.datac(!din_a[221]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_474 ),
	.cout(Xd_0__inst_mult_18_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_137 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_674 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_479 ),
	.cout(Xd_0__inst_mult_18_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_141 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[157]),
	.datac(!din_a[161]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_499 ),
	.cout(Xd_0__inst_mult_13_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_142 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_504 ),
	.cout(Xd_0__inst_mult_13_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_136 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[145]),
	.datac(!din_a[149]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_474 ),
	.cout(Xd_0__inst_mult_12_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_137 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_674 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_479 ),
	.cout(Xd_0__inst_mult_12_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_136 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[181]),
	.datac(!din_a[185]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_474 ),
	.cout(Xd_0__inst_mult_15_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_137 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_674 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_479 ),
	.cout(Xd_0__inst_mult_15_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_136 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[169]),
	.datac(!din_a[173]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_330 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_474 ),
	.cout(Xd_0__inst_mult_14_475 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_137 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_674 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_479 ),
	.cout(Xd_0__inst_mult_14_480 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_141 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[109]),
	.datac(!din_a[113]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_499 ),
	.cout(Xd_0__inst_mult_9_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_142 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_504 ),
	.cout(Xd_0__inst_mult_9_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_141 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[97]),
	.datac(!din_a[101]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_499 ),
	.cout(Xd_0__inst_mult_8_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_142 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_504 ),
	.cout(Xd_0__inst_mult_8_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_141 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[133]),
	.datac(!din_a[137]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_499 ),
	.cout(Xd_0__inst_mult_11_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_142 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_504 ),
	.cout(Xd_0__inst_mult_11_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_141 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[121]),
	.datac(!din_a[125]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_499 ),
	.cout(Xd_0__inst_mult_10_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_142 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_504 ),
	.cout(Xd_0__inst_mult_10_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_141 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[61]),
	.datac(!din_a[65]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_499 ),
	.cout(Xd_0__inst_mult_5_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_142 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_504 ),
	.cout(Xd_0__inst_mult_5_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_141 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[49]),
	.datac(!din_a[53]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_499 ),
	.cout(Xd_0__inst_mult_4_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_142 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_504 ),
	.cout(Xd_0__inst_mult_4_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_141 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[85]),
	.datac(!din_a[89]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_499 ),
	.cout(Xd_0__inst_mult_7_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_142 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_504 ),
	.cout(Xd_0__inst_mult_7_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_141 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[73]),
	.datac(!din_a[77]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_499 ),
	.cout(Xd_0__inst_mult_6_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_142 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_504 ),
	.cout(Xd_0__inst_mult_6_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_141 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[13]),
	.datac(!din_a[17]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_499 ),
	.cout(Xd_0__inst_mult_1_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_142 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_504 ),
	.cout(Xd_0__inst_mult_1_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_141 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[1]),
	.datac(!din_a[5]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_499 ),
	.cout(Xd_0__inst_mult_0_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_142 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_504 ),
	.cout(Xd_0__inst_mult_0_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_141 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[37]),
	.datac(!din_a[41]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_355 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_499 ),
	.cout(Xd_0__inst_mult_3_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_142 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_504 ),
	.cout(Xd_0__inst_mult_3_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_150 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[25]),
	.datac(!din_a[29]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_415 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_544 ),
	.cout(Xd_0__inst_mult_2_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_151 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_549 ),
	.cout(Xd_0__inst_mult_2_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_149 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[349]),
	.datac(!din_a[354]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_539 ),
	.cout(Xd_0__inst_mult_29_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_150 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_544 ),
	.cout(Xd_0__inst_mult_29_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_143 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[337]),
	.datac(!din_a[342]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_509 ),
	.cout(Xd_0__inst_mult_28_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_144 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_514 ),
	.cout(Xd_0__inst_mult_28_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_143 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[373]),
	.datac(!din_a[378]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_509 ),
	.cout(Xd_0__inst_mult_31_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_144 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_514 ),
	.cout(Xd_0__inst_mult_31_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_143 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[361]),
	.datac(!din_a[366]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_509 ),
	.cout(Xd_0__inst_mult_30_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_144 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_514 ),
	.cout(Xd_0__inst_mult_30_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_158 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[301]),
	.datac(!din_a[306]),
	.datad(!din_b[300]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_584 ),
	.cout(Xd_0__inst_mult_25_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_159 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[302]),
	.datac(!Xd_0__inst_mult_25_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_589 ),
	.cout(Xd_0__inst_mult_25_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_189 (
// Equation(s):

	.dataa(!din_a[293]),
	.datab(!din_b[289]),
	.datac(!din_a[294]),
	.datad(!din_b[288]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_739 ),
	.cout(Xd_0__inst_mult_24_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_190 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[290]),
	.datac(!Xd_0__inst_mult_24_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_744 ),
	.cout(Xd_0__inst_mult_24_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_158 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[325]),
	.datac(!din_a[330]),
	.datad(!din_b[324]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_584 ),
	.cout(Xd_0__inst_mult_27_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_159 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[326]),
	.datac(!Xd_0__inst_mult_27_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_589 ),
	.cout(Xd_0__inst_mult_27_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_189 (
// Equation(s):

	.dataa(!din_a[317]),
	.datab(!din_b[313]),
	.datac(!din_a[318]),
	.datad(!din_b[312]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_739 ),
	.cout(Xd_0__inst_mult_26_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_190 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[314]),
	.datac(!Xd_0__inst_mult_26_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_744 ),
	.cout(Xd_0__inst_mult_26_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_149 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[253]),
	.datac(!din_a[258]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_539 ),
	.cout(Xd_0__inst_mult_21_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_150 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_544 ),
	.cout(Xd_0__inst_mult_21_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_149 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[241]),
	.datac(!din_a[246]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_539 ),
	.cout(Xd_0__inst_mult_20_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_150 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_544 ),
	.cout(Xd_0__inst_mult_20_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_149 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[277]),
	.datac(!din_a[282]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_539 ),
	.cout(Xd_0__inst_mult_23_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_150 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_544 ),
	.cout(Xd_0__inst_mult_23_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_149 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[265]),
	.datac(!din_a[270]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_539 ),
	.cout(Xd_0__inst_mult_22_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_150 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_544 ),
	.cout(Xd_0__inst_mult_22_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_149 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[205]),
	.datac(!din_a[210]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_539 ),
	.cout(Xd_0__inst_mult_17_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_150 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_544 ),
	.cout(Xd_0__inst_mult_17_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_149 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[193]),
	.datac(!din_a[198]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_539 ),
	.cout(Xd_0__inst_mult_16_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_150 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_544 ),
	.cout(Xd_0__inst_mult_16_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_149 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[229]),
	.datac(!din_a[234]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_539 ),
	.cout(Xd_0__inst_mult_19_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_150 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_544 ),
	.cout(Xd_0__inst_mult_19_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_138 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[217]),
	.datac(!din_a[222]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_484 ),
	.cout(Xd_0__inst_mult_18_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_139 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_489 ),
	.cout(Xd_0__inst_mult_18_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_143 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[157]),
	.datac(!din_a[162]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_509 ),
	.cout(Xd_0__inst_mult_13_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_144 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_514 ),
	.cout(Xd_0__inst_mult_13_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_138 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[145]),
	.datac(!din_a[150]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_484 ),
	.cout(Xd_0__inst_mult_12_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_139 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_489 ),
	.cout(Xd_0__inst_mult_12_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_138 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[181]),
	.datac(!din_a[186]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_484 ),
	.cout(Xd_0__inst_mult_15_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_139 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_489 ),
	.cout(Xd_0__inst_mult_15_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_138 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[169]),
	.datac(!din_a[174]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_475 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_484 ),
	.cout(Xd_0__inst_mult_14_485 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_139 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_684 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_480 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_489 ),
	.cout(Xd_0__inst_mult_14_490 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_143 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[109]),
	.datac(!din_a[114]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_509 ),
	.cout(Xd_0__inst_mult_9_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_144 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_514 ),
	.cout(Xd_0__inst_mult_9_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_143 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[97]),
	.datac(!din_a[102]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_509 ),
	.cout(Xd_0__inst_mult_8_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_144 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_514 ),
	.cout(Xd_0__inst_mult_8_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_143 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[133]),
	.datac(!din_a[138]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_509 ),
	.cout(Xd_0__inst_mult_11_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_144 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_514 ),
	.cout(Xd_0__inst_mult_11_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_143 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[121]),
	.datac(!din_a[126]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_509 ),
	.cout(Xd_0__inst_mult_10_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_144 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_514 ),
	.cout(Xd_0__inst_mult_10_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_143 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[61]),
	.datac(!din_a[66]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_509 ),
	.cout(Xd_0__inst_mult_5_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_144 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_514 ),
	.cout(Xd_0__inst_mult_5_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_143 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[49]),
	.datac(!din_a[54]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_509 ),
	.cout(Xd_0__inst_mult_4_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_144 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_514 ),
	.cout(Xd_0__inst_mult_4_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_143 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[85]),
	.datac(!din_a[90]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_509 ),
	.cout(Xd_0__inst_mult_7_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_144 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_514 ),
	.cout(Xd_0__inst_mult_7_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_143 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[73]),
	.datac(!din_a[78]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_509 ),
	.cout(Xd_0__inst_mult_6_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_144 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_514 ),
	.cout(Xd_0__inst_mult_6_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_143 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[13]),
	.datac(!din_a[18]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_509 ),
	.cout(Xd_0__inst_mult_1_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_144 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_514 ),
	.cout(Xd_0__inst_mult_1_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_143 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[1]),
	.datac(!din_a[6]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_509 ),
	.cout(Xd_0__inst_mult_0_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_144 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_514 ),
	.cout(Xd_0__inst_mult_0_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_143 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[37]),
	.datac(!din_a[42]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_509 ),
	.cout(Xd_0__inst_mult_3_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_144 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_514 ),
	.cout(Xd_0__inst_mult_3_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_152 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[25]),
	.datac(!din_a[30]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_554 ),
	.cout(Xd_0__inst_mult_2_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_153 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_559 ),
	.cout(Xd_0__inst_mult_2_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_151 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[349]),
	.datac(!din_a[355]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_549 ),
	.cout(Xd_0__inst_mult_29_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_152 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_554 ),
	.cout(Xd_0__inst_mult_29_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_145 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[337]),
	.datac(!din_a[343]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_519 ),
	.cout(Xd_0__inst_mult_28_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_146 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_524 ),
	.cout(Xd_0__inst_mult_28_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_145 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[373]),
	.datac(!din_a[379]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_519 ),
	.cout(Xd_0__inst_mult_31_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_146 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_524 ),
	.cout(Xd_0__inst_mult_31_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_145 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[361]),
	.datac(!din_a[367]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_519 ),
	.cout(Xd_0__inst_mult_30_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_146 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_524 ),
	.cout(Xd_0__inst_mult_30_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_151 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[253]),
	.datac(!din_a[259]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_549 ),
	.cout(Xd_0__inst_mult_21_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_152 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_554 ),
	.cout(Xd_0__inst_mult_21_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_151 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[241]),
	.datac(!din_a[247]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_549 ),
	.cout(Xd_0__inst_mult_20_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_152 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_554 ),
	.cout(Xd_0__inst_mult_20_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_151 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[277]),
	.datac(!din_a[283]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_549 ),
	.cout(Xd_0__inst_mult_23_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_152 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_554 ),
	.cout(Xd_0__inst_mult_23_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_151 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[265]),
	.datac(!din_a[271]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_549 ),
	.cout(Xd_0__inst_mult_22_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_152 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_554 ),
	.cout(Xd_0__inst_mult_22_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_151 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[205]),
	.datac(!din_a[211]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_549 ),
	.cout(Xd_0__inst_mult_17_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_152 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_554 ),
	.cout(Xd_0__inst_mult_17_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_151 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[193]),
	.datac(!din_a[199]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_549 ),
	.cout(Xd_0__inst_mult_16_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_152 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_554 ),
	.cout(Xd_0__inst_mult_16_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_151 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[229]),
	.datac(!din_a[235]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_549 ),
	.cout(Xd_0__inst_mult_19_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_152 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_554 ),
	.cout(Xd_0__inst_mult_19_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_140 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[217]),
	.datac(!din_a[223]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_494 ),
	.cout(Xd_0__inst_mult_18_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_141 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_499 ),
	.cout(Xd_0__inst_mult_18_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_145 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[157]),
	.datac(!din_a[163]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_519 ),
	.cout(Xd_0__inst_mult_13_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_146 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_524 ),
	.cout(Xd_0__inst_mult_13_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_140 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[145]),
	.datac(!din_a[151]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_494 ),
	.cout(Xd_0__inst_mult_12_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_141 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_499 ),
	.cout(Xd_0__inst_mult_12_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_140 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[181]),
	.datac(!din_a[187]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_494 ),
	.cout(Xd_0__inst_mult_15_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_141 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_499 ),
	.cout(Xd_0__inst_mult_15_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_140 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[169]),
	.datac(!din_a[175]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_485 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_494 ),
	.cout(Xd_0__inst_mult_14_495 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_141 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_689 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_499 ),
	.cout(Xd_0__inst_mult_14_500 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_145 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[109]),
	.datac(!din_a[115]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_519 ),
	.cout(Xd_0__inst_mult_9_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_146 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_524 ),
	.cout(Xd_0__inst_mult_9_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_145 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[97]),
	.datac(!din_a[103]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_519 ),
	.cout(Xd_0__inst_mult_8_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_146 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_524 ),
	.cout(Xd_0__inst_mult_8_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_145 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[133]),
	.datac(!din_a[139]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_519 ),
	.cout(Xd_0__inst_mult_11_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_146 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_524 ),
	.cout(Xd_0__inst_mult_11_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_145 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[121]),
	.datac(!din_a[127]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_519 ),
	.cout(Xd_0__inst_mult_10_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_146 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_524 ),
	.cout(Xd_0__inst_mult_10_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_145 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[61]),
	.datac(!din_a[67]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_519 ),
	.cout(Xd_0__inst_mult_5_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_146 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_524 ),
	.cout(Xd_0__inst_mult_5_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_145 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[49]),
	.datac(!din_a[55]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_519 ),
	.cout(Xd_0__inst_mult_4_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_146 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_524 ),
	.cout(Xd_0__inst_mult_4_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_145 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[85]),
	.datac(!din_a[91]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_519 ),
	.cout(Xd_0__inst_mult_7_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_146 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_524 ),
	.cout(Xd_0__inst_mult_7_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_145 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[73]),
	.datac(!din_a[79]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_519 ),
	.cout(Xd_0__inst_mult_6_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_146 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_524 ),
	.cout(Xd_0__inst_mult_6_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_145 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[13]),
	.datac(!din_a[19]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_519 ),
	.cout(Xd_0__inst_mult_1_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_146 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_524 ),
	.cout(Xd_0__inst_mult_1_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_145 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[1]),
	.datac(!din_a[7]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_519 ),
	.cout(Xd_0__inst_mult_0_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_146 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_524 ),
	.cout(Xd_0__inst_mult_0_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_145 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[37]),
	.datac(!din_a[43]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_519 ),
	.cout(Xd_0__inst_mult_3_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_146 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_524 ),
	.cout(Xd_0__inst_mult_3_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_154 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[25]),
	.datac(!din_a[31]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_564 ),
	.cout(Xd_0__inst_mult_2_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_155 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_569 ),
	.cout(Xd_0__inst_mult_2_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_153 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[349]),
	.datac(!din_a[356]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_559 ),
	.cout(Xd_0__inst_mult_29_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_154 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_564 ),
	.cout(Xd_0__inst_mult_29_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_155 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_569 ),
	.cout(Xd_0__inst_mult_29_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_29_156 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[356]),
	.datac(!din_a[349]),
	.datad(!din_b[357]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_574 ),
	.cout(Xd_0__inst_mult_29_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_147 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[337]),
	.datac(!din_a[344]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_529 ),
	.cout(Xd_0__inst_mult_28_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_148 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_534 ),
	.cout(Xd_0__inst_mult_28_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_149 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_539 ),
	.cout(Xd_0__inst_mult_28_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_28_150 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[344]),
	.datac(!din_a[337]),
	.datad(!din_b[345]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_544 ),
	.cout(Xd_0__inst_mult_28_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_147 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[373]),
	.datac(!din_a[380]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_529 ),
	.cout(Xd_0__inst_mult_31_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_148 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_534 ),
	.cout(Xd_0__inst_mult_31_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_149 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_539 ),
	.cout(Xd_0__inst_mult_31_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_31_150 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[380]),
	.datac(!din_a[373]),
	.datad(!din_b[381]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_544 ),
	.cout(Xd_0__inst_mult_31_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_147 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[361]),
	.datac(!din_a[368]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_529 ),
	.cout(Xd_0__inst_mult_30_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_148 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_534 ),
	.cout(Xd_0__inst_mult_30_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_149 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_539 ),
	.cout(Xd_0__inst_mult_30_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_30_150 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[368]),
	.datac(!din_a[361]),
	.datad(!din_b[369]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_544 ),
	.cout(Xd_0__inst_mult_30_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_160 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_594 ),
	.cout(Xd_0__inst_mult_25_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_25_161 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[308]),
	.datac(!din_a[301]),
	.datad(!din_b[309]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_599 ),
	.cout(Xd_0__inst_mult_25_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_191 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_749 ),
	.cout(Xd_0__inst_mult_24_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_24_192 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[296]),
	.datac(!din_a[289]),
	.datad(!din_b[297]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_754 ),
	.cout(Xd_0__inst_mult_24_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_160 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_594 ),
	.cout(Xd_0__inst_mult_27_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_27_161 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[332]),
	.datac(!din_a[325]),
	.datad(!din_b[333]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_599 ),
	.cout(Xd_0__inst_mult_27_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_191 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_749 ),
	.cout(Xd_0__inst_mult_26_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_26_192 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[320]),
	.datac(!din_a[313]),
	.datad(!din_b[321]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_754 ),
	.cout(Xd_0__inst_mult_26_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_153 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[253]),
	.datac(!din_a[260]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_559 ),
	.cout(Xd_0__inst_mult_21_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_154 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_564 ),
	.cout(Xd_0__inst_mult_21_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_155 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_569 ),
	.cout(Xd_0__inst_mult_21_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_21_156 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[260]),
	.datac(!din_a[253]),
	.datad(!din_b[261]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_574 ),
	.cout(Xd_0__inst_mult_21_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_153 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[241]),
	.datac(!din_a[248]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_559 ),
	.cout(Xd_0__inst_mult_20_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_154 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_564 ),
	.cout(Xd_0__inst_mult_20_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_155 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_569 ),
	.cout(Xd_0__inst_mult_20_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_20_156 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[248]),
	.datac(!din_a[241]),
	.datad(!din_b[249]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_574 ),
	.cout(Xd_0__inst_mult_20_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_153 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[277]),
	.datac(!din_a[284]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_559 ),
	.cout(Xd_0__inst_mult_23_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_154 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_564 ),
	.cout(Xd_0__inst_mult_23_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_155 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_569 ),
	.cout(Xd_0__inst_mult_23_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_23_156 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[284]),
	.datac(!din_a[277]),
	.datad(!din_b[285]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_574 ),
	.cout(Xd_0__inst_mult_23_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_153 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[265]),
	.datac(!din_a[272]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_559 ),
	.cout(Xd_0__inst_mult_22_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_154 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_564 ),
	.cout(Xd_0__inst_mult_22_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_155 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_569 ),
	.cout(Xd_0__inst_mult_22_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_22_156 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[272]),
	.datac(!din_a[265]),
	.datad(!din_b[273]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_574 ),
	.cout(Xd_0__inst_mult_22_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_153 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[205]),
	.datac(!din_a[212]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_559 ),
	.cout(Xd_0__inst_mult_17_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_154 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_564 ),
	.cout(Xd_0__inst_mult_17_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_155 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_569 ),
	.cout(Xd_0__inst_mult_17_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_17_156 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[212]),
	.datac(!din_a[205]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_574 ),
	.cout(Xd_0__inst_mult_17_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_153 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[193]),
	.datac(!din_a[200]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_559 ),
	.cout(Xd_0__inst_mult_16_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_154 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_564 ),
	.cout(Xd_0__inst_mult_16_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_155 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_569 ),
	.cout(Xd_0__inst_mult_16_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_16_156 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[200]),
	.datac(!din_a[193]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_574 ),
	.cout(Xd_0__inst_mult_16_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_153 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[229]),
	.datac(!din_a[236]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_559 ),
	.cout(Xd_0__inst_mult_19_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_154 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_564 ),
	.cout(Xd_0__inst_mult_19_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_155 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_569 ),
	.cout(Xd_0__inst_mult_19_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_19_156 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[236]),
	.datac(!din_a[229]),
	.datad(!din_b[237]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_574 ),
	.cout(Xd_0__inst_mult_19_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_142 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[217]),
	.datac(!din_a[224]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_504 ),
	.cout(Xd_0__inst_mult_18_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_143 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_509 ),
	.cout(Xd_0__inst_mult_18_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_144 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_514 ),
	.cout(Xd_0__inst_mult_18_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_18_145 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[224]),
	.datac(!din_a[217]),
	.datad(!din_b[225]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_519 ),
	.cout(Xd_0__inst_mult_18_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_147 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[157]),
	.datac(!din_a[164]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_529 ),
	.cout(Xd_0__inst_mult_13_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_148 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_534 ),
	.cout(Xd_0__inst_mult_13_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_149 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_539 ),
	.cout(Xd_0__inst_mult_13_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_13_150 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[164]),
	.datac(!din_a[157]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_544 ),
	.cout(Xd_0__inst_mult_13_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_142 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[145]),
	.datac(!din_a[152]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_504 ),
	.cout(Xd_0__inst_mult_12_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_143 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_509 ),
	.cout(Xd_0__inst_mult_12_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_144 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_514 ),
	.cout(Xd_0__inst_mult_12_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_12_145 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[152]),
	.datac(!din_a[145]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_519 ),
	.cout(Xd_0__inst_mult_12_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_142 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[181]),
	.datac(!din_a[188]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_504 ),
	.cout(Xd_0__inst_mult_15_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_143 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_509 ),
	.cout(Xd_0__inst_mult_15_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_144 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_514 ),
	.cout(Xd_0__inst_mult_15_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_15_145 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[188]),
	.datac(!din_a[181]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_519 ),
	.cout(Xd_0__inst_mult_15_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_80 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[369]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_80_sumout ),
	.cout(Xd_0__inst_mult_30_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_142 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[169]),
	.datac(!din_a[176]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_495 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_504 ),
	.cout(Xd_0__inst_mult_14_505 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_143 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_694 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_500 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_509 ),
	.cout(Xd_0__inst_mult_14_510 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_144 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_699 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_514 ),
	.cout(Xd_0__inst_mult_14_515 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_14_145 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[176]),
	.datac(!din_a[169]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_519 ),
	.cout(Xd_0__inst_mult_14_520 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_80 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[285]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_71 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_80_sumout ),
	.cout(Xd_0__inst_mult_23_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_147 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[109]),
	.datac(!din_a[116]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_529 ),
	.cout(Xd_0__inst_mult_9_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_148 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_534 ),
	.cout(Xd_0__inst_mult_9_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_149 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_539 ),
	.cout(Xd_0__inst_mult_9_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_9_150 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[116]),
	.datac(!din_a[109]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_544 ),
	.cout(Xd_0__inst_mult_9_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_80 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[153]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_80_sumout ),
	.cout(Xd_0__inst_mult_12_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_147 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[97]),
	.datac(!din_a[104]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_529 ),
	.cout(Xd_0__inst_mult_8_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_148 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_534 ),
	.cout(Xd_0__inst_mult_8_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_149 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_539 ),
	.cout(Xd_0__inst_mult_8_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_8_150 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[104]),
	.datac(!din_a[97]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_544 ),
	.cout(Xd_0__inst_mult_8_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_147 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[133]),
	.datac(!din_a[140]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_529 ),
	.cout(Xd_0__inst_mult_11_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_148 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_534 ),
	.cout(Xd_0__inst_mult_11_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_149 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_539 ),
	.cout(Xd_0__inst_mult_11_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_11_150 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[140]),
	.datac(!din_a[133]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_544 ),
	.cout(Xd_0__inst_mult_11_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_147 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[121]),
	.datac(!din_a[128]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_529 ),
	.cout(Xd_0__inst_mult_10_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_148 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_534 ),
	.cout(Xd_0__inst_mult_10_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_149 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_539 ),
	.cout(Xd_0__inst_mult_10_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_10_150 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[128]),
	.datac(!din_a[121]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_544 ),
	.cout(Xd_0__inst_mult_10_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_147 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[61]),
	.datac(!din_a[68]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_529 ),
	.cout(Xd_0__inst_mult_5_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_148 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_534 ),
	.cout(Xd_0__inst_mult_5_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_149 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_539 ),
	.cout(Xd_0__inst_mult_5_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_5_150 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[68]),
	.datac(!din_a[61]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_544 ),
	.cout(Xd_0__inst_mult_5_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_147 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[49]),
	.datac(!din_a[56]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_529 ),
	.cout(Xd_0__inst_mult_4_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_148 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_534 ),
	.cout(Xd_0__inst_mult_4_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_149 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_539 ),
	.cout(Xd_0__inst_mult_4_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_4_150 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[56]),
	.datac(!din_a[49]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_544 ),
	.cout(Xd_0__inst_mult_4_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_147 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[85]),
	.datac(!din_a[92]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_529 ),
	.cout(Xd_0__inst_mult_7_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_148 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_534 ),
	.cout(Xd_0__inst_mult_7_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_149 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_539 ),
	.cout(Xd_0__inst_mult_7_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_7_150 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[92]),
	.datac(!din_a[85]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_544 ),
	.cout(Xd_0__inst_mult_7_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_147 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[73]),
	.datac(!din_a[80]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_529 ),
	.cout(Xd_0__inst_mult_6_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_148 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_534 ),
	.cout(Xd_0__inst_mult_6_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_149 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_539 ),
	.cout(Xd_0__inst_mult_6_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_6_150 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[80]),
	.datac(!din_a[73]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_544 ),
	.cout(Xd_0__inst_mult_6_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_147 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[13]),
	.datac(!din_a[20]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_529 ),
	.cout(Xd_0__inst_mult_1_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_148 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_534 ),
	.cout(Xd_0__inst_mult_1_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_149 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_539 ),
	.cout(Xd_0__inst_mult_1_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_1_150 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[20]),
	.datac(!din_a[13]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_544 ),
	.cout(Xd_0__inst_mult_1_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_147 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[1]),
	.datac(!din_a[8]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_529 ),
	.cout(Xd_0__inst_mult_0_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_148 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_534 ),
	.cout(Xd_0__inst_mult_0_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_149 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_539 ),
	.cout(Xd_0__inst_mult_0_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_0_150 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[8]),
	.datac(!din_a[1]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_544 ),
	.cout(Xd_0__inst_mult_0_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_147 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[37]),
	.datac(!din_a[44]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_529 ),
	.cout(Xd_0__inst_mult_3_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_148 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_704 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_534 ),
	.cout(Xd_0__inst_mult_3_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_149 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_539 ),
	.cout(Xd_0__inst_mult_3_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_3_150 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[44]),
	.datac(!din_a[37]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_544 ),
	.cout(Xd_0__inst_mult_3_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_156 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[25]),
	.datac(!din_a[32]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_574 ),
	.cout(Xd_0__inst_mult_2_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_157 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_579 ),
	.cout(Xd_0__inst_mult_2_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_158 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_244 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_584 ),
	.cout(Xd_0__inst_mult_2_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000E1111),
	.shared_arith("off")
) Xd_0__inst_mult_2_159 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[32]),
	.datac(!din_a[25]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_589 ),
	.cout(Xd_0__inst_mult_2_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_157 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[349]),
	.datac(!din_a[357]),
	.datad(!din_b[348]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_579 ),
	.cout(Xd_0__inst_mult_29_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_158 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[350]),
	.datac(!Xd_0__inst_mult_29_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_584 ),
	.cout(Xd_0__inst_mult_29_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_159 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_589 ),
	.cout(Xd_0__inst_mult_29_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_160 (
// Equation(s):

	.dataa(!din_a[349]),
	.datab(!din_b[356]),
	.datac(!din_a[348]),
	.datad(!din_b[357]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_594 ),
	.cout(Xd_0__inst_mult_29_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_151 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[337]),
	.datac(!din_a[345]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_549 ),
	.cout(Xd_0__inst_mult_28_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_152 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_554 ),
	.cout(Xd_0__inst_mult_28_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_153 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_559 ),
	.cout(Xd_0__inst_mult_28_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_154 (
// Equation(s):

	.dataa(!din_a[337]),
	.datab(!din_b[344]),
	.datac(!din_a[336]),
	.datad(!din_b[345]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_564 ),
	.cout(Xd_0__inst_mult_28_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_151 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[373]),
	.datac(!din_a[381]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_549 ),
	.cout(Xd_0__inst_mult_31_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_152 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_554 ),
	.cout(Xd_0__inst_mult_31_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_153 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_559 ),
	.cout(Xd_0__inst_mult_31_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_154 (
// Equation(s):

	.dataa(!din_a[373]),
	.datab(!din_b[380]),
	.datac(!din_a[372]),
	.datad(!din_b[381]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_564 ),
	.cout(Xd_0__inst_mult_31_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_151 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[361]),
	.datac(!din_a[369]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_549 ),
	.cout(Xd_0__inst_mult_30_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_152 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_554 ),
	.cout(Xd_0__inst_mult_30_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_153 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_559 ),
	.cout(Xd_0__inst_mult_30_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_154 (
// Equation(s):

	.dataa(!din_a[361]),
	.datab(!din_b[368]),
	.datac(!din_a[360]),
	.datad(!din_b[369]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_564 ),
	.cout(Xd_0__inst_mult_30_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_162 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_604 ),
	.cout(Xd_0__inst_mult_25_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_163 (
// Equation(s):

	.dataa(!din_a[301]),
	.datab(!din_b[308]),
	.datac(!din_a[300]),
	.datad(!din_b[309]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_609 ),
	.cout(Xd_0__inst_mult_25_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_24_193 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[293]),
	.datac(!Xd_0__inst_mult_24_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_759 ),
	.cout(Xd_0__inst_mult_24_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_194 (
// Equation(s):

	.dataa(!din_a[289]),
	.datab(!din_b[296]),
	.datac(!din_a[288]),
	.datad(!din_b[297]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_764 ),
	.cout(Xd_0__inst_mult_24_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_162 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_604 ),
	.cout(Xd_0__inst_mult_27_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_163 (
// Equation(s):

	.dataa(!din_a[325]),
	.datab(!din_b[332]),
	.datac(!din_a[324]),
	.datad(!din_b[333]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_609 ),
	.cout(Xd_0__inst_mult_27_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_26_193 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[317]),
	.datac(!Xd_0__inst_mult_26_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_759 ),
	.cout(Xd_0__inst_mult_26_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_194 (
// Equation(s):

	.dataa(!din_a[313]),
	.datab(!din_b[320]),
	.datac(!din_a[312]),
	.datad(!din_b[321]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_764 ),
	.cout(Xd_0__inst_mult_26_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_157 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[253]),
	.datac(!din_a[261]),
	.datad(!din_b[252]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_579 ),
	.cout(Xd_0__inst_mult_21_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_158 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[254]),
	.datac(!Xd_0__inst_mult_21_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_584 ),
	.cout(Xd_0__inst_mult_21_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_159 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_589 ),
	.cout(Xd_0__inst_mult_21_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_160 (
// Equation(s):

	.dataa(!din_a[253]),
	.datab(!din_b[260]),
	.datac(!din_a[252]),
	.datad(!din_b[261]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_594 ),
	.cout(Xd_0__inst_mult_21_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_157 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[241]),
	.datac(!din_a[249]),
	.datad(!din_b[240]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_579 ),
	.cout(Xd_0__inst_mult_20_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_158 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[242]),
	.datac(!Xd_0__inst_mult_20_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_584 ),
	.cout(Xd_0__inst_mult_20_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_159 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_589 ),
	.cout(Xd_0__inst_mult_20_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_160 (
// Equation(s):

	.dataa(!din_a[241]),
	.datab(!din_b[248]),
	.datac(!din_a[240]),
	.datad(!din_b[249]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_594 ),
	.cout(Xd_0__inst_mult_20_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_157 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[277]),
	.datac(!din_a[285]),
	.datad(!din_b[276]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_579 ),
	.cout(Xd_0__inst_mult_23_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_158 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[278]),
	.datac(!Xd_0__inst_mult_23_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_584 ),
	.cout(Xd_0__inst_mult_23_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_159 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_589 ),
	.cout(Xd_0__inst_mult_23_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_160 (
// Equation(s):

	.dataa(!din_a[277]),
	.datab(!din_b[284]),
	.datac(!din_a[276]),
	.datad(!din_b[285]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_594 ),
	.cout(Xd_0__inst_mult_23_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_157 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[265]),
	.datac(!din_a[273]),
	.datad(!din_b[264]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_579 ),
	.cout(Xd_0__inst_mult_22_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_158 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[266]),
	.datac(!Xd_0__inst_mult_22_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_584 ),
	.cout(Xd_0__inst_mult_22_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_159 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_589 ),
	.cout(Xd_0__inst_mult_22_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_160 (
// Equation(s):

	.dataa(!din_a[265]),
	.datab(!din_b[272]),
	.datac(!din_a[264]),
	.datad(!din_b[273]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_594 ),
	.cout(Xd_0__inst_mult_22_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_157 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[205]),
	.datac(!din_a[213]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_579 ),
	.cout(Xd_0__inst_mult_17_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_158 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[206]),
	.datac(!Xd_0__inst_mult_17_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_584 ),
	.cout(Xd_0__inst_mult_17_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_159 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_589 ),
	.cout(Xd_0__inst_mult_17_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_160 (
// Equation(s):

	.dataa(!din_a[205]),
	.datab(!din_b[212]),
	.datac(!din_a[204]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_594 ),
	.cout(Xd_0__inst_mult_17_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_157 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[193]),
	.datac(!din_a[201]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_579 ),
	.cout(Xd_0__inst_mult_16_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_158 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[194]),
	.datac(!Xd_0__inst_mult_16_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_584 ),
	.cout(Xd_0__inst_mult_16_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_159 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_589 ),
	.cout(Xd_0__inst_mult_16_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_160 (
// Equation(s):

	.dataa(!din_a[193]),
	.datab(!din_b[200]),
	.datac(!din_a[192]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_594 ),
	.cout(Xd_0__inst_mult_16_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_157 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[229]),
	.datac(!din_a[237]),
	.datad(!din_b[228]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_579 ),
	.cout(Xd_0__inst_mult_19_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_158 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[230]),
	.datac(!Xd_0__inst_mult_19_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_584 ),
	.cout(Xd_0__inst_mult_19_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_159 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_589 ),
	.cout(Xd_0__inst_mult_19_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_160 (
// Equation(s):

	.dataa(!din_a[229]),
	.datab(!din_b[236]),
	.datac(!din_a[228]),
	.datad(!din_b[237]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_594 ),
	.cout(Xd_0__inst_mult_19_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_146 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[217]),
	.datac(!din_a[225]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_524 ),
	.cout(Xd_0__inst_mult_18_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_147 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_529 ),
	.cout(Xd_0__inst_mult_18_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_148 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_534 ),
	.cout(Xd_0__inst_mult_18_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_149 (
// Equation(s):

	.dataa(!din_a[217]),
	.datab(!din_b[224]),
	.datac(!din_a[216]),
	.datad(!din_b[225]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_539 ),
	.cout(Xd_0__inst_mult_18_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_151 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[157]),
	.datac(!din_a[165]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_549 ),
	.cout(Xd_0__inst_mult_13_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_152 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_554 ),
	.cout(Xd_0__inst_mult_13_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_153 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_559 ),
	.cout(Xd_0__inst_mult_13_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_154 (
// Equation(s):

	.dataa(!din_a[157]),
	.datab(!din_b[164]),
	.datac(!din_a[156]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_564 ),
	.cout(Xd_0__inst_mult_13_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_146 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[145]),
	.datac(!din_a[153]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_524 ),
	.cout(Xd_0__inst_mult_12_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_147 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_529 ),
	.cout(Xd_0__inst_mult_12_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_148 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_534 ),
	.cout(Xd_0__inst_mult_12_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_149 (
// Equation(s):

	.dataa(!din_a[145]),
	.datab(!din_b[152]),
	.datac(!din_a[144]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_539 ),
	.cout(Xd_0__inst_mult_12_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_146 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[181]),
	.datac(!din_a[189]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_524 ),
	.cout(Xd_0__inst_mult_15_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_147 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_529 ),
	.cout(Xd_0__inst_mult_15_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_148 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_534 ),
	.cout(Xd_0__inst_mult_15_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_149 (
// Equation(s):

	.dataa(!din_a[181]),
	.datab(!din_b[188]),
	.datac(!din_a[180]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_539 ),
	.cout(Xd_0__inst_mult_15_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_146 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[169]),
	.datac(!din_a[177]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_505 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_524 ),
	.cout(Xd_0__inst_mult_14_525 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_147 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_709 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_510 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_529 ),
	.cout(Xd_0__inst_mult_14_530 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_148 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_714 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_515 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_534 ),
	.cout(Xd_0__inst_mult_14_535 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_149 (
// Equation(s):

	.dataa(!din_a[169]),
	.datab(!din_b[176]),
	.datac(!din_a[168]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_539 ),
	.cout(Xd_0__inst_mult_14_540 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_151 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[109]),
	.datac(!din_a[117]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_549 ),
	.cout(Xd_0__inst_mult_9_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_152 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_554 ),
	.cout(Xd_0__inst_mult_9_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_153 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_559 ),
	.cout(Xd_0__inst_mult_9_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_154 (
// Equation(s):

	.dataa(!din_a[109]),
	.datab(!din_b[116]),
	.datac(!din_a[108]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_564 ),
	.cout(Xd_0__inst_mult_9_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_151 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[97]),
	.datac(!din_a[105]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_549 ),
	.cout(Xd_0__inst_mult_8_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_152 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_554 ),
	.cout(Xd_0__inst_mult_8_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_153 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_559 ),
	.cout(Xd_0__inst_mult_8_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_154 (
// Equation(s):

	.dataa(!din_a[97]),
	.datab(!din_b[104]),
	.datac(!din_a[96]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_564 ),
	.cout(Xd_0__inst_mult_8_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_151 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[133]),
	.datac(!din_a[141]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_549 ),
	.cout(Xd_0__inst_mult_11_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_152 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_554 ),
	.cout(Xd_0__inst_mult_11_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_153 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_559 ),
	.cout(Xd_0__inst_mult_11_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_154 (
// Equation(s):

	.dataa(!din_a[133]),
	.datab(!din_b[140]),
	.datac(!din_a[132]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_564 ),
	.cout(Xd_0__inst_mult_11_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_151 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[121]),
	.datac(!din_a[129]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_549 ),
	.cout(Xd_0__inst_mult_10_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_152 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_554 ),
	.cout(Xd_0__inst_mult_10_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_153 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_559 ),
	.cout(Xd_0__inst_mult_10_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_154 (
// Equation(s):

	.dataa(!din_a[121]),
	.datab(!din_b[128]),
	.datac(!din_a[120]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_564 ),
	.cout(Xd_0__inst_mult_10_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_151 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[61]),
	.datac(!din_a[69]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_549 ),
	.cout(Xd_0__inst_mult_5_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_152 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_554 ),
	.cout(Xd_0__inst_mult_5_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_153 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_559 ),
	.cout(Xd_0__inst_mult_5_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_154 (
// Equation(s):

	.dataa(!din_a[61]),
	.datab(!din_b[68]),
	.datac(!din_a[60]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_564 ),
	.cout(Xd_0__inst_mult_5_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_151 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[49]),
	.datac(!din_a[57]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_549 ),
	.cout(Xd_0__inst_mult_4_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_152 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_554 ),
	.cout(Xd_0__inst_mult_4_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_153 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_559 ),
	.cout(Xd_0__inst_mult_4_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_154 (
// Equation(s):

	.dataa(!din_a[49]),
	.datab(!din_b[56]),
	.datac(!din_a[48]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_564 ),
	.cout(Xd_0__inst_mult_4_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_151 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[85]),
	.datac(!din_a[93]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_549 ),
	.cout(Xd_0__inst_mult_7_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_152 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_554 ),
	.cout(Xd_0__inst_mult_7_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_153 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_559 ),
	.cout(Xd_0__inst_mult_7_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_154 (
// Equation(s):

	.dataa(!din_a[85]),
	.datab(!din_b[92]),
	.datac(!din_a[84]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_564 ),
	.cout(Xd_0__inst_mult_7_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_151 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[73]),
	.datac(!din_a[81]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_549 ),
	.cout(Xd_0__inst_mult_6_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_152 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_554 ),
	.cout(Xd_0__inst_mult_6_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_153 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_559 ),
	.cout(Xd_0__inst_mult_6_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_154 (
// Equation(s):

	.dataa(!din_a[73]),
	.datab(!din_b[80]),
	.datac(!din_a[72]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_564 ),
	.cout(Xd_0__inst_mult_6_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_151 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[13]),
	.datac(!din_a[21]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_549 ),
	.cout(Xd_0__inst_mult_1_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_152 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_554 ),
	.cout(Xd_0__inst_mult_1_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_153 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_559 ),
	.cout(Xd_0__inst_mult_1_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_154 (
// Equation(s):

	.dataa(!din_a[13]),
	.datab(!din_b[20]),
	.datac(!din_a[12]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_564 ),
	.cout(Xd_0__inst_mult_1_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_151 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[1]),
	.datac(!din_a[9]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_549 ),
	.cout(Xd_0__inst_mult_0_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_152 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_554 ),
	.cout(Xd_0__inst_mult_0_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_153 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_559 ),
	.cout(Xd_0__inst_mult_0_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_154 (
// Equation(s):

	.dataa(!din_a[1]),
	.datab(!din_b[8]),
	.datac(!din_a[0]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_564 ),
	.cout(Xd_0__inst_mult_0_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_151 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[37]),
	.datac(!din_a[45]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_549 ),
	.cout(Xd_0__inst_mult_3_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_152 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_554 ),
	.cout(Xd_0__inst_mult_3_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_153 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_540 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_559 ),
	.cout(Xd_0__inst_mult_3_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_154 (
// Equation(s):

	.dataa(!din_a[37]),
	.datab(!din_b[44]),
	.datac(!din_a[36]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_564 ),
	.cout(Xd_0__inst_mult_3_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_160 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[25]),
	.datac(!din_a[33]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_594 ),
	.cout(Xd_0__inst_mult_2_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_161 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_599 ),
	.cout(Xd_0__inst_mult_2_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_162 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_239 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_604 ),
	.cout(Xd_0__inst_mult_2_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000000111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_163 (
// Equation(s):

	.dataa(!din_a[25]),
	.datab(!din_b[32]),
	.datac(!din_a[24]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_609 ),
	.cout(Xd_0__inst_mult_2_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_161 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_599 ),
	.cout(Xd_0__inst_mult_29_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_162 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[356]),
	.datac(!din_a[348]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_604 ),
	.cout(Xd_0__inst_mult_29_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_155 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[337]),
	.datac(!din_a[346]),
	.datad(!din_b[336]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_569 ),
	.cout(Xd_0__inst_mult_28_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_156 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_574 ),
	.cout(Xd_0__inst_mult_28_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_157 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_579 ),
	.cout(Xd_0__inst_mult_28_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_158 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[344]),
	.datac(!din_a[336]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_584 ),
	.cout(Xd_0__inst_mult_28_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_155 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[373]),
	.datac(!din_a[382]),
	.datad(!din_b[372]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_569 ),
	.cout(Xd_0__inst_mult_31_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_156 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_574 ),
	.cout(Xd_0__inst_mult_31_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_157 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_579 ),
	.cout(Xd_0__inst_mult_31_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_158 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[380]),
	.datac(!din_a[372]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_584 ),
	.cout(Xd_0__inst_mult_31_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_155 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[361]),
	.datac(!din_a[370]),
	.datad(!din_b[360]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_569 ),
	.cout(Xd_0__inst_mult_30_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_156 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_574 ),
	.cout(Xd_0__inst_mult_30_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_157 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_579 ),
	.cout(Xd_0__inst_mult_30_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_158 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[368]),
	.datac(!din_a[360]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_584 ),
	.cout(Xd_0__inst_mult_30_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_164 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_614 ),
	.cout(Xd_0__inst_mult_25_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_165 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[308]),
	.datac(!din_a[300]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_619 ),
	.cout(Xd_0__inst_mult_25_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_195 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[296]),
	.datac(!din_a[288]),
	.datad(!din_b[298]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_769 ),
	.cout(Xd_0__inst_mult_24_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_164 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_614 ),
	.cout(Xd_0__inst_mult_27_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_165 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[332]),
	.datac(!din_a[324]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_619 ),
	.cout(Xd_0__inst_mult_27_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_195 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[320]),
	.datac(!din_a[312]),
	.datad(!din_b[322]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_769 ),
	.cout(Xd_0__inst_mult_26_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_161 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_599 ),
	.cout(Xd_0__inst_mult_21_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_162 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[260]),
	.datac(!din_a[252]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_604 ),
	.cout(Xd_0__inst_mult_21_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_161 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_599 ),
	.cout(Xd_0__inst_mult_20_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_162 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[248]),
	.datac(!din_a[240]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_604 ),
	.cout(Xd_0__inst_mult_20_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_161 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_599 ),
	.cout(Xd_0__inst_mult_23_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_162 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[284]),
	.datac(!din_a[276]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_604 ),
	.cout(Xd_0__inst_mult_23_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_161 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_599 ),
	.cout(Xd_0__inst_mult_22_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_162 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[272]),
	.datac(!din_a[264]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_604 ),
	.cout(Xd_0__inst_mult_22_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_161 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_599 ),
	.cout(Xd_0__inst_mult_17_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_162 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[212]),
	.datac(!din_a[204]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_604 ),
	.cout(Xd_0__inst_mult_17_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_161 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_599 ),
	.cout(Xd_0__inst_mult_16_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_162 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[200]),
	.datac(!din_a[192]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_604 ),
	.cout(Xd_0__inst_mult_16_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_161 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_599 ),
	.cout(Xd_0__inst_mult_19_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_162 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[236]),
	.datac(!din_a[228]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_604 ),
	.cout(Xd_0__inst_mult_19_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_150 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[217]),
	.datac(!din_a[226]),
	.datad(!din_b[216]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_544 ),
	.cout(Xd_0__inst_mult_18_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_151 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_549 ),
	.cout(Xd_0__inst_mult_18_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_152 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_554 ),
	.cout(Xd_0__inst_mult_18_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_153 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[224]),
	.datac(!din_a[216]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_559 ),
	.cout(Xd_0__inst_mult_18_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_155 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[157]),
	.datac(!din_a[166]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_569 ),
	.cout(Xd_0__inst_mult_13_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_156 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_574 ),
	.cout(Xd_0__inst_mult_13_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_157 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_579 ),
	.cout(Xd_0__inst_mult_13_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_158 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[164]),
	.datac(!din_a[156]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_584 ),
	.cout(Xd_0__inst_mult_13_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_150 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[145]),
	.datac(!din_a[154]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_544 ),
	.cout(Xd_0__inst_mult_12_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_151 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_549 ),
	.cout(Xd_0__inst_mult_12_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_152 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_554 ),
	.cout(Xd_0__inst_mult_12_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_153 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[152]),
	.datac(!din_a[144]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_559 ),
	.cout(Xd_0__inst_mult_12_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_150 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[181]),
	.datac(!din_a[190]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_544 ),
	.cout(Xd_0__inst_mult_15_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_151 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_549 ),
	.cout(Xd_0__inst_mult_15_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_152 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_554 ),
	.cout(Xd_0__inst_mult_15_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_153 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[188]),
	.datac(!din_a[180]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_559 ),
	.cout(Xd_0__inst_mult_15_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_150 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[169]),
	.datac(!din_a[178]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_525 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_544 ),
	.cout(Xd_0__inst_mult_14_545 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_151 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_719 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_530 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_549 ),
	.cout(Xd_0__inst_mult_14_550 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_152 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_724 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_535 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_554 ),
	.cout(Xd_0__inst_mult_14_555 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_153 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[176]),
	.datac(!din_a[168]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_520 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_559 ),
	.cout(Xd_0__inst_mult_14_560 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_155 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[109]),
	.datac(!din_a[118]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_569 ),
	.cout(Xd_0__inst_mult_9_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_156 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_574 ),
	.cout(Xd_0__inst_mult_9_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_157 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_579 ),
	.cout(Xd_0__inst_mult_9_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_158 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[116]),
	.datac(!din_a[108]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_584 ),
	.cout(Xd_0__inst_mult_9_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_155 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[97]),
	.datac(!din_a[106]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_569 ),
	.cout(Xd_0__inst_mult_8_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_156 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_574 ),
	.cout(Xd_0__inst_mult_8_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_157 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_579 ),
	.cout(Xd_0__inst_mult_8_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_158 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[104]),
	.datac(!din_a[96]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_584 ),
	.cout(Xd_0__inst_mult_8_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_155 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[133]),
	.datac(!din_a[142]),
	.datad(!din_b[132]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_569 ),
	.cout(Xd_0__inst_mult_11_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_156 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_574 ),
	.cout(Xd_0__inst_mult_11_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_157 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_579 ),
	.cout(Xd_0__inst_mult_11_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_158 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[140]),
	.datac(!din_a[132]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_584 ),
	.cout(Xd_0__inst_mult_11_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_155 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[121]),
	.datac(!din_a[130]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_569 ),
	.cout(Xd_0__inst_mult_10_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_156 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_574 ),
	.cout(Xd_0__inst_mult_10_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_157 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_579 ),
	.cout(Xd_0__inst_mult_10_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_158 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[128]),
	.datac(!din_a[120]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_584 ),
	.cout(Xd_0__inst_mult_10_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_155 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[61]),
	.datac(!din_a[70]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_569 ),
	.cout(Xd_0__inst_mult_5_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_156 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_574 ),
	.cout(Xd_0__inst_mult_5_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_157 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_579 ),
	.cout(Xd_0__inst_mult_5_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_158 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[68]),
	.datac(!din_a[60]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_584 ),
	.cout(Xd_0__inst_mult_5_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_155 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[49]),
	.datac(!din_a[58]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_569 ),
	.cout(Xd_0__inst_mult_4_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_156 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_574 ),
	.cout(Xd_0__inst_mult_4_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_157 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_579 ),
	.cout(Xd_0__inst_mult_4_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_158 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[56]),
	.datac(!din_a[48]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_584 ),
	.cout(Xd_0__inst_mult_4_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_155 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[85]),
	.datac(!din_a[94]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_569 ),
	.cout(Xd_0__inst_mult_7_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_156 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_574 ),
	.cout(Xd_0__inst_mult_7_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_157 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_579 ),
	.cout(Xd_0__inst_mult_7_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_158 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[92]),
	.datac(!din_a[84]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_584 ),
	.cout(Xd_0__inst_mult_7_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_155 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[73]),
	.datac(!din_a[82]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_569 ),
	.cout(Xd_0__inst_mult_6_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_156 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_574 ),
	.cout(Xd_0__inst_mult_6_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_157 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_579 ),
	.cout(Xd_0__inst_mult_6_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_158 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[80]),
	.datac(!din_a[72]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_584 ),
	.cout(Xd_0__inst_mult_6_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_155 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[13]),
	.datac(!din_a[22]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_569 ),
	.cout(Xd_0__inst_mult_1_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_156 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_574 ),
	.cout(Xd_0__inst_mult_1_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_157 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_579 ),
	.cout(Xd_0__inst_mult_1_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_158 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[20]),
	.datac(!din_a[12]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_584 ),
	.cout(Xd_0__inst_mult_1_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_155 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[1]),
	.datac(!din_a[10]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_569 ),
	.cout(Xd_0__inst_mult_0_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_156 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_574 ),
	.cout(Xd_0__inst_mult_0_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_157 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_579 ),
	.cout(Xd_0__inst_mult_0_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_158 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[8]),
	.datac(!din_a[0]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_584 ),
	.cout(Xd_0__inst_mult_0_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_155 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[37]),
	.datac(!din_a[46]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_569 ),
	.cout(Xd_0__inst_mult_3_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_156 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_574 ),
	.cout(Xd_0__inst_mult_3_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_157 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_579 ),
	.cout(Xd_0__inst_mult_3_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_158 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[44]),
	.datac(!din_a[36]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_584 ),
	.cout(Xd_0__inst_mult_3_585 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_164 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[25]),
	.datac(!din_a[34]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_614 ),
	.cout(Xd_0__inst_mult_2_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_165 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_619 ),
	.cout(Xd_0__inst_mult_2_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_166 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_234 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_624 ),
	.cout(Xd_0__inst_mult_2_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_167 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[32]),
	.datac(!din_a[24]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_629 ),
	.cout(Xd_0__inst_mult_2_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_163 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_609 ),
	.cout(Xd_0__inst_mult_29_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_164 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_614 ),
	.cout(Xd_0__inst_mult_29_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_159 (
// Equation(s):

	.dataa(!din_a[346]),
	.datab(!din_b[337]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_589 ),
	.cout(Xd_0__inst_mult_28_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_160 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[338]),
	.datac(!Xd_0__inst_mult_28_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_594 ),
	.cout(Xd_0__inst_mult_28_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_161 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_599 ),
	.cout(Xd_0__inst_mult_28_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_162 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_604 ),
	.cout(Xd_0__inst_mult_28_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_159 (
// Equation(s):

	.dataa(!din_a[382]),
	.datab(!din_b[373]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_589 ),
	.cout(Xd_0__inst_mult_31_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_160 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[374]),
	.datac(!Xd_0__inst_mult_31_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_594 ),
	.cout(Xd_0__inst_mult_31_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_161 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_599 ),
	.cout(Xd_0__inst_mult_31_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_162 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_604 ),
	.cout(Xd_0__inst_mult_31_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_159 (
// Equation(s):

	.dataa(!din_a[370]),
	.datab(!din_b[361]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_589 ),
	.cout(Xd_0__inst_mult_30_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_160 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[362]),
	.datac(!Xd_0__inst_mult_30_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_594 ),
	.cout(Xd_0__inst_mult_30_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_161 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_599 ),
	.cout(Xd_0__inst_mult_30_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_162 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_604 ),
	.cout(Xd_0__inst_mult_30_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_166 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_624 ),
	.cout(Xd_0__inst_mult_25_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_167 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_629 ),
	.cout(Xd_0__inst_mult_25_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_166 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_624 ),
	.cout(Xd_0__inst_mult_27_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_167 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_629 ),
	.cout(Xd_0__inst_mult_27_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_163 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_609 ),
	.cout(Xd_0__inst_mult_21_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_164 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_614 ),
	.cout(Xd_0__inst_mult_21_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_163 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_609 ),
	.cout(Xd_0__inst_mult_20_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_164 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_614 ),
	.cout(Xd_0__inst_mult_20_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_163 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_609 ),
	.cout(Xd_0__inst_mult_23_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_164 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_614 ),
	.cout(Xd_0__inst_mult_23_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_163 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_609 ),
	.cout(Xd_0__inst_mult_22_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_164 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_614 ),
	.cout(Xd_0__inst_mult_22_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_163 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_609 ),
	.cout(Xd_0__inst_mult_17_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_164 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_614 ),
	.cout(Xd_0__inst_mult_17_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_163 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_609 ),
	.cout(Xd_0__inst_mult_16_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_164 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_614 ),
	.cout(Xd_0__inst_mult_16_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_163 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_609 ),
	.cout(Xd_0__inst_mult_19_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_164 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_614 ),
	.cout(Xd_0__inst_mult_19_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_154 (
// Equation(s):

	.dataa(!din_a[226]),
	.datab(!din_b[217]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_564 ),
	.cout(Xd_0__inst_mult_18_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_155 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[218]),
	.datac(!Xd_0__inst_mult_18_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_569 ),
	.cout(Xd_0__inst_mult_18_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_156 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_574 ),
	.cout(Xd_0__inst_mult_18_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_157 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_579 ),
	.cout(Xd_0__inst_mult_18_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_159 (
// Equation(s):

	.dataa(!din_a[166]),
	.datab(!din_b[157]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_589 ),
	.cout(Xd_0__inst_mult_13_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_160 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[158]),
	.datac(!Xd_0__inst_mult_13_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_594 ),
	.cout(Xd_0__inst_mult_13_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_161 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_599 ),
	.cout(Xd_0__inst_mult_13_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_162 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_604 ),
	.cout(Xd_0__inst_mult_13_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_154 (
// Equation(s):

	.dataa(!din_a[154]),
	.datab(!din_b[145]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_564 ),
	.cout(Xd_0__inst_mult_12_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_155 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[146]),
	.datac(!Xd_0__inst_mult_12_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_569 ),
	.cout(Xd_0__inst_mult_12_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_156 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_574 ),
	.cout(Xd_0__inst_mult_12_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_157 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_579 ),
	.cout(Xd_0__inst_mult_12_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_154 (
// Equation(s):

	.dataa(!din_a[190]),
	.datab(!din_b[181]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_564 ),
	.cout(Xd_0__inst_mult_15_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_155 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[182]),
	.datac(!Xd_0__inst_mult_15_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_569 ),
	.cout(Xd_0__inst_mult_15_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_156 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_574 ),
	.cout(Xd_0__inst_mult_15_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_157 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_579 ),
	.cout(Xd_0__inst_mult_15_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_154 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[169]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_545 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_564 ),
	.cout(Xd_0__inst_mult_14_565 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_155 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[170]),
	.datac(!Xd_0__inst_mult_14_729 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_550 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_569 ),
	.cout(Xd_0__inst_mult_14_570 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_156 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_734 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_555 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_574 ),
	.cout(Xd_0__inst_mult_14_575 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_157 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_579 ),
	.cout(Xd_0__inst_mult_14_580 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_159 (
// Equation(s):

	.dataa(!din_a[118]),
	.datab(!din_b[109]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_589 ),
	.cout(Xd_0__inst_mult_9_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_160 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[110]),
	.datac(!Xd_0__inst_mult_9_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_594 ),
	.cout(Xd_0__inst_mult_9_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_161 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_599 ),
	.cout(Xd_0__inst_mult_9_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_162 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_604 ),
	.cout(Xd_0__inst_mult_9_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_159 (
// Equation(s):

	.dataa(!din_a[106]),
	.datab(!din_b[97]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_589 ),
	.cout(Xd_0__inst_mult_8_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_160 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[98]),
	.datac(!Xd_0__inst_mult_8_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_594 ),
	.cout(Xd_0__inst_mult_8_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_161 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_599 ),
	.cout(Xd_0__inst_mult_8_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_162 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_604 ),
	.cout(Xd_0__inst_mult_8_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_159 (
// Equation(s):

	.dataa(!din_a[142]),
	.datab(!din_b[133]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_589 ),
	.cout(Xd_0__inst_mult_11_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_160 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[134]),
	.datac(!Xd_0__inst_mult_11_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_594 ),
	.cout(Xd_0__inst_mult_11_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_161 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_599 ),
	.cout(Xd_0__inst_mult_11_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_162 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_604 ),
	.cout(Xd_0__inst_mult_11_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_159 (
// Equation(s):

	.dataa(!din_a[130]),
	.datab(!din_b[121]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_589 ),
	.cout(Xd_0__inst_mult_10_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_160 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[122]),
	.datac(!Xd_0__inst_mult_10_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_594 ),
	.cout(Xd_0__inst_mult_10_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_161 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_599 ),
	.cout(Xd_0__inst_mult_10_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_162 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_604 ),
	.cout(Xd_0__inst_mult_10_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_159 (
// Equation(s):

	.dataa(!din_a[70]),
	.datab(!din_b[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_589 ),
	.cout(Xd_0__inst_mult_5_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_160 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[62]),
	.datac(!Xd_0__inst_mult_5_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_594 ),
	.cout(Xd_0__inst_mult_5_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_161 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_599 ),
	.cout(Xd_0__inst_mult_5_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_162 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_604 ),
	.cout(Xd_0__inst_mult_5_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_159 (
// Equation(s):

	.dataa(!din_a[58]),
	.datab(!din_b[49]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_589 ),
	.cout(Xd_0__inst_mult_4_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_160 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[50]),
	.datac(!Xd_0__inst_mult_4_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_594 ),
	.cout(Xd_0__inst_mult_4_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_161 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_599 ),
	.cout(Xd_0__inst_mult_4_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_162 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_604 ),
	.cout(Xd_0__inst_mult_4_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_159 (
// Equation(s):

	.dataa(!din_a[94]),
	.datab(!din_b[85]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_589 ),
	.cout(Xd_0__inst_mult_7_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_160 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[86]),
	.datac(!Xd_0__inst_mult_7_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_594 ),
	.cout(Xd_0__inst_mult_7_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_161 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_599 ),
	.cout(Xd_0__inst_mult_7_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_162 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_604 ),
	.cout(Xd_0__inst_mult_7_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_159 (
// Equation(s):

	.dataa(!din_a[82]),
	.datab(!din_b[73]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_589 ),
	.cout(Xd_0__inst_mult_6_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_160 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[74]),
	.datac(!Xd_0__inst_mult_6_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_594 ),
	.cout(Xd_0__inst_mult_6_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_161 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_599 ),
	.cout(Xd_0__inst_mult_6_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_162 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_604 ),
	.cout(Xd_0__inst_mult_6_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_159 (
// Equation(s):

	.dataa(!din_a[22]),
	.datab(!din_b[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_589 ),
	.cout(Xd_0__inst_mult_1_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_160 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[14]),
	.datac(!Xd_0__inst_mult_1_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_594 ),
	.cout(Xd_0__inst_mult_1_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_161 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_599 ),
	.cout(Xd_0__inst_mult_1_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_162 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_604 ),
	.cout(Xd_0__inst_mult_1_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_159 (
// Equation(s):

	.dataa(!din_a[10]),
	.datab(!din_b[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_589 ),
	.cout(Xd_0__inst_mult_0_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_160 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[2]),
	.datac(!Xd_0__inst_mult_0_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_594 ),
	.cout(Xd_0__inst_mult_0_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_161 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_599 ),
	.cout(Xd_0__inst_mult_0_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_162 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_604 ),
	.cout(Xd_0__inst_mult_0_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_159 (
// Equation(s):

	.dataa(!din_a[46]),
	.datab(!din_b[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_589 ),
	.cout(Xd_0__inst_mult_3_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_160 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[38]),
	.datac(!Xd_0__inst_mult_3_739 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_594 ),
	.cout(Xd_0__inst_mult_3_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_161 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_599 ),
	.cout(Xd_0__inst_mult_3_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_162 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_604 ),
	.cout(Xd_0__inst_mult_3_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_168 (
// Equation(s):

	.dataa(!din_a[34]),
	.datab(!din_b[25]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_634 ),
	.cout(Xd_0__inst_mult_2_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_169 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[26]),
	.datac(!Xd_0__inst_mult_2_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_639 ),
	.cout(Xd_0__inst_mult_2_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_170 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_229 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_644 ),
	.cout(Xd_0__inst_mult_2_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_171 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_649 ),
	.cout(Xd_0__inst_mult_2_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_165 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_619 ),
	.cout(Xd_0__inst_mult_29_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_166 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_624 ),
	.cout(Xd_0__inst_mult_29_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_163 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_609 ),
	.cout(Xd_0__inst_mult_28_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_164 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_614 ),
	.cout(Xd_0__inst_mult_28_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_163 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_609 ),
	.cout(Xd_0__inst_mult_31_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_164 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_614 ),
	.cout(Xd_0__inst_mult_31_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_163 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_609 ),
	.cout(Xd_0__inst_mult_30_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_164 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_614 ),
	.cout(Xd_0__inst_mult_30_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_168 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_634 ),
	.cout(Xd_0__inst_mult_25_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_169 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_639 ),
	.cout(Xd_0__inst_mult_25_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_168 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_634 ),
	.cout(Xd_0__inst_mult_27_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_169 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_639 ),
	.cout(Xd_0__inst_mult_27_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_165 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_619 ),
	.cout(Xd_0__inst_mult_21_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_166 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_624 ),
	.cout(Xd_0__inst_mult_21_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_165 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_619 ),
	.cout(Xd_0__inst_mult_20_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_166 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_624 ),
	.cout(Xd_0__inst_mult_20_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_165 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_619 ),
	.cout(Xd_0__inst_mult_23_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_166 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_624 ),
	.cout(Xd_0__inst_mult_23_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_165 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_619 ),
	.cout(Xd_0__inst_mult_22_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_166 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_624 ),
	.cout(Xd_0__inst_mult_22_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_165 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_619 ),
	.cout(Xd_0__inst_mult_17_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_166 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_624 ),
	.cout(Xd_0__inst_mult_17_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_165 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_619 ),
	.cout(Xd_0__inst_mult_16_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_166 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_624 ),
	.cout(Xd_0__inst_mult_16_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_165 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_619 ),
	.cout(Xd_0__inst_mult_19_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_166 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_624 ),
	.cout(Xd_0__inst_mult_19_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_158 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_584 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_159 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[219]),
	.datac(!Xd_0__inst_mult_18_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_589 ),
	.cout(Xd_0__inst_mult_18_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_160 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_594 ),
	.cout(Xd_0__inst_mult_18_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_161 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_599 ),
	.cout(Xd_0__inst_mult_18_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_163 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_609 ),
	.cout(Xd_0__inst_mult_13_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_164 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_614 ),
	.cout(Xd_0__inst_mult_13_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_158 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_584 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_159 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[147]),
	.datac(!Xd_0__inst_mult_12_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_589 ),
	.cout(Xd_0__inst_mult_12_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_160 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_594 ),
	.cout(Xd_0__inst_mult_12_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_161 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_599 ),
	.cout(Xd_0__inst_mult_12_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_158 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_584 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_159 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[183]),
	.datac(!Xd_0__inst_mult_15_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_589 ),
	.cout(Xd_0__inst_mult_15_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_160 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_594 ),
	.cout(Xd_0__inst_mult_15_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_161 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_599 ),
	.cout(Xd_0__inst_mult_15_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_158 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_565 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_584 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_159 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[171]),
	.datac(!Xd_0__inst_mult_14_749 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_570 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_589 ),
	.cout(Xd_0__inst_mult_14_590 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_160 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_575 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_594 ),
	.cout(Xd_0__inst_mult_14_595 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_161 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_580 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_599 ),
	.cout(Xd_0__inst_mult_14_600 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_163 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_609 ),
	.cout(Xd_0__inst_mult_9_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_164 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_614 ),
	.cout(Xd_0__inst_mult_9_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_163 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_609 ),
	.cout(Xd_0__inst_mult_8_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_164 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_614 ),
	.cout(Xd_0__inst_mult_8_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_163 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_609 ),
	.cout(Xd_0__inst_mult_11_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_164 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_614 ),
	.cout(Xd_0__inst_mult_11_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_163 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_609 ),
	.cout(Xd_0__inst_mult_10_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_164 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_614 ),
	.cout(Xd_0__inst_mult_10_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_163 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_609 ),
	.cout(Xd_0__inst_mult_5_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_164 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_614 ),
	.cout(Xd_0__inst_mult_5_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_163 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_609 ),
	.cout(Xd_0__inst_mult_4_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_164 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_614 ),
	.cout(Xd_0__inst_mult_4_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_163 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_609 ),
	.cout(Xd_0__inst_mult_7_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_164 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_614 ),
	.cout(Xd_0__inst_mult_7_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_163 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_609 ),
	.cout(Xd_0__inst_mult_6_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_164 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_614 ),
	.cout(Xd_0__inst_mult_6_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_163 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_609 ),
	.cout(Xd_0__inst_mult_1_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_164 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_614 ),
	.cout(Xd_0__inst_mult_1_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_163 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_609 ),
	.cout(Xd_0__inst_mult_0_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_164 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_614 ),
	.cout(Xd_0__inst_mult_0_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_163 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_759 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_609 ),
	.cout(Xd_0__inst_mult_3_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_164 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_614 ),
	.cout(Xd_0__inst_mult_3_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_172 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_224 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_654 ),
	.cout(Xd_0__inst_mult_2_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_173 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_659 ),
	.cout(Xd_0__inst_mult_2_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_167 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_629 ),
	.cout(Xd_0__inst_mult_29_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_168 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_634 ),
	.cout(Xd_0__inst_mult_29_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_165 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_619 ),
	.cout(Xd_0__inst_mult_28_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_166 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_624 ),
	.cout(Xd_0__inst_mult_28_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_165 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_619 ),
	.cout(Xd_0__inst_mult_31_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_166 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_624 ),
	.cout(Xd_0__inst_mult_31_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_165 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_619 ),
	.cout(Xd_0__inst_mult_30_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_166 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_624 ),
	.cout(Xd_0__inst_mult_30_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_170 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_644 ),
	.cout(Xd_0__inst_mult_25_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_171 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_649 ),
	.cout(Xd_0__inst_mult_25_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_170 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_644 ),
	.cout(Xd_0__inst_mult_27_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_171 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_649 ),
	.cout(Xd_0__inst_mult_27_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_167 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_629 ),
	.cout(Xd_0__inst_mult_21_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_168 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_634 ),
	.cout(Xd_0__inst_mult_21_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_167 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_629 ),
	.cout(Xd_0__inst_mult_20_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_168 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_634 ),
	.cout(Xd_0__inst_mult_20_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_167 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_629 ),
	.cout(Xd_0__inst_mult_23_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_168 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_634 ),
	.cout(Xd_0__inst_mult_23_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_167 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_629 ),
	.cout(Xd_0__inst_mult_22_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_168 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_634 ),
	.cout(Xd_0__inst_mult_22_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_167 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_629 ),
	.cout(Xd_0__inst_mult_17_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_168 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_634 ),
	.cout(Xd_0__inst_mult_17_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_167 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_629 ),
	.cout(Xd_0__inst_mult_16_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_168 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_634 ),
	.cout(Xd_0__inst_mult_16_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_167 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_629 ),
	.cout(Xd_0__inst_mult_19_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_168 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_634 ),
	.cout(Xd_0__inst_mult_19_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_162 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[220]),
	.datac(!Xd_0__inst_mult_18_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_604 ),
	.cout(Xd_0__inst_mult_18_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_163 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_609 ),
	.cout(Xd_0__inst_mult_18_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_164 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_614 ),
	.cout(Xd_0__inst_mult_18_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_165 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_619 ),
	.cout(Xd_0__inst_mult_13_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_166 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_624 ),
	.cout(Xd_0__inst_mult_13_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_162 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[148]),
	.datac(!Xd_0__inst_mult_12_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_604 ),
	.cout(Xd_0__inst_mult_12_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_163 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_609 ),
	.cout(Xd_0__inst_mult_12_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_164 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_614 ),
	.cout(Xd_0__inst_mult_12_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_162 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[184]),
	.datac(!Xd_0__inst_mult_15_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_604 ),
	.cout(Xd_0__inst_mult_15_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_163 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_609 ),
	.cout(Xd_0__inst_mult_15_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_164 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_614 ),
	.cout(Xd_0__inst_mult_15_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_162 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[172]),
	.datac(!Xd_0__inst_mult_14_764 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_590 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_604 ),
	.cout(Xd_0__inst_mult_14_605 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_163 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_595 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_609 ),
	.cout(Xd_0__inst_mult_14_610 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_164 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_600 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_614 ),
	.cout(Xd_0__inst_mult_14_615 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_165 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_619 ),
	.cout(Xd_0__inst_mult_9_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_166 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_624 ),
	.cout(Xd_0__inst_mult_9_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_165 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_619 ),
	.cout(Xd_0__inst_mult_8_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_166 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_624 ),
	.cout(Xd_0__inst_mult_8_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_165 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_619 ),
	.cout(Xd_0__inst_mult_11_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_166 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_624 ),
	.cout(Xd_0__inst_mult_11_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_165 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_619 ),
	.cout(Xd_0__inst_mult_10_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_166 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_624 ),
	.cout(Xd_0__inst_mult_10_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_165 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_619 ),
	.cout(Xd_0__inst_mult_5_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_166 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_624 ),
	.cout(Xd_0__inst_mult_5_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_165 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_619 ),
	.cout(Xd_0__inst_mult_4_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_166 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_624 ),
	.cout(Xd_0__inst_mult_4_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_165 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_619 ),
	.cout(Xd_0__inst_mult_7_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_166 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_624 ),
	.cout(Xd_0__inst_mult_7_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_165 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_619 ),
	.cout(Xd_0__inst_mult_6_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_166 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_624 ),
	.cout(Xd_0__inst_mult_6_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_165 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_619 ),
	.cout(Xd_0__inst_mult_1_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_166 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_624 ),
	.cout(Xd_0__inst_mult_1_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_165 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_619 ),
	.cout(Xd_0__inst_mult_0_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_166 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_624 ),
	.cout(Xd_0__inst_mult_0_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_165 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_769 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_619 ),
	.cout(Xd_0__inst_mult_3_620 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_166 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_774 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_624 ),
	.cout(Xd_0__inst_mult_3_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_174 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_219 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_664 ),
	.cout(Xd_0__inst_mult_2_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_175 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_669 ),
	.cout(Xd_0__inst_mult_2_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_169 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[353]),
	.datac(!Xd_0__inst_mult_29_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_639 ),
	.cout(Xd_0__inst_mult_29_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_170 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_644 ),
	.cout(Xd_0__inst_mult_29_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_167 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[341]),
	.datac(!Xd_0__inst_mult_28_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_629 ),
	.cout(Xd_0__inst_mult_28_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_168 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_634 ),
	.cout(Xd_0__inst_mult_28_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_167 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[377]),
	.datac(!Xd_0__inst_mult_31_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_629 ),
	.cout(Xd_0__inst_mult_31_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_168 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_634 ),
	.cout(Xd_0__inst_mult_31_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_167 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[365]),
	.datac(!Xd_0__inst_mult_30_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_629 ),
	.cout(Xd_0__inst_mult_30_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_168 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_634 ),
	.cout(Xd_0__inst_mult_30_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_172 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[305]),
	.datac(!Xd_0__inst_mult_25_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_654 ),
	.cout(Xd_0__inst_mult_25_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_173 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_659 ),
	.cout(Xd_0__inst_mult_25_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_172 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[329]),
	.datac(!Xd_0__inst_mult_27_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_654 ),
	.cout(Xd_0__inst_mult_27_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_173 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_659 ),
	.cout(Xd_0__inst_mult_27_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_169 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[257]),
	.datac(!Xd_0__inst_mult_21_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_639 ),
	.cout(Xd_0__inst_mult_21_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_170 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_644 ),
	.cout(Xd_0__inst_mult_21_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_169 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[245]),
	.datac(!Xd_0__inst_mult_20_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_639 ),
	.cout(Xd_0__inst_mult_20_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_170 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_644 ),
	.cout(Xd_0__inst_mult_20_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_169 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[281]),
	.datac(!Xd_0__inst_mult_23_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_639 ),
	.cout(Xd_0__inst_mult_23_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_170 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_644 ),
	.cout(Xd_0__inst_mult_23_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_169 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[269]),
	.datac(!Xd_0__inst_mult_22_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_639 ),
	.cout(Xd_0__inst_mult_22_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_170 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_644 ),
	.cout(Xd_0__inst_mult_22_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_169 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[209]),
	.datac(!Xd_0__inst_mult_17_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_639 ),
	.cout(Xd_0__inst_mult_17_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_170 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_644 ),
	.cout(Xd_0__inst_mult_17_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_169 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[197]),
	.datac(!Xd_0__inst_mult_16_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_639 ),
	.cout(Xd_0__inst_mult_16_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_170 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_644 ),
	.cout(Xd_0__inst_mult_16_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_169 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[233]),
	.datac(!Xd_0__inst_mult_19_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_639 ),
	.cout(Xd_0__inst_mult_19_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_170 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_644 ),
	.cout(Xd_0__inst_mult_19_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_165 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_619 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_166 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[221]),
	.datac(!Xd_0__inst_mult_18_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_624 ),
	.cout(Xd_0__inst_mult_18_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_167 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_629 ),
	.cout(Xd_0__inst_mult_18_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_167 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[161]),
	.datac(!Xd_0__inst_mult_13_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_629 ),
	.cout(Xd_0__inst_mult_13_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_168 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_634 ),
	.cout(Xd_0__inst_mult_13_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_165 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_619 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_166 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[149]),
	.datac(!Xd_0__inst_mult_12_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_624 ),
	.cout(Xd_0__inst_mult_12_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_167 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_629 ),
	.cout(Xd_0__inst_mult_12_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_165 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_619 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_166 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[185]),
	.datac(!Xd_0__inst_mult_15_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_624 ),
	.cout(Xd_0__inst_mult_15_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_167 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_629 ),
	.cout(Xd_0__inst_mult_15_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_165 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_619 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_75 (
// Equation(s):

	.dataa(!din_a[178]),
	.datab(!din_b[172]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_75_sumout ),
	.cout(Xd_0__inst_mult_14_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_166 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[173]),
	.datac(!Xd_0__inst_mult_14_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_610 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_624 ),
	.cout(Xd_0__inst_mult_14_625 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_167 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_615 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_629 ),
	.cout(Xd_0__inst_mult_14_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_167 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[113]),
	.datac(!Xd_0__inst_mult_9_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_629 ),
	.cout(Xd_0__inst_mult_9_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_168 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_634 ),
	.cout(Xd_0__inst_mult_9_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_167 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[101]),
	.datac(!Xd_0__inst_mult_8_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_629 ),
	.cout(Xd_0__inst_mult_8_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_168 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_634 ),
	.cout(Xd_0__inst_mult_8_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_167 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[137]),
	.datac(!Xd_0__inst_mult_11_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_629 ),
	.cout(Xd_0__inst_mult_11_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_168 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_634 ),
	.cout(Xd_0__inst_mult_11_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_167 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[125]),
	.datac(!Xd_0__inst_mult_10_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_629 ),
	.cout(Xd_0__inst_mult_10_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_168 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_634 ),
	.cout(Xd_0__inst_mult_10_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_167 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[65]),
	.datac(!Xd_0__inst_mult_5_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_629 ),
	.cout(Xd_0__inst_mult_5_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_168 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_634 ),
	.cout(Xd_0__inst_mult_5_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_167 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[53]),
	.datac(!Xd_0__inst_mult_4_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_629 ),
	.cout(Xd_0__inst_mult_4_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_168 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_634 ),
	.cout(Xd_0__inst_mult_4_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_167 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[89]),
	.datac(!Xd_0__inst_mult_7_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_629 ),
	.cout(Xd_0__inst_mult_7_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_168 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_634 ),
	.cout(Xd_0__inst_mult_7_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_167 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[77]),
	.datac(!Xd_0__inst_mult_6_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_629 ),
	.cout(Xd_0__inst_mult_6_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_168 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_634 ),
	.cout(Xd_0__inst_mult_6_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_167 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[17]),
	.datac(!Xd_0__inst_mult_1_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_629 ),
	.cout(Xd_0__inst_mult_1_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_168 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_634 ),
	.cout(Xd_0__inst_mult_1_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_167 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[5]),
	.datac(!Xd_0__inst_mult_0_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_629 ),
	.cout(Xd_0__inst_mult_0_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_168 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_634 ),
	.cout(Xd_0__inst_mult_0_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_167 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[41]),
	.datac(!Xd_0__inst_mult_3_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_629 ),
	.cout(Xd_0__inst_mult_3_630 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_168 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_784 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_634 ),
	.cout(Xd_0__inst_mult_3_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_176 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[29]),
	.datac(!Xd_0__inst_mult_2_214 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_674 ),
	.cout(Xd_0__inst_mult_2_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_177 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_679 ),
	.cout(Xd_0__inst_mult_2_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_171 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[354]),
	.datac(!Xd_0__inst_mult_29_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_649 ),
	.cout(Xd_0__inst_mult_29_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_172 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_654 ),
	.cout(Xd_0__inst_mult_29_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_169 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[342]),
	.datac(!Xd_0__inst_mult_28_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_639 ),
	.cout(Xd_0__inst_mult_28_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_170 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_644 ),
	.cout(Xd_0__inst_mult_28_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_169 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[378]),
	.datac(!Xd_0__inst_mult_31_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_639 ),
	.cout(Xd_0__inst_mult_31_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_170 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_644 ),
	.cout(Xd_0__inst_mult_31_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_169 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[366]),
	.datac(!Xd_0__inst_mult_30_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_639 ),
	.cout(Xd_0__inst_mult_30_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_170 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_644 ),
	.cout(Xd_0__inst_mult_30_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_174 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[306]),
	.datac(!Xd_0__inst_mult_25_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_664 ),
	.cout(Xd_0__inst_mult_25_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_175 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_669 ),
	.cout(Xd_0__inst_mult_25_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_174 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[330]),
	.datac(!Xd_0__inst_mult_27_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_664 ),
	.cout(Xd_0__inst_mult_27_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_175 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_669 ),
	.cout(Xd_0__inst_mult_27_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_171 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[258]),
	.datac(!Xd_0__inst_mult_21_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_649 ),
	.cout(Xd_0__inst_mult_21_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_172 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_654 ),
	.cout(Xd_0__inst_mult_21_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_171 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[246]),
	.datac(!Xd_0__inst_mult_20_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_649 ),
	.cout(Xd_0__inst_mult_20_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_172 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_654 ),
	.cout(Xd_0__inst_mult_20_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_171 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[282]),
	.datac(!Xd_0__inst_mult_23_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_649 ),
	.cout(Xd_0__inst_mult_23_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_172 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_654 ),
	.cout(Xd_0__inst_mult_23_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_171 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[270]),
	.datac(!Xd_0__inst_mult_22_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_649 ),
	.cout(Xd_0__inst_mult_22_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_172 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_654 ),
	.cout(Xd_0__inst_mult_22_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_171 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[210]),
	.datac(!Xd_0__inst_mult_17_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_649 ),
	.cout(Xd_0__inst_mult_17_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_172 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_654 ),
	.cout(Xd_0__inst_mult_17_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_171 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[198]),
	.datac(!Xd_0__inst_mult_16_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_649 ),
	.cout(Xd_0__inst_mult_16_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_172 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_654 ),
	.cout(Xd_0__inst_mult_16_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_171 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[234]),
	.datac(!Xd_0__inst_mult_19_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_649 ),
	.cout(Xd_0__inst_mult_19_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_172 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_654 ),
	.cout(Xd_0__inst_mult_19_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_168 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[222]),
	.datac(!Xd_0__inst_mult_18_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_634 ),
	.cout(Xd_0__inst_mult_18_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_169 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_639 ),
	.cout(Xd_0__inst_mult_18_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_169 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[162]),
	.datac(!Xd_0__inst_mult_13_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_639 ),
	.cout(Xd_0__inst_mult_13_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_170 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_644 ),
	.cout(Xd_0__inst_mult_13_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_168 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[150]),
	.datac(!Xd_0__inst_mult_12_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_634 ),
	.cout(Xd_0__inst_mult_12_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_169 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_639 ),
	.cout(Xd_0__inst_mult_12_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_168 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[186]),
	.datac(!Xd_0__inst_mult_15_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_634 ),
	.cout(Xd_0__inst_mult_15_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_169 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_639 ),
	.cout(Xd_0__inst_mult_15_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_168 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[174]),
	.datac(!Xd_0__inst_mult_14_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_625 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_634 ),
	.cout(Xd_0__inst_mult_14_635 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_169 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_639 ),
	.cout(Xd_0__inst_mult_14_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_169 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[114]),
	.datac(!Xd_0__inst_mult_9_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_639 ),
	.cout(Xd_0__inst_mult_9_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_170 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_644 ),
	.cout(Xd_0__inst_mult_9_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_169 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[102]),
	.datac(!Xd_0__inst_mult_8_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_639 ),
	.cout(Xd_0__inst_mult_8_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_170 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_644 ),
	.cout(Xd_0__inst_mult_8_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_169 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[138]),
	.datac(!Xd_0__inst_mult_11_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_639 ),
	.cout(Xd_0__inst_mult_11_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_170 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_644 ),
	.cout(Xd_0__inst_mult_11_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_169 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[126]),
	.datac(!Xd_0__inst_mult_10_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_639 ),
	.cout(Xd_0__inst_mult_10_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_170 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_644 ),
	.cout(Xd_0__inst_mult_10_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_169 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[66]),
	.datac(!Xd_0__inst_mult_5_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_639 ),
	.cout(Xd_0__inst_mult_5_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_170 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_644 ),
	.cout(Xd_0__inst_mult_5_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_169 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[54]),
	.datac(!Xd_0__inst_mult_4_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_639 ),
	.cout(Xd_0__inst_mult_4_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_170 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_644 ),
	.cout(Xd_0__inst_mult_4_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_169 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[90]),
	.datac(!Xd_0__inst_mult_7_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_639 ),
	.cout(Xd_0__inst_mult_7_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_170 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_644 ),
	.cout(Xd_0__inst_mult_7_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_169 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[78]),
	.datac(!Xd_0__inst_mult_6_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_639 ),
	.cout(Xd_0__inst_mult_6_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_170 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_644 ),
	.cout(Xd_0__inst_mult_6_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_169 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[18]),
	.datac(!Xd_0__inst_mult_1_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_639 ),
	.cout(Xd_0__inst_mult_1_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_170 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_644 ),
	.cout(Xd_0__inst_mult_1_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_169 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[6]),
	.datac(!Xd_0__inst_mult_0_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_639 ),
	.cout(Xd_0__inst_mult_0_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_170 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_644 ),
	.cout(Xd_0__inst_mult_0_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_169 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[42]),
	.datac(!Xd_0__inst_mult_3_789 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_639 ),
	.cout(Xd_0__inst_mult_3_640 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_170 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_794 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_644 ),
	.cout(Xd_0__inst_mult_3_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_178 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[30]),
	.datac(!Xd_0__inst_mult_2_210 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_684 ),
	.cout(Xd_0__inst_mult_2_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_179 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_689 ),
	.cout(Xd_0__inst_mult_2_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_173 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[355]),
	.datac(!Xd_0__inst_mult_29_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_659 ),
	.cout(Xd_0__inst_mult_29_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_174 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[356]),
	.datac(!Xd_0__inst_mult_29_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_664 ),
	.cout(Xd_0__inst_mult_29_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_171 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[343]),
	.datac(!Xd_0__inst_mult_28_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_649 ),
	.cout(Xd_0__inst_mult_28_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_172 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[344]),
	.datac(!Xd_0__inst_mult_28_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_654 ),
	.cout(Xd_0__inst_mult_28_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_171 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[379]),
	.datac(!Xd_0__inst_mult_31_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_649 ),
	.cout(Xd_0__inst_mult_31_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_172 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[380]),
	.datac(!Xd_0__inst_mult_31_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_654 ),
	.cout(Xd_0__inst_mult_31_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_171 (
// Equation(s):

	.dataa(!din_a[369]),
	.datab(!din_b[367]),
	.datac(!Xd_0__inst_mult_30_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_649 ),
	.cout(Xd_0__inst_mult_30_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_172 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[368]),
	.datac(!Xd_0__inst_mult_30_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_654 ),
	.cout(Xd_0__inst_mult_30_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_176 (
// Equation(s):

	.dataa(!din_a[309]),
	.datab(!din_b[307]),
	.datac(!Xd_0__inst_mult_25_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_674 ),
	.cout(Xd_0__inst_mult_25_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_177 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[308]),
	.datac(!Xd_0__inst_mult_25_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_679 ),
	.cout(Xd_0__inst_mult_25_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_176 (
// Equation(s):

	.dataa(!din_a[333]),
	.datab(!din_b[331]),
	.datac(!Xd_0__inst_mult_27_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_674 ),
	.cout(Xd_0__inst_mult_27_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_177 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[332]),
	.datac(!Xd_0__inst_mult_27_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_679 ),
	.cout(Xd_0__inst_mult_27_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_173 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[259]),
	.datac(!Xd_0__inst_mult_21_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_659 ),
	.cout(Xd_0__inst_mult_21_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_174 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[260]),
	.datac(!Xd_0__inst_mult_21_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_664 ),
	.cout(Xd_0__inst_mult_21_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_173 (
// Equation(s):

	.dataa(!din_a[249]),
	.datab(!din_b[247]),
	.datac(!Xd_0__inst_mult_20_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_659 ),
	.cout(Xd_0__inst_mult_20_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_174 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[248]),
	.datac(!Xd_0__inst_mult_20_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_664 ),
	.cout(Xd_0__inst_mult_20_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_173 (
// Equation(s):

	.dataa(!din_a[285]),
	.datab(!din_b[283]),
	.datac(!Xd_0__inst_mult_23_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_659 ),
	.cout(Xd_0__inst_mult_23_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_174 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[284]),
	.datac(!Xd_0__inst_mult_23_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_664 ),
	.cout(Xd_0__inst_mult_23_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_173 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[271]),
	.datac(!Xd_0__inst_mult_22_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_659 ),
	.cout(Xd_0__inst_mult_22_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_174 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[272]),
	.datac(!Xd_0__inst_mult_22_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_664 ),
	.cout(Xd_0__inst_mult_22_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_173 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[211]),
	.datac(!Xd_0__inst_mult_17_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_659 ),
	.cout(Xd_0__inst_mult_17_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_174 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[212]),
	.datac(!Xd_0__inst_mult_17_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_664 ),
	.cout(Xd_0__inst_mult_17_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_173 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[199]),
	.datac(!Xd_0__inst_mult_16_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_659 ),
	.cout(Xd_0__inst_mult_16_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_174 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[200]),
	.datac(!Xd_0__inst_mult_16_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_664 ),
	.cout(Xd_0__inst_mult_16_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_173 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[235]),
	.datac(!Xd_0__inst_mult_19_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_659 ),
	.cout(Xd_0__inst_mult_19_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_174 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[236]),
	.datac(!Xd_0__inst_mult_19_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_664 ),
	.cout(Xd_0__inst_mult_19_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_170 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[223]),
	.datac(!Xd_0__inst_mult_18_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_644 ),
	.cout(Xd_0__inst_mult_18_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_171 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[224]),
	.datac(!Xd_0__inst_mult_18_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_649 ),
	.cout(Xd_0__inst_mult_18_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_171 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[163]),
	.datac(!Xd_0__inst_mult_13_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_649 ),
	.cout(Xd_0__inst_mult_13_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_172 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[164]),
	.datac(!Xd_0__inst_mult_13_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_654 ),
	.cout(Xd_0__inst_mult_13_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_170 (
// Equation(s):

	.dataa(!din_a[153]),
	.datab(!din_b[151]),
	.datac(!Xd_0__inst_mult_12_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_644 ),
	.cout(Xd_0__inst_mult_12_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_171 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[152]),
	.datac(!Xd_0__inst_mult_12_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_649 ),
	.cout(Xd_0__inst_mult_12_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_170 (
// Equation(s):

	.dataa(!din_a[189]),
	.datab(!din_b[187]),
	.datac(!Xd_0__inst_mult_15_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_644 ),
	.cout(Xd_0__inst_mult_15_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_171 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[188]),
	.datac(!Xd_0__inst_mult_15_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_649 ),
	.cout(Xd_0__inst_mult_15_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_170 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[175]),
	.datac(!Xd_0__inst_mult_14_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_635 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_644 ),
	.cout(Xd_0__inst_mult_14_645 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_171 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[176]),
	.datac(!Xd_0__inst_mult_14_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_649 ),
	.cout(Xd_0__inst_mult_14_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_171 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[115]),
	.datac(!Xd_0__inst_mult_9_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_649 ),
	.cout(Xd_0__inst_mult_9_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_172 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[116]),
	.datac(!Xd_0__inst_mult_9_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_654 ),
	.cout(Xd_0__inst_mult_9_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_171 (
// Equation(s):

	.dataa(!din_a[105]),
	.datab(!din_b[103]),
	.datac(!Xd_0__inst_mult_8_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_649 ),
	.cout(Xd_0__inst_mult_8_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_172 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[104]),
	.datac(!Xd_0__inst_mult_8_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_654 ),
	.cout(Xd_0__inst_mult_8_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_171 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[139]),
	.datac(!Xd_0__inst_mult_11_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_649 ),
	.cout(Xd_0__inst_mult_11_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_172 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[140]),
	.datac(!Xd_0__inst_mult_11_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_654 ),
	.cout(Xd_0__inst_mult_11_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_171 (
// Equation(s):

	.dataa(!din_a[129]),
	.datab(!din_b[127]),
	.datac(!Xd_0__inst_mult_10_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_649 ),
	.cout(Xd_0__inst_mult_10_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_172 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(!Xd_0__inst_mult_10_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_654 ),
	.cout(Xd_0__inst_mult_10_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_171 (
// Equation(s):

	.dataa(!din_a[69]),
	.datab(!din_b[67]),
	.datac(!Xd_0__inst_mult_5_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_649 ),
	.cout(Xd_0__inst_mult_5_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_172 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[68]),
	.datac(!Xd_0__inst_mult_5_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_654 ),
	.cout(Xd_0__inst_mult_5_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_171 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[55]),
	.datac(!Xd_0__inst_mult_4_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_649 ),
	.cout(Xd_0__inst_mult_4_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_172 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(!Xd_0__inst_mult_4_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_654 ),
	.cout(Xd_0__inst_mult_4_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_171 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[91]),
	.datac(!Xd_0__inst_mult_7_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_649 ),
	.cout(Xd_0__inst_mult_7_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_172 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[92]),
	.datac(!Xd_0__inst_mult_7_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_654 ),
	.cout(Xd_0__inst_mult_7_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_171 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[79]),
	.datac(!Xd_0__inst_mult_6_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_649 ),
	.cout(Xd_0__inst_mult_6_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_172 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[80]),
	.datac(!Xd_0__inst_mult_6_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_654 ),
	.cout(Xd_0__inst_mult_6_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_171 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[19]),
	.datac(!Xd_0__inst_mult_1_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_649 ),
	.cout(Xd_0__inst_mult_1_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_172 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[20]),
	.datac(!Xd_0__inst_mult_1_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_654 ),
	.cout(Xd_0__inst_mult_1_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_171 (
// Equation(s):

	.dataa(!din_a[9]),
	.datab(!din_b[7]),
	.datac(!Xd_0__inst_mult_0_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_649 ),
	.cout(Xd_0__inst_mult_0_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_172 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(!Xd_0__inst_mult_0_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_654 ),
	.cout(Xd_0__inst_mult_0_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_171 (
// Equation(s):

	.dataa(!din_a[45]),
	.datab(!din_b[43]),
	.datac(!Xd_0__inst_mult_3_799 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_640 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_649 ),
	.cout(Xd_0__inst_mult_3_650 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_172 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(!Xd_0__inst_mult_3_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_654 ),
	.cout(Xd_0__inst_mult_3_655 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_180 (
// Equation(s):

	.dataa(!din_a[33]),
	.datab(!din_b[31]),
	.datac(!Xd_0__inst_mult_2_205 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_694 ),
	.cout(Xd_0__inst_mult_2_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_181 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[32]),
	.datac(!Xd_0__inst_mult_2_804 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_699 ),
	.cout(Xd_0__inst_mult_2_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_176 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[357]),
	.datac(!Xd_0__inst_mult_29_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_674 ),
	.cout(Xd_0__inst_mult_29_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_174 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[345]),
	.datac(!Xd_0__inst_mult_28_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_664 ),
	.cout(Xd_0__inst_mult_28_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_174 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[381]),
	.datac(!Xd_0__inst_mult_31_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_664 ),
	.cout(Xd_0__inst_mult_31_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_174 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[369]),
	.datac(!Xd_0__inst_mult_30_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_664 ),
	.cout(Xd_0__inst_mult_30_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_179 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[309]),
	.datac(!Xd_0__inst_mult_25_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_689 ),
	.cout(Xd_0__inst_mult_25_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_179 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[333]),
	.datac(!Xd_0__inst_mult_27_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_689 ),
	.cout(Xd_0__inst_mult_27_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_176 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[261]),
	.datac(!Xd_0__inst_mult_21_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_674 ),
	.cout(Xd_0__inst_mult_21_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_176 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[249]),
	.datac(!Xd_0__inst_mult_20_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_674 ),
	.cout(Xd_0__inst_mult_20_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_176 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[285]),
	.datac(!Xd_0__inst_mult_23_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_674 ),
	.cout(Xd_0__inst_mult_23_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_176 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[273]),
	.datac(!Xd_0__inst_mult_22_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_674 ),
	.cout(Xd_0__inst_mult_22_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_176 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[213]),
	.datac(!Xd_0__inst_mult_17_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_674 ),
	.cout(Xd_0__inst_mult_17_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_176 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[201]),
	.datac(!Xd_0__inst_mult_16_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_674 ),
	.cout(Xd_0__inst_mult_16_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_176 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[237]),
	.datac(!Xd_0__inst_mult_19_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_674 ),
	.cout(Xd_0__inst_mult_19_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_172 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_654 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_173 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[225]),
	.datac(!Xd_0__inst_mult_18_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_659 ),
	.cout(Xd_0__inst_mult_18_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_174 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[165]),
	.datac(!Xd_0__inst_mult_13_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_664 ),
	.cout(Xd_0__inst_mult_13_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_172 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_654 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_173 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[153]),
	.datac(!Xd_0__inst_mult_12_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_659 ),
	.cout(Xd_0__inst_mult_12_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_172 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_654 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_173 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[189]),
	.datac(!Xd_0__inst_mult_15_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_659 ),
	.cout(Xd_0__inst_mult_15_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_172 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_645 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_654 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_173 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[177]),
	.datac(!Xd_0__inst_mult_14_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_659 ),
	.cout(Xd_0__inst_mult_14_660 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_174 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[117]),
	.datac(!Xd_0__inst_mult_9_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_664 ),
	.cout(Xd_0__inst_mult_9_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_174 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[105]),
	.datac(!Xd_0__inst_mult_8_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_664 ),
	.cout(Xd_0__inst_mult_8_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_174 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[141]),
	.datac(!Xd_0__inst_mult_11_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_664 ),
	.cout(Xd_0__inst_mult_11_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_174 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[129]),
	.datac(!Xd_0__inst_mult_10_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_664 ),
	.cout(Xd_0__inst_mult_10_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_174 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[69]),
	.datac(!Xd_0__inst_mult_5_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_664 ),
	.cout(Xd_0__inst_mult_5_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_174 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[57]),
	.datac(!Xd_0__inst_mult_4_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_664 ),
	.cout(Xd_0__inst_mult_4_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_174 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[93]),
	.datac(!Xd_0__inst_mult_7_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_664 ),
	.cout(Xd_0__inst_mult_7_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_174 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[81]),
	.datac(!Xd_0__inst_mult_6_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_664 ),
	.cout(Xd_0__inst_mult_6_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_174 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[21]),
	.datac(!Xd_0__inst_mult_1_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_664 ),
	.cout(Xd_0__inst_mult_1_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_174 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[9]),
	.datac(!Xd_0__inst_mult_0_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_664 ),
	.cout(Xd_0__inst_mult_0_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_173 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_659 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_174 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[45]),
	.datac(!Xd_0__inst_mult_3_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_655 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_664 ),
	.cout(Xd_0__inst_mult_3_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_182 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_704 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_183 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[33]),
	.datac(!Xd_0__inst_mult_2_809 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_709 ),
	.cout(Xd_0__inst_mult_2_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_29_177 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[358]),
	.datac(!Xd_0__inst_mult_29_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_679 ),
	.cout(Xd_0__inst_mult_29_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_80 (
// Equation(s):

	.dataa(!din_a[357]),
	.datab(!din_b[357]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_36 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_80_sumout ),
	.cout(Xd_0__inst_mult_29_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_28_175 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[346]),
	.datac(!Xd_0__inst_mult_28_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_669 ),
	.cout(Xd_0__inst_mult_28_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_80 (
// Equation(s):

	.dataa(!din_a[345]),
	.datab(!din_b[345]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_80_sumout ),
	.cout(Xd_0__inst_mult_28_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_31_175 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[382]),
	.datac(!Xd_0__inst_mult_31_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_669 ),
	.cout(Xd_0__inst_mult_31_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_80 (
// Equation(s):

	.dataa(!din_a[381]),
	.datab(!din_b[381]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_80_sumout ),
	.cout(Xd_0__inst_mult_31_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_30_175 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[370]),
	.datac(!Xd_0__inst_mult_30_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_669 ),
	.cout(Xd_0__inst_mult_30_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_25_180 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[310]),
	.datac(!Xd_0__inst_mult_25_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_694 ),
	.cout(Xd_0__inst_mult_25_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_27_180 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[334]),
	.datac(!Xd_0__inst_mult_18_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_694 ),
	.cout(Xd_0__inst_mult_27_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_21_177 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[262]),
	.datac(!Xd_0__inst_mult_21_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_679 ),
	.cout(Xd_0__inst_mult_21_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_80 (
// Equation(s):

	.dataa(!din_a[261]),
	.datab(!din_b[261]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_41 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_80_sumout ),
	.cout(Xd_0__inst_mult_21_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_20_177 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[250]),
	.datac(!Xd_0__inst_mult_20_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_679 ),
	.cout(Xd_0__inst_mult_20_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_23_177 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[286]),
	.datac(!Xd_0__inst_mult_23_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_679 ),
	.cout(Xd_0__inst_mult_23_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_22_177 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[274]),
	.datac(!Xd_0__inst_mult_22_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_679 ),
	.cout(Xd_0__inst_mult_22_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_80 (
// Equation(s):

	.dataa(!din_a[273]),
	.datab(!din_b[273]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_80_sumout ),
	.cout(Xd_0__inst_mult_22_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_17_177 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[214]),
	.datac(!Xd_0__inst_mult_17_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_679 ),
	.cout(Xd_0__inst_mult_17_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_80 (
// Equation(s):

	.dataa(!din_a[213]),
	.datab(!din_b[213]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_80_sumout ),
	.cout(Xd_0__inst_mult_17_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_16_177 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[202]),
	.datac(!Xd_0__inst_mult_16_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_679 ),
	.cout(Xd_0__inst_mult_16_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_75 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[201]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_75_sumout ),
	.cout(Xd_0__inst_mult_16_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_19_177 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[238]),
	.datac(!Xd_0__inst_mult_19_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_679 ),
	.cout(Xd_0__inst_mult_19_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_75 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[237]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_75_sumout ),
	.cout(Xd_0__inst_mult_19_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_18_174 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[226]),
	.datac(!Xd_0__inst_mult_15_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_664 ),
	.cout(Xd_0__inst_mult_18_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_75 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[225]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_75_sumout ),
	.cout(Xd_0__inst_mult_18_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_13_175 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[166]),
	.datac(!Xd_0__inst_mult_12_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_669 ),
	.cout(Xd_0__inst_mult_13_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_75 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_75_sumout ),
	.cout(Xd_0__inst_mult_13_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_12_174 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[154]),
	.datac(!Xd_0__inst_mult_2_779 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_664 ),
	.cout(Xd_0__inst_mult_12_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_15_174 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[190]),
	.datac(!Xd_0__inst_mult_3_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_664 ),
	.cout(Xd_0__inst_mult_15_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_14_174 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[178]),
	.datac(!Xd_0__inst_mult_0_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_660 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_664 ),
	.cout(Xd_0__inst_mult_14_665 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_9_175 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[118]),
	.datac(!Xd_0__inst_mult_1_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_669 ),
	.cout(Xd_0__inst_mult_9_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_75 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_75_sumout ),
	.cout(Xd_0__inst_mult_9_76 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_8_175 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[106]),
	.datac(!Xd_0__inst_mult_6_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_669 ),
	.cout(Xd_0__inst_mult_8_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_11_175 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[142]),
	.datac(!Xd_0__inst_mult_7_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_669 ),
	.cout(Xd_0__inst_mult_11_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_10_175 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[130]),
	.datac(!Xd_0__inst_mult_4_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_669 ),
	.cout(Xd_0__inst_mult_10_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_5_175 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[70]),
	.datac(!Xd_0__inst_mult_5_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_669 ),
	.cout(Xd_0__inst_mult_5_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_4_175 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[58]),
	.datac(!Xd_0__inst_mult_10_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_669 ),
	.cout(Xd_0__inst_mult_4_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_7_175 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[94]),
	.datac(!Xd_0__inst_mult_11_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_669 ),
	.cout(Xd_0__inst_mult_7_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_6_175 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[82]),
	.datac(!Xd_0__inst_mult_8_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_669 ),
	.cout(Xd_0__inst_mult_6_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_1_175 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[22]),
	.datac(!Xd_0__inst_mult_9_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_669 ),
	.cout(Xd_0__inst_mult_1_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_0_175 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[10]),
	.datac(!Xd_0__inst_mult_14_744 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_669 ),
	.cout(Xd_0__inst_mult_0_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_3_175 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[46]),
	.datac(!Xd_0__inst_mult_27_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_669 ),
	.cout(Xd_0__inst_mult_3_670 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000001011E1E),
	.shared_arith("off")
) Xd_0__inst_mult_2_184 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[34]),
	.datac(!Xd_0__inst_mult_13_754 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_714 ),
	.cout(Xd_0__inst_mult_2_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_181 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_699 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_181 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_699 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_80 (
// Equation(s):

	.dataa(!din_a[201]),
	.datab(!din_b[202]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_80_sumout ),
	.cout(Xd_0__inst_mult_16_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_178 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_684 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_80 (
// Equation(s):

	.dataa(!din_a[237]),
	.datab(!din_b[238]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_80_sumout ),
	.cout(Xd_0__inst_mult_19_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_80 (
// Equation(s):

	.dataa(!din_a[225]),
	.datab(!din_b[226]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_80_sumout ),
	.cout(Xd_0__inst_mult_18_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_80 (
// Equation(s):

	.dataa(!din_a[165]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_80_sumout ),
	.cout(Xd_0__inst_mult_13_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_175 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_665 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_669 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_80 (
// Equation(s):

	.dataa(!din_a[177]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_80_sumout ),
	.cout(Xd_0__inst_mult_14_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_80 (
// Equation(s):

	.dataa(!din_a[117]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_80_sumout ),
	.cout(Xd_0__inst_mult_9_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_80 (
// Equation(s):

	.dataa(!din_a[141]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_76 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_80_sumout ),
	.cout(Xd_0__inst_mult_11_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_80 (
// Equation(s):

	.dataa(!din_a[57]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_80_sumout ),
	.cout(Xd_0__inst_mult_4_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_80 (
// Equation(s):

	.dataa(!din_a[93]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_80_sumout ),
	.cout(Xd_0__inst_mult_7_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_80 (
// Equation(s):

	.dataa(!din_a[81]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_80_sumout ),
	.cout(Xd_0__inst_mult_6_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_80 (
// Equation(s):

	.dataa(!din_a[21]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_81 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_80_sumout ),
	.cout(Xd_0__inst_mult_1_81 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_176 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_670 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_674 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_2_185 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_719 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_177 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[112]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_679 ),
	.cout(Xd_0__inst_mult_9_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_177 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[100]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_679 ),
	.cout(Xd_0__inst_mult_8_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_179 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[255]),
	.datac(!din_a[258]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_689 ),
	.cout(Xd_0__inst_mult_21_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_177 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[136]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_679 ),
	.cout(Xd_0__inst_mult_11_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_177 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[124]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_679 ),
	.cout(Xd_0__inst_mult_10_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_179 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[243]),
	.datac(!din_a[246]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_689 ),
	.cout(Xd_0__inst_mult_20_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_182 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[303]),
	.datac(!din_a[303]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_704 ),
	.cout(Xd_0__inst_mult_25_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_177 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[40]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_679 ),
	.cout(Xd_0__inst_mult_3_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_177 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_679 ),
	.cout(Xd_0__inst_mult_0_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_179 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[279]),
	.datac(!din_a[282]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_689 ),
	.cout(Xd_0__inst_mult_23_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_177 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_679 ),
	.cout(Xd_0__inst_mult_6_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_177 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_679 ),
	.cout(Xd_0__inst_mult_1_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_179 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[267]),
	.datac(!din_a[270]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_689 ),
	.cout(Xd_0__inst_mult_22_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_196 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[291]),
	.datac(!din_a[291]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_774 ),
	.cout(Xd_0__inst_mult_24_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_196 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[318]),
	.datac(!din_a[315]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_774 ),
	.cout(Xd_0__inst_mult_26_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_177 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_679 ),
	.cout(Xd_0__inst_mult_7_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_177 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[52]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_679 ),
	.cout(Xd_0__inst_mult_4_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_179 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[231]),
	.datac(!din_a[234]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_689 ),
	.cout(Xd_0__inst_mult_19_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_177 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[364]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_679 ),
	.cout(Xd_0__inst_mult_30_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_177 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[64]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_679 ),
	.cout(Xd_0__inst_mult_5_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_179 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[207]),
	.datac(!din_a[210]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_689 ),
	.cout(Xd_0__inst_mult_17_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_182 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[327]),
	.datac(!din_a[327]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_704 ),
	.cout(Xd_0__inst_mult_27_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_177 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[160]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_679 ),
	.cout(Xd_0__inst_mult_13_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_186 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_724 ),
	.cout(Xd_0__inst_mult_2_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_179 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[195]),
	.datac(!din_a[198]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_689 ),
	.cout(Xd_0__inst_mult_16_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_177 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[340]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_679 ),
	.cout(Xd_0__inst_mult_28_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_177 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[376]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_679 ),
	.cout(Xd_0__inst_mult_31_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_179 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[351]),
	.datac(!din_a[354]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_689 ),
	.cout(Xd_0__inst_mult_29_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_197 (
// Equation(s):

	.dataa(!din_a[316]),
	.datab(!din_b[315]),
	.datac(!din_a[315]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_779 ),
	.cout(Xd_0__inst_mult_26_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_197 (
// Equation(s):

	.dataa(!din_a[292]),
	.datab(!din_b[294]),
	.datac(!din_a[291]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_779 ),
	.cout(Xd_0__inst_mult_24_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_180 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[351]),
	.datac(!din_a[349]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_694 ),
	.cout(Xd_0__inst_mult_29_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_29_181 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[351]),
	.datac(!din_a[349]),
	.datad(!din_b[350]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_178 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[339]),
	.datac(!din_a[337]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_684 ),
	.cout(Xd_0__inst_mult_28_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_28_179 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[339]),
	.datac(!din_a[337]),
	.datad(!din_b[338]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_178 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[375]),
	.datac(!din_a[373]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_684 ),
	.cout(Xd_0__inst_mult_31_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_31_179 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[375]),
	.datac(!din_a[373]),
	.datad(!din_b[374]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_178 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[363]),
	.datac(!din_a[361]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_684 ),
	.cout(Xd_0__inst_mult_30_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_30_179 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[363]),
	.datac(!din_a[361]),
	.datad(!din_b[362]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_183 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[303]),
	.datac(!din_a[301]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_709 ),
	.cout(Xd_0__inst_mult_25_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_25_184 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[303]),
	.datac(!din_a[301]),
	.datad(!din_b[302]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_198 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[291]),
	.datac(!din_a[289]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_784 ),
	.cout(Xd_0__inst_mult_24_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_24_199 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[291]),
	.datac(!din_a[289]),
	.datad(!din_b[290]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_183 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[327]),
	.datac(!din_a[325]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_460 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_709 ),
	.cout(Xd_0__inst_mult_27_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_27_184 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[327]),
	.datac(!din_a[325]),
	.datad(!din_b[326]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_198 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[315]),
	.datac(!din_a[313]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_650 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_784 ),
	.cout(Xd_0__inst_mult_26_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_26_199 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[315]),
	.datac(!din_a[313]),
	.datad(!din_b[314]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_180 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[255]),
	.datac(!din_a[253]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_694 ),
	.cout(Xd_0__inst_mult_21_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_21_181 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[255]),
	.datac(!din_a[253]),
	.datad(!din_b[254]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_180 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[243]),
	.datac(!din_a[241]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_694 ),
	.cout(Xd_0__inst_mult_20_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_20_181 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[243]),
	.datac(!din_a[241]),
	.datad(!din_b[242]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_180 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[279]),
	.datac(!din_a[277]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_694 ),
	.cout(Xd_0__inst_mult_23_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_23_181 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[279]),
	.datac(!din_a[277]),
	.datad(!din_b[278]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_180 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[267]),
	.datac(!din_a[265]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_694 ),
	.cout(Xd_0__inst_mult_22_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_22_181 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[267]),
	.datac(!din_a[265]),
	.datad(!din_b[266]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_180 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[207]),
	.datac(!din_a[205]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_694 ),
	.cout(Xd_0__inst_mult_17_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_17_181 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[207]),
	.datac(!din_a[205]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_180 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[195]),
	.datac(!din_a[193]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_694 ),
	.cout(Xd_0__inst_mult_16_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_16_181 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[195]),
	.datac(!din_a[193]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_180 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[231]),
	.datac(!din_a[229]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_400 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_694 ),
	.cout(Xd_0__inst_mult_19_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_19_181 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[231]),
	.datac(!din_a[229]),
	.datad(!din_b[230]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_176 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[219]),
	.datac(!din_a[217]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_674 ),
	.cout(Xd_0__inst_mult_18_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_18_177 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[219]),
	.datac(!din_a[217]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_178 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[159]),
	.datac(!din_a[157]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_684 ),
	.cout(Xd_0__inst_mult_13_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_13_179 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[159]),
	.datac(!din_a[157]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_176 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[147]),
	.datac(!din_a[145]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_674 ),
	.cout(Xd_0__inst_mult_12_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_12_177 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[147]),
	.datac(!din_a[145]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_176 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[183]),
	.datac(!din_a[181]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_674 ),
	.cout(Xd_0__inst_mult_15_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_15_177 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[183]),
	.datac(!din_a[181]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_176 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[171]),
	.datac(!din_a[169]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_335 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_674 ),
	.cout(Xd_0__inst_mult_14_675 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_14_177 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[171]),
	.datac(!din_a[169]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_680 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_178 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[111]),
	.datac(!din_a[109]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_684 ),
	.cout(Xd_0__inst_mult_9_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_9_179 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[111]),
	.datac(!din_a[109]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_178 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[99]),
	.datac(!din_a[97]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_684 ),
	.cout(Xd_0__inst_mult_8_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_8_179 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[99]),
	.datac(!din_a[97]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_178 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[135]),
	.datac(!din_a[133]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_684 ),
	.cout(Xd_0__inst_mult_11_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_11_179 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[135]),
	.datac(!din_a[133]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_178 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[123]),
	.datac(!din_a[121]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_684 ),
	.cout(Xd_0__inst_mult_10_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_10_179 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[123]),
	.datac(!din_a[121]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_178 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[63]),
	.datac(!din_a[61]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_684 ),
	.cout(Xd_0__inst_mult_5_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_5_179 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[63]),
	.datac(!din_a[61]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_178 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[51]),
	.datac(!din_a[49]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_684 ),
	.cout(Xd_0__inst_mult_4_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_4_179 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[51]),
	.datac(!din_a[49]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_178 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[87]),
	.datac(!din_a[85]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_684 ),
	.cout(Xd_0__inst_mult_7_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_7_179 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[87]),
	.datac(!din_a[85]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_178 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[75]),
	.datac(!din_a[73]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_684 ),
	.cout(Xd_0__inst_mult_6_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_6_179 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[75]),
	.datac(!din_a[73]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_178 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[15]),
	.datac(!din_a[13]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_684 ),
	.cout(Xd_0__inst_mult_1_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_1_179 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[15]),
	.datac(!din_a[13]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_178 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[3]),
	.datac(!din_a[1]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_684 ),
	.cout(Xd_0__inst_mult_0_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_0_179 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[3]),
	.datac(!din_a[1]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_178 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[39]),
	.datac(!din_a[37]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_360 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_684 ),
	.cout(Xd_0__inst_mult_3_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_3_179 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[39]),
	.datac(!din_a[37]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_187 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[27]),
	.datac(!din_a[25]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_420 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_729 ),
	.cout(Xd_0__inst_mult_2_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_2_188 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[27]),
	.datac(!din_a[25]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_182 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[351]),
	.datac(!din_a[350]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_704 ),
	.cout(Xd_0__inst_mult_29_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_180 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[339]),
	.datac(!din_a[338]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_694 ),
	.cout(Xd_0__inst_mult_28_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_180 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[375]),
	.datac(!din_a[374]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_694 ),
	.cout(Xd_0__inst_mult_31_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_180 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[363]),
	.datac(!din_a[362]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_694 ),
	.cout(Xd_0__inst_mult_30_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_185 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[303]),
	.datac(!din_a[302]),
	.datad(!din_b[304]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_719 ),
	.cout(Xd_0__inst_mult_25_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_200 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[291]),
	.datac(!din_a[290]),
	.datad(!din_b[292]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_794 ),
	.cout(Xd_0__inst_mult_24_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_185 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[327]),
	.datac(!din_a[326]),
	.datad(!din_b[328]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_719 ),
	.cout(Xd_0__inst_mult_27_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_200 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[315]),
	.datac(!din_a[314]),
	.datad(!din_b[316]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_794 ),
	.cout(Xd_0__inst_mult_26_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_182 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[255]),
	.datac(!din_a[254]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_704 ),
	.cout(Xd_0__inst_mult_21_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_182 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[243]),
	.datac(!din_a[242]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_704 ),
	.cout(Xd_0__inst_mult_20_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_182 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[279]),
	.datac(!din_a[278]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_704 ),
	.cout(Xd_0__inst_mult_23_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_182 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[267]),
	.datac(!din_a[266]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_704 ),
	.cout(Xd_0__inst_mult_22_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_182 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[207]),
	.datac(!din_a[206]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_704 ),
	.cout(Xd_0__inst_mult_17_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_182 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[195]),
	.datac(!din_a[194]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_704 ),
	.cout(Xd_0__inst_mult_16_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_182 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[231]),
	.datac(!din_a[230]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_704 ),
	.cout(Xd_0__inst_mult_19_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_178 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[219]),
	.datac(!din_a[218]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_684 ),
	.cout(Xd_0__inst_mult_18_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_180 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[159]),
	.datac(!din_a[158]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_694 ),
	.cout(Xd_0__inst_mult_13_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_178 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[147]),
	.datac(!din_a[146]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_684 ),
	.cout(Xd_0__inst_mult_12_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_178 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[183]),
	.datac(!din_a[182]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_684 ),
	.cout(Xd_0__inst_mult_15_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_178 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[171]),
	.datac(!din_a[170]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_675 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_684 ),
	.cout(Xd_0__inst_mult_14_685 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_180 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[111]),
	.datac(!din_a[110]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_694 ),
	.cout(Xd_0__inst_mult_9_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_180 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[99]),
	.datac(!din_a[98]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_694 ),
	.cout(Xd_0__inst_mult_8_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_180 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[135]),
	.datac(!din_a[134]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_694 ),
	.cout(Xd_0__inst_mult_11_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_180 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[123]),
	.datac(!din_a[122]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_694 ),
	.cout(Xd_0__inst_mult_10_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_180 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[63]),
	.datac(!din_a[62]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_694 ),
	.cout(Xd_0__inst_mult_5_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_180 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_694 ),
	.cout(Xd_0__inst_mult_4_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_180 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[87]),
	.datac(!din_a[86]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_694 ),
	.cout(Xd_0__inst_mult_7_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_180 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[75]),
	.datac(!din_a[74]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_694 ),
	.cout(Xd_0__inst_mult_6_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_180 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[15]),
	.datac(!din_a[14]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_694 ),
	.cout(Xd_0__inst_mult_1_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_180 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[3]),
	.datac(!din_a[2]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_694 ),
	.cout(Xd_0__inst_mult_0_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_180 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[39]),
	.datac(!din_a[38]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_694 ),
	.cout(Xd_0__inst_mult_3_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_189 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[27]),
	.datac(!din_a[26]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_739 ),
	.cout(Xd_0__inst_mult_2_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_183 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[351]),
	.datac(!din_a[351]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_709 ),
	.cout(Xd_0__inst_mult_29_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_181 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[339]),
	.datac(!din_a[339]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_699 ),
	.cout(Xd_0__inst_mult_28_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_181 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[375]),
	.datac(!din_a[375]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_699 ),
	.cout(Xd_0__inst_mult_31_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_181 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[363]),
	.datac(!din_a[363]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_699 ),
	.cout(Xd_0__inst_mult_30_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_183 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[255]),
	.datac(!din_a[255]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_709 ),
	.cout(Xd_0__inst_mult_21_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_183 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[243]),
	.datac(!din_a[243]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_709 ),
	.cout(Xd_0__inst_mult_20_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_183 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[279]),
	.datac(!din_a[279]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_709 ),
	.cout(Xd_0__inst_mult_23_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_183 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[267]),
	.datac(!din_a[267]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_709 ),
	.cout(Xd_0__inst_mult_22_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_183 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[207]),
	.datac(!din_a[207]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_709 ),
	.cout(Xd_0__inst_mult_17_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_183 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[195]),
	.datac(!din_a[195]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_709 ),
	.cout(Xd_0__inst_mult_16_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_183 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[231]),
	.datac(!din_a[231]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_709 ),
	.cout(Xd_0__inst_mult_19_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_179 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[219]),
	.datac(!din_a[219]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_689 ),
	.cout(Xd_0__inst_mult_18_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_181 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[159]),
	.datac(!din_a[159]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_699 ),
	.cout(Xd_0__inst_mult_13_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_179 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[147]),
	.datac(!din_a[147]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_689 ),
	.cout(Xd_0__inst_mult_12_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_179 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[183]),
	.datac(!din_a[183]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_689 ),
	.cout(Xd_0__inst_mult_15_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_179 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[171]),
	.datac(!din_a[171]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_685 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_689 ),
	.cout(Xd_0__inst_mult_14_690 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_181 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[111]),
	.datac(!din_a[111]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_699 ),
	.cout(Xd_0__inst_mult_9_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_181 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[99]),
	.datac(!din_a[99]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_699 ),
	.cout(Xd_0__inst_mult_8_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_181 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[135]),
	.datac(!din_a[135]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_699 ),
	.cout(Xd_0__inst_mult_11_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_181 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[123]),
	.datac(!din_a[123]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_699 ),
	.cout(Xd_0__inst_mult_10_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_181 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[63]),
	.datac(!din_a[63]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_699 ),
	.cout(Xd_0__inst_mult_5_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_181 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[51]),
	.datac(!din_a[51]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_699 ),
	.cout(Xd_0__inst_mult_4_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_181 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[87]),
	.datac(!din_a[87]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_699 ),
	.cout(Xd_0__inst_mult_7_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_181 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[75]),
	.datac(!din_a[75]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_699 ),
	.cout(Xd_0__inst_mult_6_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_181 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[15]),
	.datac(!din_a[15]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_699 ),
	.cout(Xd_0__inst_mult_1_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_181 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[3]),
	.datac(!din_a[3]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_699 ),
	.cout(Xd_0__inst_mult_0_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_181 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[39]),
	.datac(!din_a[39]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_699 ),
	.cout(Xd_0__inst_mult_3_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_190 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[27]),
	.datac(!din_a[27]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_744 ),
	.cout(Xd_0__inst_mult_2_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_184 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[351]),
	.datac(!din_a[352]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_714 ),
	.cout(Xd_0__inst_mult_29_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_185 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[354]),
	.datac(!din_a[349]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_719 ),
	.cout(Xd_0__inst_mult_29_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_29_186 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[354]),
	.datac(!din_a[349]),
	.datad(!din_b[353]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_182 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[339]),
	.datac(!din_a[340]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_704 ),
	.cout(Xd_0__inst_mult_28_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_183 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[342]),
	.datac(!din_a[337]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_709 ),
	.cout(Xd_0__inst_mult_28_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_28_184 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[342]),
	.datac(!din_a[337]),
	.datad(!din_b[341]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_182 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[375]),
	.datac(!din_a[376]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_704 ),
	.cout(Xd_0__inst_mult_31_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_183 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[378]),
	.datac(!din_a[373]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_709 ),
	.cout(Xd_0__inst_mult_31_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_31_184 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[378]),
	.datac(!din_a[373]),
	.datad(!din_b[377]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_182 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[363]),
	.datac(!din_a[364]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_704 ),
	.cout(Xd_0__inst_mult_30_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_183 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[366]),
	.datac(!din_a[361]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_709 ),
	.cout(Xd_0__inst_mult_30_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_30_184 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[366]),
	.datac(!din_a[361]),
	.datad(!din_b[365]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_186 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[306]),
	.datac(!din_a[301]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_724 ),
	.cout(Xd_0__inst_mult_25_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_25_187 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[306]),
	.datac(!din_a[301]),
	.datad(!din_b[305]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_201 (
// Equation(s):

	.dataa(!din_a[290]),
	.datab(!din_b[294]),
	.datac(!din_a[289]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_799 ),
	.cout(Xd_0__inst_mult_24_800 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_24_202 (
// Equation(s):

	.dataa(!din_a[288]),
	.datab(!din_b[294]),
	.datac(!din_a[289]),
	.datad(!din_b[293]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_186 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[330]),
	.datac(!din_a[325]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_490 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_724 ),
	.cout(Xd_0__inst_mult_27_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_27_187 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[330]),
	.datac(!din_a[325]),
	.datad(!din_b[329]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_201 (
// Equation(s):

	.dataa(!din_a[314]),
	.datab(!din_b[318]),
	.datac(!din_a[313]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_680 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_799 ),
	.cout(Xd_0__inst_mult_26_800 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_26_202 (
// Equation(s):

	.dataa(!din_a[312]),
	.datab(!din_b[318]),
	.datac(!din_a[313]),
	.datad(!din_b[317]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_184 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[255]),
	.datac(!din_a[256]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_714 ),
	.cout(Xd_0__inst_mult_21_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_185 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[258]),
	.datac(!din_a[253]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_719 ),
	.cout(Xd_0__inst_mult_21_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_21_186 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[258]),
	.datac(!din_a[253]),
	.datad(!din_b[257]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_184 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[243]),
	.datac(!din_a[244]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_714 ),
	.cout(Xd_0__inst_mult_20_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_185 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[246]),
	.datac(!din_a[241]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_719 ),
	.cout(Xd_0__inst_mult_20_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_20_186 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[246]),
	.datac(!din_a[241]),
	.datad(!din_b[245]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_184 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[279]),
	.datac(!din_a[280]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_714 ),
	.cout(Xd_0__inst_mult_23_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_185 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[282]),
	.datac(!din_a[277]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_719 ),
	.cout(Xd_0__inst_mult_23_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_23_186 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[282]),
	.datac(!din_a[277]),
	.datad(!din_b[281]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_184 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[267]),
	.datac(!din_a[268]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_714 ),
	.cout(Xd_0__inst_mult_22_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_185 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[270]),
	.datac(!din_a[265]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_719 ),
	.cout(Xd_0__inst_mult_22_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_22_186 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[270]),
	.datac(!din_a[265]),
	.datad(!din_b[269]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_184 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[207]),
	.datac(!din_a[208]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_714 ),
	.cout(Xd_0__inst_mult_17_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_185 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[210]),
	.datac(!din_a[205]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_719 ),
	.cout(Xd_0__inst_mult_17_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_17_186 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[210]),
	.datac(!din_a[205]),
	.datad(!din_b[209]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_184 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[195]),
	.datac(!din_a[196]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_714 ),
	.cout(Xd_0__inst_mult_16_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_185 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[198]),
	.datac(!din_a[193]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_719 ),
	.cout(Xd_0__inst_mult_16_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_16_186 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[198]),
	.datac(!din_a[193]),
	.datad(!din_b[197]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_184 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[231]),
	.datac(!din_a[232]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_714 ),
	.cout(Xd_0__inst_mult_19_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_185 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[234]),
	.datac(!din_a[229]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_430 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_719 ),
	.cout(Xd_0__inst_mult_19_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_19_186 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[234]),
	.datac(!din_a[229]),
	.datad(!din_b[233]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_180 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[219]),
	.datac(!din_a[220]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_694 ),
	.cout(Xd_0__inst_mult_18_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_181 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[222]),
	.datac(!din_a[217]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_699 ),
	.cout(Xd_0__inst_mult_18_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_18_182 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[222]),
	.datac(!din_a[217]),
	.datad(!din_b[221]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_182 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[159]),
	.datac(!din_a[160]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_704 ),
	.cout(Xd_0__inst_mult_13_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_183 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[162]),
	.datac(!din_a[157]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_709 ),
	.cout(Xd_0__inst_mult_13_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_13_184 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[162]),
	.datac(!din_a[157]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_180 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[147]),
	.datac(!din_a[148]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_694 ),
	.cout(Xd_0__inst_mult_12_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_181 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[150]),
	.datac(!din_a[145]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_699 ),
	.cout(Xd_0__inst_mult_12_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_12_182 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[150]),
	.datac(!din_a[145]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_180 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[183]),
	.datac(!din_a[184]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_694 ),
	.cout(Xd_0__inst_mult_15_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_181 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[186]),
	.datac(!din_a[181]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_699 ),
	.cout(Xd_0__inst_mult_15_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_15_182 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[186]),
	.datac(!din_a[181]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_180 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[171]),
	.datac(!din_a[172]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_690 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_694 ),
	.cout(Xd_0__inst_mult_14_695 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_181 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[174]),
	.datac(!din_a[169]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_365 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_699 ),
	.cout(Xd_0__inst_mult_14_700 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_14_182 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[174]),
	.datac(!din_a[169]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_182 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[111]),
	.datac(!din_a[112]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_704 ),
	.cout(Xd_0__inst_mult_9_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_183 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[114]),
	.datac(!din_a[109]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_709 ),
	.cout(Xd_0__inst_mult_9_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_9_184 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[114]),
	.datac(!din_a[109]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_182 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[99]),
	.datac(!din_a[100]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_704 ),
	.cout(Xd_0__inst_mult_8_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_183 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[102]),
	.datac(!din_a[97]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_709 ),
	.cout(Xd_0__inst_mult_8_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_8_184 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[102]),
	.datac(!din_a[97]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_182 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[135]),
	.datac(!din_a[136]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_704 ),
	.cout(Xd_0__inst_mult_11_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_183 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[138]),
	.datac(!din_a[133]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_709 ),
	.cout(Xd_0__inst_mult_11_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_11_184 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[138]),
	.datac(!din_a[133]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_182 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[123]),
	.datac(!din_a[124]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_704 ),
	.cout(Xd_0__inst_mult_10_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_183 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[126]),
	.datac(!din_a[121]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_709 ),
	.cout(Xd_0__inst_mult_10_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_10_184 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[126]),
	.datac(!din_a[121]),
	.datad(!din_b[125]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_182 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[63]),
	.datac(!din_a[64]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_704 ),
	.cout(Xd_0__inst_mult_5_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_183 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[66]),
	.datac(!din_a[61]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_709 ),
	.cout(Xd_0__inst_mult_5_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_5_184 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[66]),
	.datac(!din_a[61]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_182 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[51]),
	.datac(!din_a[52]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_704 ),
	.cout(Xd_0__inst_mult_4_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_183 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[54]),
	.datac(!din_a[49]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_709 ),
	.cout(Xd_0__inst_mult_4_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_4_184 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[54]),
	.datac(!din_a[49]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_182 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[87]),
	.datac(!din_a[88]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_704 ),
	.cout(Xd_0__inst_mult_7_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_183 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[90]),
	.datac(!din_a[85]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_709 ),
	.cout(Xd_0__inst_mult_7_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_7_184 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[90]),
	.datac(!din_a[85]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_182 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[75]),
	.datac(!din_a[76]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_704 ),
	.cout(Xd_0__inst_mult_6_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_183 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[78]),
	.datac(!din_a[73]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_709 ),
	.cout(Xd_0__inst_mult_6_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_6_184 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[78]),
	.datac(!din_a[73]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_182 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[15]),
	.datac(!din_a[16]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_704 ),
	.cout(Xd_0__inst_mult_1_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_183 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[18]),
	.datac(!din_a[13]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_709 ),
	.cout(Xd_0__inst_mult_1_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_1_184 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[18]),
	.datac(!din_a[13]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_182 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[3]),
	.datac(!din_a[4]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_704 ),
	.cout(Xd_0__inst_mult_0_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_183 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[6]),
	.datac(!din_a[1]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_709 ),
	.cout(Xd_0__inst_mult_0_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_0_184 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[6]),
	.datac(!din_a[1]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_182 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[39]),
	.datac(!din_a[40]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_704 ),
	.cout(Xd_0__inst_mult_3_705 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_183 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[42]),
	.datac(!din_a[37]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_390 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_709 ),
	.cout(Xd_0__inst_mult_3_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_3_184 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[42]),
	.datac(!din_a[37]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_191 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[27]),
	.datac(!din_a[28]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_749 ),
	.cout(Xd_0__inst_mult_2_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_2_192 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[30]),
	.datac(!din_a[25]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(gnd),
	.sharein(),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_187 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[351]),
	.datac(!din_a[353]),
	.datad(!din_b[352]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_729 ),
	.cout(Xd_0__inst_mult_29_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_188 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[354]),
	.datac(!din_a[350]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_734 ),
	.cout(Xd_0__inst_mult_29_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_185 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[339]),
	.datac(!din_a[341]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_719 ),
	.cout(Xd_0__inst_mult_28_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_186 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[342]),
	.datac(!din_a[338]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_724 ),
	.cout(Xd_0__inst_mult_28_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_185 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[375]),
	.datac(!din_a[377]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_719 ),
	.cout(Xd_0__inst_mult_31_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_186 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[378]),
	.datac(!din_a[374]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_724 ),
	.cout(Xd_0__inst_mult_31_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_185 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[363]),
	.datac(!din_a[365]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_719 ),
	.cout(Xd_0__inst_mult_30_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_186 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[366]),
	.datac(!din_a[362]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_724 ),
	.cout(Xd_0__inst_mult_30_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_188 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[306]),
	.datac(!din_a[302]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_734 ),
	.cout(Xd_0__inst_mult_25_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_24_203 (
// Equation(s):

	.dataa(!din_a[291]),
	.datab(!din_b[294]),
	.datac(!din_a[290]),
	.datad(!din_b[295]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_24_800 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_24_809 ),
	.cout(Xd_0__inst_mult_24_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_188 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[330]),
	.datac(!din_a[326]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_734 ),
	.cout(Xd_0__inst_mult_27_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_26_203 (
// Equation(s):

	.dataa(!din_a[315]),
	.datab(!din_b[318]),
	.datac(!din_a[314]),
	.datad(!din_b[319]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_26_800 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_26_809 ),
	.cout(Xd_0__inst_mult_26_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_187 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[255]),
	.datac(!din_a[257]),
	.datad(!din_b[256]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_729 ),
	.cout(Xd_0__inst_mult_21_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_188 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[258]),
	.datac(!din_a[254]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_734 ),
	.cout(Xd_0__inst_mult_21_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_187 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[243]),
	.datac(!din_a[245]),
	.datad(!din_b[244]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_729 ),
	.cout(Xd_0__inst_mult_20_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_188 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[246]),
	.datac(!din_a[242]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_734 ),
	.cout(Xd_0__inst_mult_20_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_187 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[279]),
	.datac(!din_a[281]),
	.datad(!din_b[280]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_729 ),
	.cout(Xd_0__inst_mult_23_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_188 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[282]),
	.datac(!din_a[278]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_734 ),
	.cout(Xd_0__inst_mult_23_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_187 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[267]),
	.datac(!din_a[269]),
	.datad(!din_b[268]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_729 ),
	.cout(Xd_0__inst_mult_22_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_188 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[270]),
	.datac(!din_a[266]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_734 ),
	.cout(Xd_0__inst_mult_22_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_187 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[207]),
	.datac(!din_a[209]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_729 ),
	.cout(Xd_0__inst_mult_17_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_188 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[210]),
	.datac(!din_a[206]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_734 ),
	.cout(Xd_0__inst_mult_17_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_187 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[195]),
	.datac(!din_a[197]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_729 ),
	.cout(Xd_0__inst_mult_16_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_188 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[198]),
	.datac(!din_a[194]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_734 ),
	.cout(Xd_0__inst_mult_16_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_187 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[231]),
	.datac(!din_a[233]),
	.datad(!din_b[232]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_729 ),
	.cout(Xd_0__inst_mult_19_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_188 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[234]),
	.datac(!din_a[230]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_734 ),
	.cout(Xd_0__inst_mult_19_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_183 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[219]),
	.datac(!din_a[221]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_709 ),
	.cout(Xd_0__inst_mult_18_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_184 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[222]),
	.datac(!din_a[218]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_714 ),
	.cout(Xd_0__inst_mult_18_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_185 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[159]),
	.datac(!din_a[161]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_719 ),
	.cout(Xd_0__inst_mult_13_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_186 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[162]),
	.datac(!din_a[158]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_724 ),
	.cout(Xd_0__inst_mult_13_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_183 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[147]),
	.datac(!din_a[149]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_709 ),
	.cout(Xd_0__inst_mult_12_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_184 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[150]),
	.datac(!din_a[146]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_714 ),
	.cout(Xd_0__inst_mult_12_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_183 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[183]),
	.datac(!din_a[185]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_709 ),
	.cout(Xd_0__inst_mult_15_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_184 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[186]),
	.datac(!din_a[182]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_714 ),
	.cout(Xd_0__inst_mult_15_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_183 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[171]),
	.datac(!din_a[173]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_695 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_709 ),
	.cout(Xd_0__inst_mult_14_710 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_184 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[174]),
	.datac(!din_a[170]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_700 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_714 ),
	.cout(Xd_0__inst_mult_14_715 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_185 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[111]),
	.datac(!din_a[113]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_719 ),
	.cout(Xd_0__inst_mult_9_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_186 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[114]),
	.datac(!din_a[110]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_724 ),
	.cout(Xd_0__inst_mult_9_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_185 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[99]),
	.datac(!din_a[101]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_719 ),
	.cout(Xd_0__inst_mult_8_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_186 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[102]),
	.datac(!din_a[98]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_724 ),
	.cout(Xd_0__inst_mult_8_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_185 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[135]),
	.datac(!din_a[137]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_719 ),
	.cout(Xd_0__inst_mult_11_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_186 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[138]),
	.datac(!din_a[134]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_724 ),
	.cout(Xd_0__inst_mult_11_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_185 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[123]),
	.datac(!din_a[125]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_719 ),
	.cout(Xd_0__inst_mult_10_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_186 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[126]),
	.datac(!din_a[122]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_724 ),
	.cout(Xd_0__inst_mult_10_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_185 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[63]),
	.datac(!din_a[65]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_719 ),
	.cout(Xd_0__inst_mult_5_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_186 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[66]),
	.datac(!din_a[62]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_724 ),
	.cout(Xd_0__inst_mult_5_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_185 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[51]),
	.datac(!din_a[53]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_719 ),
	.cout(Xd_0__inst_mult_4_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_186 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[54]),
	.datac(!din_a[50]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_724 ),
	.cout(Xd_0__inst_mult_4_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_185 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[87]),
	.datac(!din_a[89]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_719 ),
	.cout(Xd_0__inst_mult_7_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_186 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[90]),
	.datac(!din_a[86]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_724 ),
	.cout(Xd_0__inst_mult_7_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_185 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[75]),
	.datac(!din_a[77]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_719 ),
	.cout(Xd_0__inst_mult_6_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_186 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[78]),
	.datac(!din_a[74]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_724 ),
	.cout(Xd_0__inst_mult_6_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_185 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[15]),
	.datac(!din_a[17]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_719 ),
	.cout(Xd_0__inst_mult_1_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_186 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[18]),
	.datac(!din_a[14]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_724 ),
	.cout(Xd_0__inst_mult_1_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_185 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[3]),
	.datac(!din_a[5]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_719 ),
	.cout(Xd_0__inst_mult_0_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_186 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[6]),
	.datac(!din_a[2]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_724 ),
	.cout(Xd_0__inst_mult_0_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_185 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[39]),
	.datac(!din_a[41]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_705 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_719 ),
	.cout(Xd_0__inst_mult_3_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_186 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[42]),
	.datac(!din_a[38]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_724 ),
	.cout(Xd_0__inst_mult_3_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_193 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[27]),
	.datac(!din_a[29]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_759 ),
	.cout(Xd_0__inst_mult_2_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_189 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[354]),
	.datac(!din_a[351]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_739 ),
	.cout(Xd_0__inst_mult_29_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_187 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[339]),
	.datac(!din_a[342]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_729 ),
	.cout(Xd_0__inst_mult_28_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_188 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[342]),
	.datac(!din_a[339]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_734 ),
	.cout(Xd_0__inst_mult_28_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_187 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[375]),
	.datac(!din_a[378]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_729 ),
	.cout(Xd_0__inst_mult_31_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_188 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[378]),
	.datac(!din_a[375]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_734 ),
	.cout(Xd_0__inst_mult_31_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_187 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[363]),
	.datac(!din_a[366]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_729 ),
	.cout(Xd_0__inst_mult_30_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_188 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[366]),
	.datac(!din_a[363]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_734 ),
	.cout(Xd_0__inst_mult_30_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_189 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[306]),
	.datac(!din_a[303]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_739 ),
	.cout(Xd_0__inst_mult_25_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_189 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[330]),
	.datac(!din_a[327]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_739 ),
	.cout(Xd_0__inst_mult_27_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_189 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[258]),
	.datac(!din_a[255]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_739 ),
	.cout(Xd_0__inst_mult_21_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_189 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[246]),
	.datac(!din_a[243]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_739 ),
	.cout(Xd_0__inst_mult_20_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_189 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[282]),
	.datac(!din_a[279]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_739 ),
	.cout(Xd_0__inst_mult_23_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_189 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[270]),
	.datac(!din_a[267]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_739 ),
	.cout(Xd_0__inst_mult_22_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_189 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[210]),
	.datac(!din_a[207]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_739 ),
	.cout(Xd_0__inst_mult_17_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_189 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[198]),
	.datac(!din_a[195]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_739 ),
	.cout(Xd_0__inst_mult_16_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_189 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[234]),
	.datac(!din_a[231]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_739 ),
	.cout(Xd_0__inst_mult_19_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_185 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[219]),
	.datac(!din_a[222]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_719 ),
	.cout(Xd_0__inst_mult_18_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_186 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[222]),
	.datac(!din_a[219]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_724 ),
	.cout(Xd_0__inst_mult_18_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_187 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[159]),
	.datac(!din_a[162]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_729 ),
	.cout(Xd_0__inst_mult_13_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_188 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[162]),
	.datac(!din_a[159]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_734 ),
	.cout(Xd_0__inst_mult_13_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_185 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[147]),
	.datac(!din_a[150]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_719 ),
	.cout(Xd_0__inst_mult_12_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_186 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[150]),
	.datac(!din_a[147]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_724 ),
	.cout(Xd_0__inst_mult_12_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_185 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[183]),
	.datac(!din_a[186]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_719 ),
	.cout(Xd_0__inst_mult_15_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_186 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[186]),
	.datac(!din_a[183]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_724 ),
	.cout(Xd_0__inst_mult_15_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_185 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[171]),
	.datac(!din_a[174]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_710 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_719 ),
	.cout(Xd_0__inst_mult_14_720 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_186 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[174]),
	.datac(!din_a[171]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_715 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_724 ),
	.cout(Xd_0__inst_mult_14_725 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_187 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[111]),
	.datac(!din_a[114]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_729 ),
	.cout(Xd_0__inst_mult_9_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_188 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[114]),
	.datac(!din_a[111]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_734 ),
	.cout(Xd_0__inst_mult_9_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_187 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[99]),
	.datac(!din_a[102]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_729 ),
	.cout(Xd_0__inst_mult_8_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_188 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[102]),
	.datac(!din_a[99]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_734 ),
	.cout(Xd_0__inst_mult_8_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_187 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[135]),
	.datac(!din_a[138]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_729 ),
	.cout(Xd_0__inst_mult_11_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_188 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[138]),
	.datac(!din_a[135]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_734 ),
	.cout(Xd_0__inst_mult_11_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_187 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[123]),
	.datac(!din_a[126]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_729 ),
	.cout(Xd_0__inst_mult_10_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_188 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[126]),
	.datac(!din_a[123]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_734 ),
	.cout(Xd_0__inst_mult_10_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_187 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[63]),
	.datac(!din_a[66]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_729 ),
	.cout(Xd_0__inst_mult_5_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_188 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[66]),
	.datac(!din_a[63]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_734 ),
	.cout(Xd_0__inst_mult_5_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_187 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[51]),
	.datac(!din_a[54]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_729 ),
	.cout(Xd_0__inst_mult_4_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_188 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[54]),
	.datac(!din_a[51]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_734 ),
	.cout(Xd_0__inst_mult_4_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_187 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[87]),
	.datac(!din_a[90]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_729 ),
	.cout(Xd_0__inst_mult_7_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_188 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[90]),
	.datac(!din_a[87]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_734 ),
	.cout(Xd_0__inst_mult_7_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_187 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[75]),
	.datac(!din_a[78]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_729 ),
	.cout(Xd_0__inst_mult_6_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_188 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[78]),
	.datac(!din_a[75]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_734 ),
	.cout(Xd_0__inst_mult_6_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_187 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[15]),
	.datac(!din_a[18]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_729 ),
	.cout(Xd_0__inst_mult_1_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_188 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[18]),
	.datac(!din_a[15]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_734 ),
	.cout(Xd_0__inst_mult_1_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_187 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[3]),
	.datac(!din_a[6]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_729 ),
	.cout(Xd_0__inst_mult_0_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_188 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[6]),
	.datac(!din_a[3]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_734 ),
	.cout(Xd_0__inst_mult_0_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_187 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[39]),
	.datac(!din_a[42]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_729 ),
	.cout(Xd_0__inst_mult_3_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_188 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[42]),
	.datac(!din_a[39]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_734 ),
	.cout(Xd_0__inst_mult_3_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_194 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[27]),
	.datac(!din_a[30]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_764 ),
	.cout(Xd_0__inst_mult_2_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_190 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[354]),
	.datac(!din_a[352]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_744 ),
	.cout(Xd_0__inst_mult_29_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_191 (
// Equation(s):

	.dataa(!din_a[350]),
	.datab(!din_b[357]),
	.datac(!din_a[349]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_749 ),
	.cout(Xd_0__inst_mult_29_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_29_192 (
// Equation(s):

	.dataa(!din_a[348]),
	.datab(!din_b[357]),
	.datac(!din_a[349]),
	.datad(!din_b[356]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_754 ),
	.cout(Xd_0__inst_mult_29_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_189 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[339]),
	.datac(!din_a[343]),
	.datad(!din_b[340]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_739 ),
	.cout(Xd_0__inst_mult_28_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_190 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[342]),
	.datac(!din_a[340]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_744 ),
	.cout(Xd_0__inst_mult_28_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_191 (
// Equation(s):

	.dataa(!din_a[338]),
	.datab(!din_b[345]),
	.datac(!din_a[337]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_749 ),
	.cout(Xd_0__inst_mult_28_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_28_192 (
// Equation(s):

	.dataa(!din_a[336]),
	.datab(!din_b[345]),
	.datac(!din_a[337]),
	.datad(!din_b[344]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_754 ),
	.cout(Xd_0__inst_mult_28_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_189 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[375]),
	.datac(!din_a[379]),
	.datad(!din_b[376]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_739 ),
	.cout(Xd_0__inst_mult_31_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_190 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[378]),
	.datac(!din_a[376]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_744 ),
	.cout(Xd_0__inst_mult_31_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_191 (
// Equation(s):

	.dataa(!din_a[374]),
	.datab(!din_b[381]),
	.datac(!din_a[373]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_749 ),
	.cout(Xd_0__inst_mult_31_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_31_192 (
// Equation(s):

	.dataa(!din_a[372]),
	.datab(!din_b[381]),
	.datac(!din_a[373]),
	.datad(!din_b[380]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_754 ),
	.cout(Xd_0__inst_mult_31_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_189 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[363]),
	.datac(!din_a[367]),
	.datad(!din_b[364]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_739 ),
	.cout(Xd_0__inst_mult_30_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_190 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[366]),
	.datac(!din_a[364]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_744 ),
	.cout(Xd_0__inst_mult_30_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_191 (
// Equation(s):

	.dataa(!din_a[362]),
	.datab(!din_b[369]),
	.datac(!din_a[361]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_749 ),
	.cout(Xd_0__inst_mult_30_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_30_192 (
// Equation(s):

	.dataa(!din_a[360]),
	.datab(!din_b[369]),
	.datac(!din_a[361]),
	.datad(!din_b[368]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_754 ),
	.cout(Xd_0__inst_mult_30_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_190 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[306]),
	.datac(!din_a[304]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_744 ),
	.cout(Xd_0__inst_mult_25_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_191 (
// Equation(s):

	.dataa(!din_a[302]),
	.datab(!din_b[309]),
	.datac(!din_a[301]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_749 ),
	.cout(Xd_0__inst_mult_25_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_25_192 (
// Equation(s):

	.dataa(!din_a[300]),
	.datab(!din_b[309]),
	.datac(!din_a[301]),
	.datad(!din_b[308]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_754 ),
	.cout(Xd_0__inst_mult_25_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_190 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[330]),
	.datac(!din_a[328]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_744 ),
	.cout(Xd_0__inst_mult_27_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_191 (
// Equation(s):

	.dataa(!din_a[326]),
	.datab(!din_b[333]),
	.datac(!din_a[325]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_620 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_749 ),
	.cout(Xd_0__inst_mult_27_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_27_192 (
// Equation(s):

	.dataa(!din_a[324]),
	.datab(!din_b[333]),
	.datac(!din_a[325]),
	.datad(!din_b[332]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_754 ),
	.cout(Xd_0__inst_mult_27_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_190 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[258]),
	.datac(!din_a[256]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_744 ),
	.cout(Xd_0__inst_mult_21_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_191 (
// Equation(s):

	.dataa(!din_a[254]),
	.datab(!din_b[261]),
	.datac(!din_a[253]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_749 ),
	.cout(Xd_0__inst_mult_21_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_21_192 (
// Equation(s):

	.dataa(!din_a[252]),
	.datab(!din_b[261]),
	.datac(!din_a[253]),
	.datad(!din_b[260]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_754 ),
	.cout(Xd_0__inst_mult_21_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_190 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[246]),
	.datac(!din_a[244]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_744 ),
	.cout(Xd_0__inst_mult_20_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_191 (
// Equation(s):

	.dataa(!din_a[242]),
	.datab(!din_b[249]),
	.datac(!din_a[241]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_749 ),
	.cout(Xd_0__inst_mult_20_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_20_192 (
// Equation(s):

	.dataa(!din_a[240]),
	.datab(!din_b[249]),
	.datac(!din_a[241]),
	.datad(!din_b[248]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_754 ),
	.cout(Xd_0__inst_mult_20_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_190 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[282]),
	.datac(!din_a[280]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_744 ),
	.cout(Xd_0__inst_mult_23_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_191 (
// Equation(s):

	.dataa(!din_a[278]),
	.datab(!din_b[285]),
	.datac(!din_a[277]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_749 ),
	.cout(Xd_0__inst_mult_23_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_23_192 (
// Equation(s):

	.dataa(!din_a[276]),
	.datab(!din_b[285]),
	.datac(!din_a[277]),
	.datad(!din_b[284]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_754 ),
	.cout(Xd_0__inst_mult_23_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_190 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[270]),
	.datac(!din_a[268]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_744 ),
	.cout(Xd_0__inst_mult_22_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_191 (
// Equation(s):

	.dataa(!din_a[266]),
	.datab(!din_b[273]),
	.datac(!din_a[265]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_749 ),
	.cout(Xd_0__inst_mult_22_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_22_192 (
// Equation(s):

	.dataa(!din_a[264]),
	.datab(!din_b[273]),
	.datac(!din_a[265]),
	.datad(!din_b[272]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_754 ),
	.cout(Xd_0__inst_mult_22_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_190 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[210]),
	.datac(!din_a[208]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_744 ),
	.cout(Xd_0__inst_mult_17_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_191 (
// Equation(s):

	.dataa(!din_a[206]),
	.datab(!din_b[213]),
	.datac(!din_a[205]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_749 ),
	.cout(Xd_0__inst_mult_17_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_17_192 (
// Equation(s):

	.dataa(!din_a[204]),
	.datab(!din_b[213]),
	.datac(!din_a[205]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_754 ),
	.cout(Xd_0__inst_mult_17_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_190 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[198]),
	.datac(!din_a[196]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_744 ),
	.cout(Xd_0__inst_mult_16_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_191 (
// Equation(s):

	.dataa(!din_a[194]),
	.datab(!din_b[201]),
	.datac(!din_a[193]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_749 ),
	.cout(Xd_0__inst_mult_16_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_16_192 (
// Equation(s):

	.dataa(!din_a[192]),
	.datab(!din_b[201]),
	.datac(!din_a[193]),
	.datad(!din_b[200]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_754 ),
	.cout(Xd_0__inst_mult_16_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_190 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[234]),
	.datac(!din_a[232]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_744 ),
	.cout(Xd_0__inst_mult_19_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_191 (
// Equation(s):

	.dataa(!din_a[230]),
	.datab(!din_b[237]),
	.datac(!din_a[229]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_605 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_749 ),
	.cout(Xd_0__inst_mult_19_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_19_192 (
// Equation(s):

	.dataa(!din_a[228]),
	.datab(!din_b[237]),
	.datac(!din_a[229]),
	.datad(!din_b[236]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_754 ),
	.cout(Xd_0__inst_mult_19_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_187 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[219]),
	.datac(!din_a[223]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_729 ),
	.cout(Xd_0__inst_mult_18_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_188 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[222]),
	.datac(!din_a[220]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_734 ),
	.cout(Xd_0__inst_mult_18_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_189 (
// Equation(s):

	.dataa(!din_a[218]),
	.datab(!din_b[225]),
	.datac(!din_a[217]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_739 ),
	.cout(Xd_0__inst_mult_18_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_18_190 (
// Equation(s):

	.dataa(!din_a[216]),
	.datab(!din_b[225]),
	.datac(!din_a[217]),
	.datad(!din_b[224]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_744 ),
	.cout(Xd_0__inst_mult_18_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_189 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[159]),
	.datac(!din_a[163]),
	.datad(!din_b[160]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_739 ),
	.cout(Xd_0__inst_mult_13_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_190 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[162]),
	.datac(!din_a[160]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_744 ),
	.cout(Xd_0__inst_mult_13_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_191 (
// Equation(s):

	.dataa(!din_a[158]),
	.datab(!din_b[165]),
	.datac(!din_a[157]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_749 ),
	.cout(Xd_0__inst_mult_13_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_13_192 (
// Equation(s):

	.dataa(!din_a[156]),
	.datab(!din_b[165]),
	.datac(!din_a[157]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_754 ),
	.cout(Xd_0__inst_mult_13_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_187 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[147]),
	.datac(!din_a[151]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_729 ),
	.cout(Xd_0__inst_mult_12_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_188 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[150]),
	.datac(!din_a[148]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_734 ),
	.cout(Xd_0__inst_mult_12_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_189 (
// Equation(s):

	.dataa(!din_a[146]),
	.datab(!din_b[153]),
	.datac(!din_a[145]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_739 ),
	.cout(Xd_0__inst_mult_12_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_12_190 (
// Equation(s):

	.dataa(!din_a[144]),
	.datab(!din_b[153]),
	.datac(!din_a[145]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_744 ),
	.cout(Xd_0__inst_mult_12_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_187 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[183]),
	.datac(!din_a[187]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_729 ),
	.cout(Xd_0__inst_mult_15_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_188 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[186]),
	.datac(!din_a[184]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_734 ),
	.cout(Xd_0__inst_mult_15_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_189 (
// Equation(s):

	.dataa(!din_a[182]),
	.datab(!din_b[189]),
	.datac(!din_a[181]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_739 ),
	.cout(Xd_0__inst_mult_15_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_15_190 (
// Equation(s):

	.dataa(!din_a[180]),
	.datab(!din_b[189]),
	.datac(!din_a[181]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_744 ),
	.cout(Xd_0__inst_mult_15_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_187 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[171]),
	.datac(!din_a[175]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_720 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_729 ),
	.cout(Xd_0__inst_mult_14_730 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_188 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[174]),
	.datac(!din_a[172]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_725 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_734 ),
	.cout(Xd_0__inst_mult_14_735 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_189 (
// Equation(s):

	.dataa(!din_a[170]),
	.datab(!din_b[177]),
	.datac(!din_a[169]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_560 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_739 ),
	.cout(Xd_0__inst_mult_14_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_14_190 (
// Equation(s):

	.dataa(!din_a[168]),
	.datab(!din_b[177]),
	.datac(!din_a[169]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_744 ),
	.cout(Xd_0__inst_mult_14_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_189 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[111]),
	.datac(!din_a[115]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_739 ),
	.cout(Xd_0__inst_mult_9_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_190 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[114]),
	.datac(!din_a[112]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_744 ),
	.cout(Xd_0__inst_mult_9_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_191 (
// Equation(s):

	.dataa(!din_a[110]),
	.datab(!din_b[117]),
	.datac(!din_a[109]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_749 ),
	.cout(Xd_0__inst_mult_9_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_9_192 (
// Equation(s):

	.dataa(!din_a[108]),
	.datab(!din_b[117]),
	.datac(!din_a[109]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_754 ),
	.cout(Xd_0__inst_mult_9_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_189 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[99]),
	.datac(!din_a[103]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_739 ),
	.cout(Xd_0__inst_mult_8_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_190 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[102]),
	.datac(!din_a[100]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_744 ),
	.cout(Xd_0__inst_mult_8_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_191 (
// Equation(s):

	.dataa(!din_a[98]),
	.datab(!din_b[105]),
	.datac(!din_a[97]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_749 ),
	.cout(Xd_0__inst_mult_8_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_8_192 (
// Equation(s):

	.dataa(!din_a[96]),
	.datab(!din_b[105]),
	.datac(!din_a[97]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_754 ),
	.cout(Xd_0__inst_mult_8_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_189 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[135]),
	.datac(!din_a[139]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_739 ),
	.cout(Xd_0__inst_mult_11_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_190 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[138]),
	.datac(!din_a[136]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_744 ),
	.cout(Xd_0__inst_mult_11_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_191 (
// Equation(s):

	.dataa(!din_a[134]),
	.datab(!din_b[141]),
	.datac(!din_a[133]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_749 ),
	.cout(Xd_0__inst_mult_11_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_11_192 (
// Equation(s):

	.dataa(!din_a[132]),
	.datab(!din_b[141]),
	.datac(!din_a[133]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_754 ),
	.cout(Xd_0__inst_mult_11_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_189 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[123]),
	.datac(!din_a[127]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_739 ),
	.cout(Xd_0__inst_mult_10_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_190 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[126]),
	.datac(!din_a[124]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_744 ),
	.cout(Xd_0__inst_mult_10_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_191 (
// Equation(s):

	.dataa(!din_a[122]),
	.datab(!din_b[129]),
	.datac(!din_a[121]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_749 ),
	.cout(Xd_0__inst_mult_10_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_10_192 (
// Equation(s):

	.dataa(!din_a[120]),
	.datab(!din_b[129]),
	.datac(!din_a[121]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_754 ),
	.cout(Xd_0__inst_mult_10_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_189 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[63]),
	.datac(!din_a[67]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_739 ),
	.cout(Xd_0__inst_mult_5_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_190 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[66]),
	.datac(!din_a[64]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_744 ),
	.cout(Xd_0__inst_mult_5_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_191 (
// Equation(s):

	.dataa(!din_a[62]),
	.datab(!din_b[69]),
	.datac(!din_a[61]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_749 ),
	.cout(Xd_0__inst_mult_5_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_5_192 (
// Equation(s):

	.dataa(!din_a[60]),
	.datab(!din_b[69]),
	.datac(!din_a[61]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_754 ),
	.cout(Xd_0__inst_mult_5_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_189 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[51]),
	.datac(!din_a[55]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_739 ),
	.cout(Xd_0__inst_mult_4_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_190 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[54]),
	.datac(!din_a[52]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_744 ),
	.cout(Xd_0__inst_mult_4_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_191 (
// Equation(s):

	.dataa(!din_a[50]),
	.datab(!din_b[57]),
	.datac(!din_a[49]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_749 ),
	.cout(Xd_0__inst_mult_4_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_4_192 (
// Equation(s):

	.dataa(!din_a[48]),
	.datab(!din_b[57]),
	.datac(!din_a[49]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_754 ),
	.cout(Xd_0__inst_mult_4_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_189 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[87]),
	.datac(!din_a[91]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_739 ),
	.cout(Xd_0__inst_mult_7_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_190 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[90]),
	.datac(!din_a[88]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_744 ),
	.cout(Xd_0__inst_mult_7_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_191 (
// Equation(s):

	.dataa(!din_a[86]),
	.datab(!din_b[93]),
	.datac(!din_a[85]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_749 ),
	.cout(Xd_0__inst_mult_7_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_7_192 (
// Equation(s):

	.dataa(!din_a[84]),
	.datab(!din_b[93]),
	.datac(!din_a[85]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_754 ),
	.cout(Xd_0__inst_mult_7_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_189 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[75]),
	.datac(!din_a[79]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_739 ),
	.cout(Xd_0__inst_mult_6_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_190 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[78]),
	.datac(!din_a[76]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_744 ),
	.cout(Xd_0__inst_mult_6_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_191 (
// Equation(s):

	.dataa(!din_a[74]),
	.datab(!din_b[81]),
	.datac(!din_a[73]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_749 ),
	.cout(Xd_0__inst_mult_6_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_6_192 (
// Equation(s):

	.dataa(!din_a[72]),
	.datab(!din_b[81]),
	.datac(!din_a[73]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_754 ),
	.cout(Xd_0__inst_mult_6_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_189 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[15]),
	.datac(!din_a[19]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_739 ),
	.cout(Xd_0__inst_mult_1_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_190 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[18]),
	.datac(!din_a[16]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_744 ),
	.cout(Xd_0__inst_mult_1_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_191 (
// Equation(s):

	.dataa(!din_a[14]),
	.datab(!din_b[21]),
	.datac(!din_a[13]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_749 ),
	.cout(Xd_0__inst_mult_1_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_1_192 (
// Equation(s):

	.dataa(!din_a[12]),
	.datab(!din_b[21]),
	.datac(!din_a[13]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_754 ),
	.cout(Xd_0__inst_mult_1_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_189 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[3]),
	.datac(!din_a[7]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_739 ),
	.cout(Xd_0__inst_mult_0_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_190 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[6]),
	.datac(!din_a[4]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_744 ),
	.cout(Xd_0__inst_mult_0_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_191 (
// Equation(s):

	.dataa(!din_a[2]),
	.datab(!din_b[9]),
	.datac(!din_a[1]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_749 ),
	.cout(Xd_0__inst_mult_0_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_0_192 (
// Equation(s):

	.dataa(!din_a[0]),
	.datab(!din_b[9]),
	.datac(!din_a[1]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_754 ),
	.cout(Xd_0__inst_mult_0_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_189 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[39]),
	.datac(!din_a[43]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_739 ),
	.cout(Xd_0__inst_mult_3_740 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_190 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[42]),
	.datac(!din_a[40]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_744 ),
	.cout(Xd_0__inst_mult_3_745 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_191 (
// Equation(s):

	.dataa(!din_a[38]),
	.datab(!din_b[45]),
	.datac(!din_a[37]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_585 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_749 ),
	.cout(Xd_0__inst_mult_3_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_3_192 (
// Equation(s):

	.dataa(!din_a[36]),
	.datab(!din_b[45]),
	.datac(!din_a[37]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_754 ),
	.cout(Xd_0__inst_mult_3_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_195 (
// Equation(s):

	.dataa(!din_a[32]),
	.datab(!din_b[27]),
	.datac(!din_a[31]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_769 ),
	.cout(Xd_0__inst_mult_2_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_196 (
// Equation(s):

	.dataa(!din_a[26]),
	.datab(!din_b[33]),
	.datac(!din_a[25]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_630 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_774 ),
	.cout(Xd_0__inst_mult_2_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000010000),
	.shared_arith("off")
) Xd_0__inst_mult_2_197 (
// Equation(s):

	.dataa(!din_a[24]),
	.datab(!din_b[33]),
	.datac(!din_a[25]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_810 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_779 ),
	.cout(Xd_0__inst_mult_2_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_193 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[354]),
	.datac(!din_a[353]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_759 ),
	.cout(Xd_0__inst_mult_29_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_194 (
// Equation(s):

	.dataa(!din_a[351]),
	.datab(!din_b[357]),
	.datac(!din_a[350]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_764 ),
	.cout(Xd_0__inst_mult_29_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_193 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[342]),
	.datac(!din_a[341]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_759 ),
	.cout(Xd_0__inst_mult_28_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_194 (
// Equation(s):

	.dataa(!din_a[339]),
	.datab(!din_b[345]),
	.datac(!din_a[338]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_764 ),
	.cout(Xd_0__inst_mult_28_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_193 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[378]),
	.datac(!din_a[377]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_759 ),
	.cout(Xd_0__inst_mult_31_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_194 (
// Equation(s):

	.dataa(!din_a[375]),
	.datab(!din_b[381]),
	.datac(!din_a[374]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_764 ),
	.cout(Xd_0__inst_mult_31_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_193 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[366]),
	.datac(!din_a[365]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_759 ),
	.cout(Xd_0__inst_mult_30_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_194 (
// Equation(s):

	.dataa(!din_a[363]),
	.datab(!din_b[369]),
	.datac(!din_a[362]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_764 ),
	.cout(Xd_0__inst_mult_30_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_193 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[306]),
	.datac(!din_a[305]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_759 ),
	.cout(Xd_0__inst_mult_25_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_194 (
// Equation(s):

	.dataa(!din_a[303]),
	.datab(!din_b[309]),
	.datac(!din_a[302]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_764 ),
	.cout(Xd_0__inst_mult_25_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_193 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[330]),
	.datac(!din_a[329]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_759 ),
	.cout(Xd_0__inst_mult_27_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_194 (
// Equation(s):

	.dataa(!din_a[327]),
	.datab(!din_b[333]),
	.datac(!din_a[326]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_764 ),
	.cout(Xd_0__inst_mult_27_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_193 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[258]),
	.datac(!din_a[257]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_759 ),
	.cout(Xd_0__inst_mult_21_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_194 (
// Equation(s):

	.dataa(!din_a[255]),
	.datab(!din_b[261]),
	.datac(!din_a[254]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_764 ),
	.cout(Xd_0__inst_mult_21_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_193 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[246]),
	.datac(!din_a[245]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_759 ),
	.cout(Xd_0__inst_mult_20_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_194 (
// Equation(s):

	.dataa(!din_a[243]),
	.datab(!din_b[249]),
	.datac(!din_a[242]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_764 ),
	.cout(Xd_0__inst_mult_20_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_193 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[282]),
	.datac(!din_a[281]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_759 ),
	.cout(Xd_0__inst_mult_23_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_194 (
// Equation(s):

	.dataa(!din_a[279]),
	.datab(!din_b[285]),
	.datac(!din_a[278]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_764 ),
	.cout(Xd_0__inst_mult_23_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_193 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[270]),
	.datac(!din_a[269]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_759 ),
	.cout(Xd_0__inst_mult_22_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_194 (
// Equation(s):

	.dataa(!din_a[267]),
	.datab(!din_b[273]),
	.datac(!din_a[266]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_764 ),
	.cout(Xd_0__inst_mult_22_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_193 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[210]),
	.datac(!din_a[209]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_759 ),
	.cout(Xd_0__inst_mult_17_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_194 (
// Equation(s):

	.dataa(!din_a[207]),
	.datab(!din_b[213]),
	.datac(!din_a[206]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_764 ),
	.cout(Xd_0__inst_mult_17_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_193 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[198]),
	.datac(!din_a[197]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_759 ),
	.cout(Xd_0__inst_mult_16_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_194 (
// Equation(s):

	.dataa(!din_a[195]),
	.datab(!din_b[201]),
	.datac(!din_a[194]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_764 ),
	.cout(Xd_0__inst_mult_16_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_193 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[234]),
	.datac(!din_a[233]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_759 ),
	.cout(Xd_0__inst_mult_19_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_194 (
// Equation(s):

	.dataa(!din_a[231]),
	.datab(!din_b[237]),
	.datac(!din_a[230]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_764 ),
	.cout(Xd_0__inst_mult_19_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_191 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[220]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_749 ),
	.cout(Xd_0__inst_mult_18_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_192 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[222]),
	.datac(!din_a[221]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_754 ),
	.cout(Xd_0__inst_mult_18_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_193 (
// Equation(s):

	.dataa(!din_a[219]),
	.datab(!din_b[225]),
	.datac(!din_a[218]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_759 ),
	.cout(Xd_0__inst_mult_18_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_193 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[162]),
	.datac(!din_a[161]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_759 ),
	.cout(Xd_0__inst_mult_13_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_194 (
// Equation(s):

	.dataa(!din_a[159]),
	.datab(!din_b[165]),
	.datac(!din_a[158]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_764 ),
	.cout(Xd_0__inst_mult_13_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_191 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[148]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_749 ),
	.cout(Xd_0__inst_mult_12_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_192 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[150]),
	.datac(!din_a[149]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_754 ),
	.cout(Xd_0__inst_mult_12_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_193 (
// Equation(s):

	.dataa(!din_a[147]),
	.datab(!din_b[153]),
	.datac(!din_a[146]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_759 ),
	.cout(Xd_0__inst_mult_12_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_191 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[184]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_749 ),
	.cout(Xd_0__inst_mult_15_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_192 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[186]),
	.datac(!din_a[185]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_754 ),
	.cout(Xd_0__inst_mult_15_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_193 (
// Equation(s):

	.dataa(!din_a[183]),
	.datab(!din_b[189]),
	.datac(!din_a[182]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_759 ),
	.cout(Xd_0__inst_mult_15_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_191 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[172]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_730 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_749 ),
	.cout(Xd_0__inst_mult_14_750 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_192 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[174]),
	.datac(!din_a[173]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_735 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_754 ),
	.cout(Xd_0__inst_mult_14_755 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_193 (
// Equation(s):

	.dataa(!din_a[171]),
	.datab(!din_b[177]),
	.datac(!din_a[170]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_740 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_759 ),
	.cout(Xd_0__inst_mult_14_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_193 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[114]),
	.datac(!din_a[113]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_759 ),
	.cout(Xd_0__inst_mult_9_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_194 (
// Equation(s):

	.dataa(!din_a[111]),
	.datab(!din_b[117]),
	.datac(!din_a[110]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_764 ),
	.cout(Xd_0__inst_mult_9_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_193 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[102]),
	.datac(!din_a[101]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_759 ),
	.cout(Xd_0__inst_mult_8_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_194 (
// Equation(s):

	.dataa(!din_a[99]),
	.datab(!din_b[105]),
	.datac(!din_a[98]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_764 ),
	.cout(Xd_0__inst_mult_8_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_193 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[138]),
	.datac(!din_a[137]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_759 ),
	.cout(Xd_0__inst_mult_11_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_194 (
// Equation(s):

	.dataa(!din_a[135]),
	.datab(!din_b[141]),
	.datac(!din_a[134]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_764 ),
	.cout(Xd_0__inst_mult_11_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_193 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[126]),
	.datac(!din_a[125]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_759 ),
	.cout(Xd_0__inst_mult_10_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_194 (
// Equation(s):

	.dataa(!din_a[123]),
	.datab(!din_b[129]),
	.datac(!din_a[122]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_764 ),
	.cout(Xd_0__inst_mult_10_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_193 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[66]),
	.datac(!din_a[65]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_759 ),
	.cout(Xd_0__inst_mult_5_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_194 (
// Equation(s):

	.dataa(!din_a[63]),
	.datab(!din_b[69]),
	.datac(!din_a[62]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_764 ),
	.cout(Xd_0__inst_mult_5_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_193 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[54]),
	.datac(!din_a[53]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_759 ),
	.cout(Xd_0__inst_mult_4_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_194 (
// Equation(s):

	.dataa(!din_a[51]),
	.datab(!din_b[57]),
	.datac(!din_a[50]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_764 ),
	.cout(Xd_0__inst_mult_4_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_193 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[90]),
	.datac(!din_a[89]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_759 ),
	.cout(Xd_0__inst_mult_7_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_194 (
// Equation(s):

	.dataa(!din_a[87]),
	.datab(!din_b[93]),
	.datac(!din_a[86]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_764 ),
	.cout(Xd_0__inst_mult_7_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_193 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[78]),
	.datac(!din_a[77]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_759 ),
	.cout(Xd_0__inst_mult_6_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_194 (
// Equation(s):

	.dataa(!din_a[75]),
	.datab(!din_b[81]),
	.datac(!din_a[74]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_764 ),
	.cout(Xd_0__inst_mult_6_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_193 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[18]),
	.datac(!din_a[17]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_759 ),
	.cout(Xd_0__inst_mult_1_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_194 (
// Equation(s):

	.dataa(!din_a[15]),
	.datab(!din_b[21]),
	.datac(!din_a[14]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_764 ),
	.cout(Xd_0__inst_mult_1_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_193 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[6]),
	.datac(!din_a[5]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_759 ),
	.cout(Xd_0__inst_mult_0_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_194 (
// Equation(s):

	.dataa(!din_a[3]),
	.datab(!din_b[9]),
	.datac(!din_a[2]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_764 ),
	.cout(Xd_0__inst_mult_0_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_193 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[42]),
	.datac(!din_a[41]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_745 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_759 ),
	.cout(Xd_0__inst_mult_3_760 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_194 (
// Equation(s):

	.dataa(!din_a[39]),
	.datab(!din_b[45]),
	.datac(!din_a[38]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_764 ),
	.cout(Xd_0__inst_mult_3_765 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_198 (
// Equation(s):

	.dataa(!din_a[27]),
	.datab(!din_b[33]),
	.datac(!din_a[26]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_784 ),
	.cout(Xd_0__inst_mult_2_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_195 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[354]),
	.datac(!din_a[354]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_769 ),
	.cout(Xd_0__inst_mult_29_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_196 (
// Equation(s):

	.dataa(!din_a[352]),
	.datab(!din_b[357]),
	.datac(!din_a[351]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_774 ),
	.cout(Xd_0__inst_mult_29_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_195 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[342]),
	.datac(!din_a[342]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_769 ),
	.cout(Xd_0__inst_mult_28_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_196 (
// Equation(s):

	.dataa(!din_a[340]),
	.datab(!din_b[345]),
	.datac(!din_a[339]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_774 ),
	.cout(Xd_0__inst_mult_28_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_195 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[378]),
	.datac(!din_a[378]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_769 ),
	.cout(Xd_0__inst_mult_31_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_196 (
// Equation(s):

	.dataa(!din_a[376]),
	.datab(!din_b[381]),
	.datac(!din_a[375]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_774 ),
	.cout(Xd_0__inst_mult_31_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_195 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[366]),
	.datac(!din_a[366]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_769 ),
	.cout(Xd_0__inst_mult_30_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_196 (
// Equation(s):

	.dataa(!din_a[364]),
	.datab(!din_b[369]),
	.datac(!din_a[363]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_774 ),
	.cout(Xd_0__inst_mult_30_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_195 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[306]),
	.datac(!din_a[306]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_769 ),
	.cout(Xd_0__inst_mult_25_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_196 (
// Equation(s):

	.dataa(!din_a[304]),
	.datab(!din_b[309]),
	.datac(!din_a[303]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_774 ),
	.cout(Xd_0__inst_mult_25_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_195 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[330]),
	.datac(!din_a[330]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_769 ),
	.cout(Xd_0__inst_mult_27_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_196 (
// Equation(s):

	.dataa(!din_a[328]),
	.datab(!din_b[333]),
	.datac(!din_a[327]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_774 ),
	.cout(Xd_0__inst_mult_27_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_195 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[258]),
	.datac(!din_a[258]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_769 ),
	.cout(Xd_0__inst_mult_21_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_196 (
// Equation(s):

	.dataa(!din_a[256]),
	.datab(!din_b[261]),
	.datac(!din_a[255]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_774 ),
	.cout(Xd_0__inst_mult_21_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_195 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[246]),
	.datac(!din_a[246]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_769 ),
	.cout(Xd_0__inst_mult_20_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_196 (
// Equation(s):

	.dataa(!din_a[244]),
	.datab(!din_b[249]),
	.datac(!din_a[243]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_774 ),
	.cout(Xd_0__inst_mult_20_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_195 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[282]),
	.datac(!din_a[282]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_769 ),
	.cout(Xd_0__inst_mult_23_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_196 (
// Equation(s):

	.dataa(!din_a[280]),
	.datab(!din_b[285]),
	.datac(!din_a[279]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_774 ),
	.cout(Xd_0__inst_mult_23_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_195 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[270]),
	.datac(!din_a[270]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_769 ),
	.cout(Xd_0__inst_mult_22_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_196 (
// Equation(s):

	.dataa(!din_a[268]),
	.datab(!din_b[273]),
	.datac(!din_a[267]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_774 ),
	.cout(Xd_0__inst_mult_22_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_195 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[210]),
	.datac(!din_a[210]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_769 ),
	.cout(Xd_0__inst_mult_17_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_196 (
// Equation(s):

	.dataa(!din_a[208]),
	.datab(!din_b[213]),
	.datac(!din_a[207]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_774 ),
	.cout(Xd_0__inst_mult_17_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_195 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[198]),
	.datac(!din_a[198]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_769 ),
	.cout(Xd_0__inst_mult_16_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_196 (
// Equation(s):

	.dataa(!din_a[196]),
	.datab(!din_b[201]),
	.datac(!din_a[195]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_774 ),
	.cout(Xd_0__inst_mult_16_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_195 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[234]),
	.datac(!din_a[234]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_769 ),
	.cout(Xd_0__inst_mult_19_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_196 (
// Equation(s):

	.dataa(!din_a[232]),
	.datab(!din_b[237]),
	.datac(!din_a[231]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_774 ),
	.cout(Xd_0__inst_mult_19_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_194 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_764 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_195 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[222]),
	.datac(!din_a[222]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_769 ),
	.cout(Xd_0__inst_mult_18_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_196 (
// Equation(s):

	.dataa(!din_a[220]),
	.datab(!din_b[225]),
	.datac(!din_a[219]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_774 ),
	.cout(Xd_0__inst_mult_18_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_195 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[162]),
	.datac(!din_a[162]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_769 ),
	.cout(Xd_0__inst_mult_13_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_196 (
// Equation(s):

	.dataa(!din_a[160]),
	.datab(!din_b[165]),
	.datac(!din_a[159]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_774 ),
	.cout(Xd_0__inst_mult_13_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_194 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_764 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_195 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[150]),
	.datac(!din_a[150]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_769 ),
	.cout(Xd_0__inst_mult_12_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_196 (
// Equation(s):

	.dataa(!din_a[148]),
	.datab(!din_b[153]),
	.datac(!din_a[147]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_774 ),
	.cout(Xd_0__inst_mult_12_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_194 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_764 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_195 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[186]),
	.datac(!din_a[186]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_769 ),
	.cout(Xd_0__inst_mult_15_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_196 (
// Equation(s):

	.dataa(!din_a[184]),
	.datab(!din_b[189]),
	.datac(!din_a[183]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_774 ),
	.cout(Xd_0__inst_mult_15_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_194 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_750 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_764 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_195 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[174]),
	.datac(!din_a[174]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_755 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_769 ),
	.cout(Xd_0__inst_mult_14_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_196 (
// Equation(s):

	.dataa(!din_a[172]),
	.datab(!din_b[177]),
	.datac(!din_a[171]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_774 ),
	.cout(Xd_0__inst_mult_14_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_195 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[114]),
	.datac(!din_a[114]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_769 ),
	.cout(Xd_0__inst_mult_9_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_196 (
// Equation(s):

	.dataa(!din_a[112]),
	.datab(!din_b[117]),
	.datac(!din_a[111]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_774 ),
	.cout(Xd_0__inst_mult_9_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_195 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[102]),
	.datac(!din_a[102]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_769 ),
	.cout(Xd_0__inst_mult_8_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_196 (
// Equation(s):

	.dataa(!din_a[100]),
	.datab(!din_b[105]),
	.datac(!din_a[99]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_774 ),
	.cout(Xd_0__inst_mult_8_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_195 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[138]),
	.datac(!din_a[138]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_769 ),
	.cout(Xd_0__inst_mult_11_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_196 (
// Equation(s):

	.dataa(!din_a[136]),
	.datab(!din_b[141]),
	.datac(!din_a[135]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_774 ),
	.cout(Xd_0__inst_mult_11_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_195 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[126]),
	.datac(!din_a[126]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_769 ),
	.cout(Xd_0__inst_mult_10_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_196 (
// Equation(s):

	.dataa(!din_a[124]),
	.datab(!din_b[129]),
	.datac(!din_a[123]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_774 ),
	.cout(Xd_0__inst_mult_10_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_195 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[66]),
	.datac(!din_a[66]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_769 ),
	.cout(Xd_0__inst_mult_5_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_196 (
// Equation(s):

	.dataa(!din_a[64]),
	.datab(!din_b[69]),
	.datac(!din_a[63]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_774 ),
	.cout(Xd_0__inst_mult_5_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_195 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[54]),
	.datac(!din_a[54]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_769 ),
	.cout(Xd_0__inst_mult_4_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_196 (
// Equation(s):

	.dataa(!din_a[52]),
	.datab(!din_b[57]),
	.datac(!din_a[51]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_774 ),
	.cout(Xd_0__inst_mult_4_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_195 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[90]),
	.datac(!din_a[90]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_769 ),
	.cout(Xd_0__inst_mult_7_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_196 (
// Equation(s):

	.dataa(!din_a[88]),
	.datab(!din_b[93]),
	.datac(!din_a[87]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_774 ),
	.cout(Xd_0__inst_mult_7_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_195 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[78]),
	.datac(!din_a[78]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_769 ),
	.cout(Xd_0__inst_mult_6_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_196 (
// Equation(s):

	.dataa(!din_a[76]),
	.datab(!din_b[81]),
	.datac(!din_a[75]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_774 ),
	.cout(Xd_0__inst_mult_6_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_195 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[18]),
	.datac(!din_a[18]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_769 ),
	.cout(Xd_0__inst_mult_1_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_196 (
// Equation(s):

	.dataa(!din_a[16]),
	.datab(!din_b[21]),
	.datac(!din_a[15]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_774 ),
	.cout(Xd_0__inst_mult_1_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_195 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[6]),
	.datac(!din_a[6]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_769 ),
	.cout(Xd_0__inst_mult_0_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_196 (
// Equation(s):

	.dataa(!din_a[4]),
	.datab(!din_b[9]),
	.datac(!din_a[3]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_774 ),
	.cout(Xd_0__inst_mult_0_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_195 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[42]),
	.datac(!din_a[42]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_760 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_769 ),
	.cout(Xd_0__inst_mult_3_770 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_196 (
// Equation(s):

	.dataa(!din_a[40]),
	.datab(!din_b[45]),
	.datac(!din_a[39]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_765 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_774 ),
	.cout(Xd_0__inst_mult_3_775 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_199 (
// Equation(s):

	.dataa(!din_a[28]),
	.datab(!din_b[33]),
	.datac(!din_a[27]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_789 ),
	.cout(Xd_0__inst_mult_2_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_197 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[354]),
	.datac(!din_a[355]),
	.datad(!din_b[355]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_779 ),
	.cout(Xd_0__inst_mult_29_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_198 (
// Equation(s):

	.dataa(!din_a[353]),
	.datab(!din_b[357]),
	.datac(!din_a[352]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_784 ),
	.cout(Xd_0__inst_mult_29_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_197 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[342]),
	.datac(!din_a[343]),
	.datad(!din_b[343]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_779 ),
	.cout(Xd_0__inst_mult_28_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_198 (
// Equation(s):

	.dataa(!din_a[341]),
	.datab(!din_b[345]),
	.datac(!din_a[340]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_784 ),
	.cout(Xd_0__inst_mult_28_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_197 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[378]),
	.datac(!din_a[379]),
	.datad(!din_b[379]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_779 ),
	.cout(Xd_0__inst_mult_31_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_198 (
// Equation(s):

	.dataa(!din_a[377]),
	.datab(!din_b[381]),
	.datac(!din_a[376]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_784 ),
	.cout(Xd_0__inst_mult_31_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_197 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[366]),
	.datac(!din_a[367]),
	.datad(!din_b[367]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_779 ),
	.cout(Xd_0__inst_mult_30_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_198 (
// Equation(s):

	.dataa(!din_a[365]),
	.datab(!din_b[369]),
	.datac(!din_a[364]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_784 ),
	.cout(Xd_0__inst_mult_30_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_197 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[306]),
	.datac(!din_a[307]),
	.datad(!din_b[307]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_779 ),
	.cout(Xd_0__inst_mult_25_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_198 (
// Equation(s):

	.dataa(!din_a[305]),
	.datab(!din_b[309]),
	.datac(!din_a[304]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_784 ),
	.cout(Xd_0__inst_mult_25_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_197 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[330]),
	.datac(!din_a[331]),
	.datad(!din_b[331]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_779 ),
	.cout(Xd_0__inst_mult_27_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_198 (
// Equation(s):

	.dataa(!din_a[329]),
	.datab(!din_b[333]),
	.datac(!din_a[328]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_784 ),
	.cout(Xd_0__inst_mult_27_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_197 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[258]),
	.datac(!din_a[259]),
	.datad(!din_b[259]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_779 ),
	.cout(Xd_0__inst_mult_21_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_198 (
// Equation(s):

	.dataa(!din_a[257]),
	.datab(!din_b[261]),
	.datac(!din_a[256]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_784 ),
	.cout(Xd_0__inst_mult_21_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_197 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[246]),
	.datac(!din_a[247]),
	.datad(!din_b[247]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_779 ),
	.cout(Xd_0__inst_mult_20_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_198 (
// Equation(s):

	.dataa(!din_a[245]),
	.datab(!din_b[249]),
	.datac(!din_a[244]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_784 ),
	.cout(Xd_0__inst_mult_20_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_197 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[282]),
	.datac(!din_a[283]),
	.datad(!din_b[283]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_779 ),
	.cout(Xd_0__inst_mult_23_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_198 (
// Equation(s):

	.dataa(!din_a[281]),
	.datab(!din_b[285]),
	.datac(!din_a[280]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_784 ),
	.cout(Xd_0__inst_mult_23_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_197 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[270]),
	.datac(!din_a[271]),
	.datad(!din_b[271]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_779 ),
	.cout(Xd_0__inst_mult_22_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_198 (
// Equation(s):

	.dataa(!din_a[269]),
	.datab(!din_b[273]),
	.datac(!din_a[268]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_784 ),
	.cout(Xd_0__inst_mult_22_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_197 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[210]),
	.datac(!din_a[211]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_779 ),
	.cout(Xd_0__inst_mult_17_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_198 (
// Equation(s):

	.dataa(!din_a[209]),
	.datab(!din_b[213]),
	.datac(!din_a[208]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_784 ),
	.cout(Xd_0__inst_mult_17_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_197 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[198]),
	.datac(!din_a[199]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_779 ),
	.cout(Xd_0__inst_mult_16_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_198 (
// Equation(s):

	.dataa(!din_a[197]),
	.datab(!din_b[201]),
	.datac(!din_a[196]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_784 ),
	.cout(Xd_0__inst_mult_16_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_197 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[234]),
	.datac(!din_a[235]),
	.datad(!din_b[235]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_779 ),
	.cout(Xd_0__inst_mult_19_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_198 (
// Equation(s):

	.dataa(!din_a[233]),
	.datab(!din_b[237]),
	.datac(!din_a[232]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_784 ),
	.cout(Xd_0__inst_mult_19_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_197 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[222]),
	.datac(!din_a[223]),
	.datad(!din_b[223]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_779 ),
	.cout(Xd_0__inst_mult_18_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_198 (
// Equation(s):

	.dataa(!din_a[221]),
	.datab(!din_b[225]),
	.datac(!din_a[220]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_784 ),
	.cout(Xd_0__inst_mult_18_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_197 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[162]),
	.datac(!din_a[163]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_779 ),
	.cout(Xd_0__inst_mult_13_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_198 (
// Equation(s):

	.dataa(!din_a[161]),
	.datab(!din_b[165]),
	.datac(!din_a[160]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_784 ),
	.cout(Xd_0__inst_mult_13_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_197 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[150]),
	.datac(!din_a[151]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_779 ),
	.cout(Xd_0__inst_mult_12_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_198 (
// Equation(s):

	.dataa(!din_a[149]),
	.datab(!din_b[153]),
	.datac(!din_a[148]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_784 ),
	.cout(Xd_0__inst_mult_12_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_197 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[186]),
	.datac(!din_a[187]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_779 ),
	.cout(Xd_0__inst_mult_15_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_198 (
// Equation(s):

	.dataa(!din_a[185]),
	.datab(!din_b[189]),
	.datac(!din_a[184]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_784 ),
	.cout(Xd_0__inst_mult_15_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_197 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[174]),
	.datac(!din_a[175]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_779 ),
	.cout(Xd_0__inst_mult_14_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_198 (
// Equation(s):

	.dataa(!din_a[173]),
	.datab(!din_b[177]),
	.datac(!din_a[172]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_784 ),
	.cout(Xd_0__inst_mult_14_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_197 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[114]),
	.datac(!din_a[115]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_779 ),
	.cout(Xd_0__inst_mult_9_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_198 (
// Equation(s):

	.dataa(!din_a[113]),
	.datab(!din_b[117]),
	.datac(!din_a[112]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_784 ),
	.cout(Xd_0__inst_mult_9_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_197 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[102]),
	.datac(!din_a[103]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_779 ),
	.cout(Xd_0__inst_mult_8_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_198 (
// Equation(s):

	.dataa(!din_a[101]),
	.datab(!din_b[105]),
	.datac(!din_a[100]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_784 ),
	.cout(Xd_0__inst_mult_8_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_197 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[138]),
	.datac(!din_a[139]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_779 ),
	.cout(Xd_0__inst_mult_11_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_198 (
// Equation(s):

	.dataa(!din_a[137]),
	.datab(!din_b[141]),
	.datac(!din_a[136]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_784 ),
	.cout(Xd_0__inst_mult_11_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_197 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[126]),
	.datac(!din_a[127]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_779 ),
	.cout(Xd_0__inst_mult_10_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_198 (
// Equation(s):

	.dataa(!din_a[125]),
	.datab(!din_b[129]),
	.datac(!din_a[124]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_784 ),
	.cout(Xd_0__inst_mult_10_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_197 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[66]),
	.datac(!din_a[67]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_779 ),
	.cout(Xd_0__inst_mult_5_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_198 (
// Equation(s):

	.dataa(!din_a[65]),
	.datab(!din_b[69]),
	.datac(!din_a[64]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_784 ),
	.cout(Xd_0__inst_mult_5_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_197 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[54]),
	.datac(!din_a[55]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_779 ),
	.cout(Xd_0__inst_mult_4_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_198 (
// Equation(s):

	.dataa(!din_a[53]),
	.datab(!din_b[57]),
	.datac(!din_a[52]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_784 ),
	.cout(Xd_0__inst_mult_4_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_197 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[90]),
	.datac(!din_a[91]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_779 ),
	.cout(Xd_0__inst_mult_7_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_198 (
// Equation(s):

	.dataa(!din_a[89]),
	.datab(!din_b[93]),
	.datac(!din_a[88]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_784 ),
	.cout(Xd_0__inst_mult_7_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_197 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[78]),
	.datac(!din_a[79]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_779 ),
	.cout(Xd_0__inst_mult_6_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_198 (
// Equation(s):

	.dataa(!din_a[77]),
	.datab(!din_b[81]),
	.datac(!din_a[76]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_784 ),
	.cout(Xd_0__inst_mult_6_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_197 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[18]),
	.datac(!din_a[19]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_779 ),
	.cout(Xd_0__inst_mult_1_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_198 (
// Equation(s):

	.dataa(!din_a[17]),
	.datab(!din_b[21]),
	.datac(!din_a[16]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_784 ),
	.cout(Xd_0__inst_mult_1_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_197 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[6]),
	.datac(!din_a[7]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_779 ),
	.cout(Xd_0__inst_mult_0_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_198 (
// Equation(s):

	.dataa(!din_a[5]),
	.datab(!din_b[9]),
	.datac(!din_a[4]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_784 ),
	.cout(Xd_0__inst_mult_0_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_197 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[42]),
	.datac(!din_a[43]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_770 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_779 ),
	.cout(Xd_0__inst_mult_3_780 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_198 (
// Equation(s):

	.dataa(!din_a[41]),
	.datab(!din_b[45]),
	.datac(!din_a[40]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_775 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_784 ),
	.cout(Xd_0__inst_mult_3_785 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_200 (
// Equation(s):

	.dataa(!din_a[29]),
	.datab(!din_b[33]),
	.datac(!din_a[28]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_794 ),
	.cout(Xd_0__inst_mult_2_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_199 (
// Equation(s):

	.dataa(!din_a[356]),
	.datab(!din_b[355]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_789 ),
	.cout(Xd_0__inst_mult_29_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_200 (
// Equation(s):

	.dataa(!din_a[354]),
	.datab(!din_b[357]),
	.datac(!din_a[353]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_794 ),
	.cout(Xd_0__inst_mult_29_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_199 (
// Equation(s):

	.dataa(!din_a[344]),
	.datab(!din_b[343]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_789 ),
	.cout(Xd_0__inst_mult_28_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_200 (
// Equation(s):

	.dataa(!din_a[342]),
	.datab(!din_b[345]),
	.datac(!din_a[341]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_794 ),
	.cout(Xd_0__inst_mult_28_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_199 (
// Equation(s):

	.dataa(!din_a[380]),
	.datab(!din_b[379]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_789 ),
	.cout(Xd_0__inst_mult_31_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_200 (
// Equation(s):

	.dataa(!din_a[378]),
	.datab(!din_b[381]),
	.datac(!din_a[377]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_794 ),
	.cout(Xd_0__inst_mult_31_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_199 (
// Equation(s):

	.dataa(!din_a[368]),
	.datab(!din_b[367]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_789 ),
	.cout(Xd_0__inst_mult_30_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_200 (
// Equation(s):

	.dataa(!din_a[366]),
	.datab(!din_b[369]),
	.datac(!din_a[365]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_794 ),
	.cout(Xd_0__inst_mult_30_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_199 (
// Equation(s):

	.dataa(!din_a[308]),
	.datab(!din_b[307]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_789 ),
	.cout(Xd_0__inst_mult_25_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_200 (
// Equation(s):

	.dataa(!din_a[306]),
	.datab(!din_b[309]),
	.datac(!din_a[305]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_794 ),
	.cout(Xd_0__inst_mult_25_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_199 (
// Equation(s):

	.dataa(!din_a[332]),
	.datab(!din_b[331]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_789 ),
	.cout(Xd_0__inst_mult_27_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_200 (
// Equation(s):

	.dataa(!din_a[330]),
	.datab(!din_b[333]),
	.datac(!din_a[329]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_794 ),
	.cout(Xd_0__inst_mult_27_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_199 (
// Equation(s):

	.dataa(!din_a[260]),
	.datab(!din_b[259]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_789 ),
	.cout(Xd_0__inst_mult_21_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_200 (
// Equation(s):

	.dataa(!din_a[258]),
	.datab(!din_b[261]),
	.datac(!din_a[257]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_794 ),
	.cout(Xd_0__inst_mult_21_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_199 (
// Equation(s):

	.dataa(!din_a[248]),
	.datab(!din_b[247]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_789 ),
	.cout(Xd_0__inst_mult_20_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_200 (
// Equation(s):

	.dataa(!din_a[246]),
	.datab(!din_b[249]),
	.datac(!din_a[245]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_794 ),
	.cout(Xd_0__inst_mult_20_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_199 (
// Equation(s):

	.dataa(!din_a[284]),
	.datab(!din_b[283]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_789 ),
	.cout(Xd_0__inst_mult_23_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_200 (
// Equation(s):

	.dataa(!din_a[282]),
	.datab(!din_b[285]),
	.datac(!din_a[281]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_794 ),
	.cout(Xd_0__inst_mult_23_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_199 (
// Equation(s):

	.dataa(!din_a[272]),
	.datab(!din_b[271]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_789 ),
	.cout(Xd_0__inst_mult_22_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_200 (
// Equation(s):

	.dataa(!din_a[270]),
	.datab(!din_b[273]),
	.datac(!din_a[269]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_794 ),
	.cout(Xd_0__inst_mult_22_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_199 (
// Equation(s):

	.dataa(!din_a[212]),
	.datab(!din_b[211]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_789 ),
	.cout(Xd_0__inst_mult_17_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_200 (
// Equation(s):

	.dataa(!din_a[210]),
	.datab(!din_b[213]),
	.datac(!din_a[209]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_794 ),
	.cout(Xd_0__inst_mult_17_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_199 (
// Equation(s):

	.dataa(!din_a[200]),
	.datab(!din_b[199]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_789 ),
	.cout(Xd_0__inst_mult_16_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_200 (
// Equation(s):

	.dataa(!din_a[198]),
	.datab(!din_b[201]),
	.datac(!din_a[197]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_794 ),
	.cout(Xd_0__inst_mult_16_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_199 (
// Equation(s):

	.dataa(!din_a[236]),
	.datab(!din_b[235]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_789 ),
	.cout(Xd_0__inst_mult_19_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_200 (
// Equation(s):

	.dataa(!din_a[234]),
	.datab(!din_b[237]),
	.datac(!din_a[233]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_794 ),
	.cout(Xd_0__inst_mult_19_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_199 (
// Equation(s):

	.dataa(!din_a[224]),
	.datab(!din_b[223]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_789 ),
	.cout(Xd_0__inst_mult_18_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_200 (
// Equation(s):

	.dataa(!din_a[222]),
	.datab(!din_b[225]),
	.datac(!din_a[221]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_794 ),
	.cout(Xd_0__inst_mult_18_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_199 (
// Equation(s):

	.dataa(!din_a[164]),
	.datab(!din_b[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_789 ),
	.cout(Xd_0__inst_mult_13_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_200 (
// Equation(s):

	.dataa(!din_a[162]),
	.datab(!din_b[165]),
	.datac(!din_a[161]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_794 ),
	.cout(Xd_0__inst_mult_13_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_199 (
// Equation(s):

	.dataa(!din_a[152]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_789 ),
	.cout(Xd_0__inst_mult_12_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_200 (
// Equation(s):

	.dataa(!din_a[150]),
	.datab(!din_b[153]),
	.datac(!din_a[149]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_794 ),
	.cout(Xd_0__inst_mult_12_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_199 (
// Equation(s):

	.dataa(!din_a[188]),
	.datab(!din_b[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_789 ),
	.cout(Xd_0__inst_mult_15_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_200 (
// Equation(s):

	.dataa(!din_a[186]),
	.datab(!din_b[189]),
	.datac(!din_a[185]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_794 ),
	.cout(Xd_0__inst_mult_15_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_199 (
// Equation(s):

	.dataa(!din_a[176]),
	.datab(!din_b[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_789 ),
	.cout(Xd_0__inst_mult_14_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_200 (
// Equation(s):

	.dataa(!din_a[174]),
	.datab(!din_b[177]),
	.datac(!din_a[173]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_794 ),
	.cout(Xd_0__inst_mult_14_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_199 (
// Equation(s):

	.dataa(!din_a[116]),
	.datab(!din_b[115]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_789 ),
	.cout(Xd_0__inst_mult_9_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_200 (
// Equation(s):

	.dataa(!din_a[114]),
	.datab(!din_b[117]),
	.datac(!din_a[113]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_794 ),
	.cout(Xd_0__inst_mult_9_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_199 (
// Equation(s):

	.dataa(!din_a[104]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_789 ),
	.cout(Xd_0__inst_mult_8_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_200 (
// Equation(s):

	.dataa(!din_a[102]),
	.datab(!din_b[105]),
	.datac(!din_a[101]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_794 ),
	.cout(Xd_0__inst_mult_8_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_199 (
// Equation(s):

	.dataa(!din_a[140]),
	.datab(!din_b[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_789 ),
	.cout(Xd_0__inst_mult_11_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_200 (
// Equation(s):

	.dataa(!din_a[138]),
	.datab(!din_b[141]),
	.datac(!din_a[137]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_794 ),
	.cout(Xd_0__inst_mult_11_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_199 (
// Equation(s):

	.dataa(!din_a[128]),
	.datab(!din_b[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_789 ),
	.cout(Xd_0__inst_mult_10_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_200 (
// Equation(s):

	.dataa(!din_a[126]),
	.datab(!din_b[129]),
	.datac(!din_a[125]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_794 ),
	.cout(Xd_0__inst_mult_10_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_199 (
// Equation(s):

	.dataa(!din_a[68]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_789 ),
	.cout(Xd_0__inst_mult_5_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_200 (
// Equation(s):

	.dataa(!din_a[66]),
	.datab(!din_b[69]),
	.datac(!din_a[65]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_794 ),
	.cout(Xd_0__inst_mult_5_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_199 (
// Equation(s):

	.dataa(!din_a[56]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_789 ),
	.cout(Xd_0__inst_mult_4_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_200 (
// Equation(s):

	.dataa(!din_a[54]),
	.datab(!din_b[57]),
	.datac(!din_a[53]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_794 ),
	.cout(Xd_0__inst_mult_4_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_199 (
// Equation(s):

	.dataa(!din_a[92]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_789 ),
	.cout(Xd_0__inst_mult_7_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_200 (
// Equation(s):

	.dataa(!din_a[90]),
	.datab(!din_b[93]),
	.datac(!din_a[89]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_794 ),
	.cout(Xd_0__inst_mult_7_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_199 (
// Equation(s):

	.dataa(!din_a[80]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_789 ),
	.cout(Xd_0__inst_mult_6_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_200 (
// Equation(s):

	.dataa(!din_a[78]),
	.datab(!din_b[81]),
	.datac(!din_a[77]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_794 ),
	.cout(Xd_0__inst_mult_6_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_199 (
// Equation(s):

	.dataa(!din_a[20]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_789 ),
	.cout(Xd_0__inst_mult_1_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_200 (
// Equation(s):

	.dataa(!din_a[18]),
	.datab(!din_b[21]),
	.datac(!din_a[17]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_794 ),
	.cout(Xd_0__inst_mult_1_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_199 (
// Equation(s):

	.dataa(!din_a[8]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_789 ),
	.cout(Xd_0__inst_mult_0_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_200 (
// Equation(s):

	.dataa(!din_a[6]),
	.datab(!din_b[9]),
	.datac(!din_a[5]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_794 ),
	.cout(Xd_0__inst_mult_0_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_199 (
// Equation(s):

	.dataa(!din_a[44]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_780 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_789 ),
	.cout(Xd_0__inst_mult_3_790 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_200 (
// Equation(s):

	.dataa(!din_a[42]),
	.datab(!din_b[45]),
	.datac(!din_a[41]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_785 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_794 ),
	.cout(Xd_0__inst_mult_3_795 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_201 (
// Equation(s):

	.dataa(!din_a[30]),
	.datab(!din_b[33]),
	.datac(!din_a[29]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_799 ),
	.cout(Xd_0__inst_mult_2_800 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_29_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_29_202 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[357]),
	.datac(!din_a[354]),
	.datad(!din_b[358]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_804 ),
	.cout(Xd_0__inst_mult_29_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_28_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_28_202 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[345]),
	.datac(!din_a[342]),
	.datad(!din_b[346]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_804 ),
	.cout(Xd_0__inst_mult_28_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_31_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_31_202 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[381]),
	.datac(!din_a[378]),
	.datad(!din_b[382]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_804 ),
	.cout(Xd_0__inst_mult_31_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_30_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_30_202 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[369]),
	.datac(!din_a[366]),
	.datad(!din_b[370]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_804 ),
	.cout(Xd_0__inst_mult_30_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_25_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_25_202 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[309]),
	.datac(!din_a[306]),
	.datad(!din_b[310]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_804 ),
	.cout(Xd_0__inst_mult_25_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_27_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_27_202 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[333]),
	.datac(!din_a[330]),
	.datad(!din_b[334]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_804 ),
	.cout(Xd_0__inst_mult_27_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_21_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_21_202 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[261]),
	.datac(!din_a[258]),
	.datad(!din_b[262]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_804 ),
	.cout(Xd_0__inst_mult_21_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_20_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_20_202 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[249]),
	.datac(!din_a[246]),
	.datad(!din_b[250]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_804 ),
	.cout(Xd_0__inst_mult_20_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_23_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_23_202 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[285]),
	.datac(!din_a[282]),
	.datad(!din_b[286]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_804 ),
	.cout(Xd_0__inst_mult_23_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_22_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_22_202 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[273]),
	.datac(!din_a[270]),
	.datad(!din_b[274]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_804 ),
	.cout(Xd_0__inst_mult_22_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_17_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_17_202 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[213]),
	.datac(!din_a[210]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_804 ),
	.cout(Xd_0__inst_mult_17_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_16_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_16_202 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[201]),
	.datac(!din_a[198]),
	.datad(!din_b[202]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_804 ),
	.cout(Xd_0__inst_mult_16_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_19_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_19_202 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[237]),
	.datac(!din_a[234]),
	.datad(!din_b[238]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_804 ),
	.cout(Xd_0__inst_mult_19_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_18_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_18_202 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[225]),
	.datac(!din_a[222]),
	.datad(!din_b[226]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_804 ),
	.cout(Xd_0__inst_mult_18_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_13_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_13_202 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[165]),
	.datac(!din_a[162]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_804 ),
	.cout(Xd_0__inst_mult_13_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_12_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_12_202 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[153]),
	.datac(!din_a[150]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_804 ),
	.cout(Xd_0__inst_mult_12_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_15_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_15_202 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[189]),
	.datac(!din_a[186]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_804 ),
	.cout(Xd_0__inst_mult_15_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_14_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_14_202 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[177]),
	.datac(!din_a[174]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_804 ),
	.cout(Xd_0__inst_mult_14_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_9_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_9_202 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[117]),
	.datac(!din_a[114]),
	.datad(!din_b[118]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_804 ),
	.cout(Xd_0__inst_mult_9_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_8_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_8_202 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[105]),
	.datac(!din_a[102]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_804 ),
	.cout(Xd_0__inst_mult_8_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_11_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_11_202 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[141]),
	.datac(!din_a[138]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_804 ),
	.cout(Xd_0__inst_mult_11_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_10_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_10_202 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[129]),
	.datac(!din_a[126]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_804 ),
	.cout(Xd_0__inst_mult_10_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_5_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_5_202 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[69]),
	.datac(!din_a[66]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_804 ),
	.cout(Xd_0__inst_mult_5_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_4_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_4_202 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[57]),
	.datac(!din_a[54]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_804 ),
	.cout(Xd_0__inst_mult_4_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_7_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_7_202 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[93]),
	.datac(!din_a[90]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_804 ),
	.cout(Xd_0__inst_mult_7_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_6_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_6_202 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[81]),
	.datac(!din_a[78]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_804 ),
	.cout(Xd_0__inst_mult_6_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_1_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_1_202 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[21]),
	.datac(!din_a[18]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_804 ),
	.cout(Xd_0__inst_mult_1_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_0_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_0_202 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[9]),
	.datac(!din_a[6]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_804 ),
	.cout(Xd_0__inst_mult_0_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("off")
) Xd_0__inst_mult_3_201 (
// Equation(s):

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_790 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_799 ),
	.cout(),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_3_202 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[45]),
	.datac(!din_a[42]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_795 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_804 ),
	.cout(Xd_0__inst_mult_3_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000000001111E),
	.shared_arith("off")
) Xd_0__inst_mult_2_202 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[33]),
	.datac(!din_a[30]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_800 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_804 ),
	.cout(Xd_0__inst_mult_2_805 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_29_203 (
// Equation(s):

	.dataa(!din_a[355]),
	.datab(!din_b[358]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_29_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_29_809 ),
	.cout(Xd_0__inst_mult_29_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_28_203 (
// Equation(s):

	.dataa(!din_a[343]),
	.datab(!din_b[346]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_28_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_28_809 ),
	.cout(Xd_0__inst_mult_28_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_31_203 (
// Equation(s):

	.dataa(!din_a[379]),
	.datab(!din_b[382]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_31_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_31_809 ),
	.cout(Xd_0__inst_mult_31_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_30_203 (
// Equation(s):

	.dataa(!din_a[367]),
	.datab(!din_b[370]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_30_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_30_809 ),
	.cout(Xd_0__inst_mult_30_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_25_203 (
// Equation(s):

	.dataa(!din_a[307]),
	.datab(!din_b[310]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_25_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_25_809 ),
	.cout(Xd_0__inst_mult_25_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_27_203 (
// Equation(s):

	.dataa(!din_a[331]),
	.datab(!din_b[334]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_27_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_27_809 ),
	.cout(Xd_0__inst_mult_27_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_21_203 (
// Equation(s):

	.dataa(!din_a[259]),
	.datab(!din_b[262]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_21_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_21_809 ),
	.cout(Xd_0__inst_mult_21_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_20_203 (
// Equation(s):

	.dataa(!din_a[247]),
	.datab(!din_b[250]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_20_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_20_809 ),
	.cout(Xd_0__inst_mult_20_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_23_203 (
// Equation(s):

	.dataa(!din_a[283]),
	.datab(!din_b[286]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_23_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_23_809 ),
	.cout(Xd_0__inst_mult_23_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_22_203 (
// Equation(s):

	.dataa(!din_a[271]),
	.datab(!din_b[274]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_22_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_22_809 ),
	.cout(Xd_0__inst_mult_22_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_17_203 (
// Equation(s):

	.dataa(!din_a[211]),
	.datab(!din_b[214]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_17_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_17_809 ),
	.cout(Xd_0__inst_mult_17_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_16_203 (
// Equation(s):

	.dataa(!din_a[199]),
	.datab(!din_b[202]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_16_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_16_809 ),
	.cout(Xd_0__inst_mult_16_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_19_203 (
// Equation(s):

	.dataa(!din_a[235]),
	.datab(!din_b[238]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_19_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_19_809 ),
	.cout(Xd_0__inst_mult_19_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_18_203 (
// Equation(s):

	.dataa(!din_a[223]),
	.datab(!din_b[226]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_18_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_18_809 ),
	.cout(Xd_0__inst_mult_18_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_13_203 (
// Equation(s):

	.dataa(!din_a[163]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_13_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_13_809 ),
	.cout(Xd_0__inst_mult_13_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_12_203 (
// Equation(s):

	.dataa(!din_a[151]),
	.datab(!din_b[154]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_12_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_12_809 ),
	.cout(Xd_0__inst_mult_12_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_15_203 (
// Equation(s):

	.dataa(!din_a[187]),
	.datab(!din_b[190]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_15_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_15_809 ),
	.cout(Xd_0__inst_mult_15_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_14_203 (
// Equation(s):

	.dataa(!din_a[175]),
	.datab(!din_b[178]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_14_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_14_809 ),
	.cout(Xd_0__inst_mult_14_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_9_203 (
// Equation(s):

	.dataa(!din_a[115]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_9_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_9_809 ),
	.cout(Xd_0__inst_mult_9_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_8_203 (
// Equation(s):

	.dataa(!din_a[103]),
	.datab(!din_b[106]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_8_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_8_809 ),
	.cout(Xd_0__inst_mult_8_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_11_203 (
// Equation(s):

	.dataa(!din_a[139]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_11_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_11_809 ),
	.cout(Xd_0__inst_mult_11_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_10_203 (
// Equation(s):

	.dataa(!din_a[127]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_10_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_10_809 ),
	.cout(Xd_0__inst_mult_10_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_5_203 (
// Equation(s):

	.dataa(!din_a[67]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_5_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_5_809 ),
	.cout(Xd_0__inst_mult_5_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_4_203 (
// Equation(s):

	.dataa(!din_a[55]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_4_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_4_809 ),
	.cout(Xd_0__inst_mult_4_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_7_203 (
// Equation(s):

	.dataa(!din_a[91]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_7_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_7_809 ),
	.cout(Xd_0__inst_mult_7_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_6_203 (
// Equation(s):

	.dataa(!din_a[79]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_6_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_6_809 ),
	.cout(Xd_0__inst_mult_6_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_1_203 (
// Equation(s):

	.dataa(!din_a[19]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_1_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_1_809 ),
	.cout(Xd_0__inst_mult_1_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_0_203 (
// Equation(s):

	.dataa(!din_a[7]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_0_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_0_809 ),
	.cout(Xd_0__inst_mult_0_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_3_203 (
// Equation(s):

	.dataa(!din_a[43]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_3_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_3_809 ),
	.cout(Xd_0__inst_mult_3_810 ),
	.shareout());

fourteennm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("off")
) Xd_0__inst_mult_2_203 (
// Equation(s):

	.dataa(!din_a[31]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.datah(gnd),
	.cin(Xd_0__inst_mult_2_805 ),
	.sharein(),
	.combout(),
	.sumout(Xd_0__inst_mult_2_809 ),
	.cout(Xd_0__inst_mult_2_810 ),
	.shareout());

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [20]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [21]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [22]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [23]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [24]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [25]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_26_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_131_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [26]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_inst_dout_27_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_136_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [27]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_1__26_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_1_131_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__26__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_inst_first_level_0__26_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_131_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__26__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_3__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_3_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_2__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_1__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_1_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_inst_first_level_0__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__25__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_7__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_7__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_7__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_6__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_6__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_6__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_5__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_5__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_5__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_4__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_4__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_4__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_3__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_3__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_3__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_2__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_2__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_2__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_1__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_1__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_1__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum2_0__24_ (
	.clk(clk),
	.d(Xd_0__inst_a2_0__adder2_inst_add_0_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum2_0__24__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__22__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_14__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_15__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_12__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_13__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_10__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_11__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_8__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_9__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_6__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_7__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_4__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_5__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_3__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sum1_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_add_0_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__23__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_31_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [31]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_27_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [27]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_23_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [23]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_19_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_r_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sign [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_30_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [30]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_28_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [28]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_29_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [29]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_31_ (
	.clk(clk),
	.d(Xd_0__inst_i29_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [31]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_26_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [26]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_24_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [24]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_25_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [25]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_27_ (
	.clk(clk),
	.d(Xd_0__inst_i29_6_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [27]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_22_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [22]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_20_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [20]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_21_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [21]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_23_ (
	.clk(clk),
	.d(Xd_0__inst_i29_11_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [23]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_18_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_16_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_17_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_19_ (
	.clk(clk),
	.d(Xd_0__inst_i29_16_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [19]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_15_ (
	.clk(clk),
	.d(Xd_0__inst_i29_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [15]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_11_ (
	.clk(clk),
	.d(Xd_0__inst_i29_26_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [11]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i29_31_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i29_36_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_210 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__10__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_234 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__11__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__12__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__13__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__14__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__15__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__16__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__17__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__18__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_274 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__19__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__20__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_29__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_28__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_31__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_30__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_25__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_24__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_27__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_26__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_21__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_20__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_23__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_22__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_17__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_16__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_19__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_18__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_13__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_12__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_15__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_14__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_9__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_8__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_11__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_10__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__21__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_30_ (
	.clk(clk),
	.d(Xd_0__inst_i29_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [30]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_28_ (
	.clk(clk),
	.d(Xd_0__inst_i29_46_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [28]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_29_ (
	.clk(clk),
	.d(Xd_0__inst_i29_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [29]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_26_ (
	.clk(clk),
	.d(Xd_0__inst_i29_56_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [26]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_24_ (
	.clk(clk),
	.d(Xd_0__inst_i29_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [24]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_25_ (
	.clk(clk),
	.d(Xd_0__inst_i29_66_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [25]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_22_ (
	.clk(clk),
	.d(Xd_0__inst_i29_71_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [22]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_20_ (
	.clk(clk),
	.d(Xd_0__inst_i29_76_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [20]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_21_ (
	.clk(clk),
	.d(Xd_0__inst_i29_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [21]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_18_ (
	.clk(clk),
	.d(Xd_0__inst_i29_86_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [18]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_16_ (
	.clk(clk),
	.d(Xd_0__inst_i29_91_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [16]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_17_ (
	.clk(clk),
	.d(Xd_0__inst_i29_96_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [17]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_14_ (
	.clk(clk),
	.d(Xd_0__inst_i29_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [14]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_12_ (
	.clk(clk),
	.d(Xd_0__inst_i29_106_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [12]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_13_ (
	.clk(clk),
	.d(Xd_0__inst_i29_111_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [13]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_10_ (
	.clk(clk),
	.d(Xd_0__inst_i29_116_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [10]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_8_ (
	.clk(clk),
	.d(Xd_0__inst_i29_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [8]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_9_ (
	.clk(clk),
	.d(Xd_0__inst_i29_126_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [9]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i29_131_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i29_136_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i29_141_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i29_146_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i29_151_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i29_156_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_559 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_559 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_564 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_564 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_294 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_569 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_569 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__3__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_29__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_28__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_31__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_30__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_25__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_24__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_574 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_27__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_26__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_574 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_21__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_20__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_23__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_22__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_17__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_16__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_19__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_18__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_319 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_product1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__4__q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_654 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_659 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_654 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_659 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_339 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_664 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_669 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_664 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_669 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_674 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_679 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_674 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_679 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_254 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_594 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_684 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_619 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_684 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_374 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_529 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_689 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_554 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_689 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_694 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_694 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_389 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_394 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_354 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_619 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_599 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_369 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_399 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_514 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_309 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_554 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_514 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_534 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_409 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_414 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_519 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_269 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_519 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_419 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_424 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_329 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_16_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_17_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_524 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_239 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_379 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_524 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_359 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_429 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_434 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_299 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_349 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_18_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_19_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_22 (
	.clk(clk),
	.d(din_a[358]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_23 (
	.clk(clk),
	.d(din_b[353]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_22 (
	.clk(clk),
	.d(din_a[346]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_23 (
	.clk(clk),
	.d(din_b[341]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_22 (
	.clk(clk),
	.d(din_a[382]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_23 (
	.clk(clk),
	.d(din_b[377]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_22 (
	.clk(clk),
	.d(din_a[370]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_23 (
	.clk(clk),
	.d(din_b[365]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_529 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_22 (
	.clk(clk),
	.d(din_a[310]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_23 (
	.clk(clk),
	.d(din_b[305]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_219 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_334 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_22 (
	.clk(clk),
	.d(din_a[298]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_23 (
	.clk(clk),
	.d(din_b[293]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_529 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_22 (
	.clk(clk),
	.d(din_a[334]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_23 (
	.clk(clk),
	.d(din_b[329]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_314 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_22 (
	.clk(clk),
	.d(din_a[322]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_23 (
	.clk(clk),
	.d(din_b[317]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_22 (
	.clk(clk),
	.d(din_a[262]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_23 (
	.clk(clk),
	.d(din_b[257]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_22 (
	.clk(clk),
	.d(din_a[250]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_23 (
	.clk(clk),
	.d(din_b[245]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_22 (
	.clk(clk),
	.d(din_a[286]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_23 (
	.clk(clk),
	.d(din_b[281]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_22 (
	.clk(clk),
	.d(din_a[274]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_23 (
	.clk(clk),
	.d(din_b[269]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_22 (
	.clk(clk),
	.d(din_a[214]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_23 (
	.clk(clk),
	.d(din_b[209]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_22 (
	.clk(clk),
	.d(din_a[202]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_23 (
	.clk(clk),
	.d(din_b[197]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_484 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_22 (
	.clk(clk),
	.d(din_a[238]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_23 (
	.clk(clk),
	.d(din_b[233]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_22 (
	.clk(clk),
	.d(din_a[226]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_23 (
	.clk(clk),
	.d(din_b[221]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_22 (
	.clk(clk),
	.d(din_a[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_23 (
	.clk(clk),
	.d(din_b[161]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_22 (
	.clk(clk),
	.d(din_a[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_23 (
	.clk(clk),
	.d(din_b[149]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_22 (
	.clk(clk),
	.d(din_a[190]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_23 (
	.clk(clk),
	.d(din_b[185]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_439 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_444 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_22 (
	.clk(clk),
	.d(din_a[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_23 (
	.clk(clk),
	.d(din_b[173]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_22 (
	.clk(clk),
	.d(din_a[118]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_23 (
	.clk(clk),
	.d(din_b[113]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_22 (
	.clk(clk),
	.d(din_a[106]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_23 (
	.clk(clk),
	.d(din_b[101]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_22 (
	.clk(clk),
	.d(din_a[142]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_23 (
	.clk(clk),
	.d(din_b[137]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_22 (
	.clk(clk),
	.d(din_a[130]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_23 (
	.clk(clk),
	.d(din_b[125]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_22 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_23 (
	.clk(clk),
	.d(din_b[65]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_22 (
	.clk(clk),
	.d(din_a[58]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_23 (
	.clk(clk),
	.d(din_b[53]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_22 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_23 (
	.clk(clk),
	.d(din_b[89]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_22 (
	.clk(clk),
	.d(din_a[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_23 (
	.clk(clk),
	.d(din_b[77]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_22 (
	.clk(clk),
	.d(din_a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_23 (
	.clk(clk),
	.d(din_b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_22 (
	.clk(clk),
	.d(din_a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_23 (
	.clk(clk),
	.d(din_b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_22 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_23 (
	.clk(clk),
	.d(din_b[41]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_20_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_21_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_22 (
	.clk(clk),
	.d(din_a[34]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_22_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_23 (
	.clk(clk),
	.d(din_b[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_23_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_534 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_289 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_534 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_279 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_489 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_449 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_24_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_25_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_539 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_259 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_539 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_249 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_494 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_454 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_26_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_27_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_544 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_229 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_544 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_499 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_459 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_514 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_28_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_29_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_549 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_549 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_214 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_504 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_464 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_474 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_519 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_30_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_31_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_29_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_28_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_31_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_30_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_554 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_25_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_24_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_554 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_27_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_205 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_26_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_80_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_21_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_20_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_23_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_22_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_17_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_16_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_509 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_19_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_18_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_13_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_12_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_15_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_40_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_469 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_14_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_9_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_8_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_11_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_10_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_5_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_4_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_7_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_60_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_6_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_1_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_70_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_0_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_75_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_479 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_3_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_33_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_524 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_32_q ));

fourteennm_ff #(
	.is_wysiwyg("true"),
	.power_up()
) Xd_0__inst_mult_2_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_50_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.sclr1(gnd),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_33_q ));

assign dout[0] = Xd_0__inst_inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_inst_dout [15];

assign dout[16] = Xd_0__inst_inst_inst_inst_dout [16];

assign dout[17] = Xd_0__inst_inst_inst_inst_dout [17];

assign dout[18] = Xd_0__inst_inst_inst_inst_dout [18];

assign dout[19] = Xd_0__inst_inst_inst_inst_dout [19];

assign dout[20] = Xd_0__inst_inst_inst_inst_dout [20];

assign dout[21] = Xd_0__inst_inst_inst_inst_dout [21];

assign dout[22] = Xd_0__inst_inst_inst_inst_dout [22];

assign dout[23] = Xd_0__inst_inst_inst_inst_dout [23];

assign dout[24] = Xd_0__inst_inst_inst_inst_dout [24];

assign dout[25] = Xd_0__inst_inst_inst_inst_dout [25];

assign dout[26] = Xd_0__inst_inst_inst_inst_dout [26];

assign dout[27] = Xd_0__inst_inst_inst_inst_dout [27];

endmodule
