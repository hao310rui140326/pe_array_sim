// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:27:55"

// 
// Device: Altera 10AX115S2F45I1SG Package FBGA1932
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_a10_7x7x32 (
	dout,
	clk,
	din_a,
	din_b);
output 	[17:0] dout;
input 	clk;
input 	[223:0] din_a;
input 	[223:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_6 ;
wire Xd_0__inst_inst_inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_10 ;
wire Xd_0__inst_inst_inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_14 ;
wire Xd_0__inst_inst_inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_18 ;
wire Xd_0__inst_inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_26 ;
wire Xd_0__inst_inst_inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_30 ;
wire Xd_0__inst_inst_inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_34 ;
wire Xd_0__inst_inst_inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_38 ;
wire Xd_0__inst_inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_46 ;
wire Xd_0__inst_inst_inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_50 ;
wire Xd_0__inst_inst_inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_54 ;
wire Xd_0__inst_inst_inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_58 ;
wire Xd_0__inst_inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_inst_add_0_65_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_66 ;
wire Xd_0__inst_inst_inst_inst_add_0_69_sumout ;
wire Xd_0__inst_i19_1_sumout ;
wire Xd_0__inst_i19_2 ;
wire Xd_0__inst_inst_inst_add_3_1_sumout ;
wire Xd_0__inst_inst_inst_add_3_2 ;
wire Xd_0__inst_inst_inst_add_3_3 ;
wire Xd_0__inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_add_0_3 ;
wire Xd_0__inst_i19_5_sumout ;
wire Xd_0__inst_i19_6 ;
wire Xd_0__inst_inst_inst_add_3_5_sumout ;
wire Xd_0__inst_inst_inst_add_3_6 ;
wire Xd_0__inst_inst_inst_add_3_7 ;
wire Xd_0__inst_inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_inst_add_0_6 ;
wire Xd_0__inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_add_3_9_sumout ;
wire Xd_0__inst_inst_inst_add_3_10 ;
wire Xd_0__inst_inst_inst_add_3_11 ;
wire Xd_0__inst_inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_inst_add_0_10 ;
wire Xd_0__inst_inst_inst_add_0_11 ;
wire Xd_0__inst_inst_inst_add_3_13_sumout ;
wire Xd_0__inst_inst_inst_add_3_14 ;
wire Xd_0__inst_inst_inst_add_3_15 ;
wire Xd_0__inst_inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_inst_add_0_14 ;
wire Xd_0__inst_inst_inst_add_0_15 ;
wire Xd_0__inst_inst_inst_add_3_17_sumout ;
wire Xd_0__inst_inst_inst_add_3_18 ;
wire Xd_0__inst_inst_inst_add_3_19 ;
wire Xd_0__inst_inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_inst_add_0_18 ;
wire Xd_0__inst_inst_inst_add_0_19 ;
wire Xd_0__inst_inst_inst_add_3_21_sumout ;
wire Xd_0__inst_inst_inst_add_3_22 ;
wire Xd_0__inst_inst_inst_add_3_23 ;
wire Xd_0__inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_add_0_23 ;
wire Xd_0__inst_inst_inst_add_3_25_sumout ;
wire Xd_0__inst_inst_inst_add_3_26 ;
wire Xd_0__inst_inst_inst_add_3_27 ;
wire Xd_0__inst_inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_inst_add_0_26 ;
wire Xd_0__inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_add_3_29_sumout ;
wire Xd_0__inst_inst_inst_add_3_30 ;
wire Xd_0__inst_inst_inst_add_3_31 ;
wire Xd_0__inst_inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_inst_add_0_30 ;
wire Xd_0__inst_inst_inst_add_0_31 ;
wire Xd_0__inst_inst_inst_add_3_33_sumout ;
wire Xd_0__inst_inst_inst_add_3_34 ;
wire Xd_0__inst_inst_inst_add_3_35 ;
wire Xd_0__inst_inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_inst_add_0_34 ;
wire Xd_0__inst_inst_inst_add_0_35 ;
wire Xd_0__inst_inst_inst_add_3_37_sumout ;
wire Xd_0__inst_inst_inst_add_3_38 ;
wire Xd_0__inst_inst_inst_add_3_39 ;
wire Xd_0__inst_inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_inst_add_0_38 ;
wire Xd_0__inst_inst_inst_add_0_39 ;
wire Xd_0__inst_inst_inst_add_3_41_sumout ;
wire Xd_0__inst_inst_inst_add_3_42 ;
wire Xd_0__inst_inst_inst_add_3_43 ;
wire Xd_0__inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_add_0_43 ;
wire Xd_0__inst_inst_inst_add_3_45_sumout ;
wire Xd_0__inst_inst_inst_add_3_46 ;
wire Xd_0__inst_inst_inst_add_3_47 ;
wire Xd_0__inst_inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_inst_add_0_46 ;
wire Xd_0__inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_add_3_49_sumout ;
wire Xd_0__inst_inst_inst_add_3_50 ;
wire Xd_0__inst_inst_inst_add_3_51 ;
wire Xd_0__inst_inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_inst_add_0_50 ;
wire Xd_0__inst_inst_inst_add_0_51 ;
wire Xd_0__inst_inst_inst_add_3_53_sumout ;
wire Xd_0__inst_inst_inst_add_3_54 ;
wire Xd_0__inst_inst_inst_add_3_55 ;
wire Xd_0__inst_inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_inst_add_0_54 ;
wire Xd_0__inst_inst_inst_add_0_55 ;
wire Xd_0__inst_inst_inst_add_3_57_sumout ;
wire Xd_0__inst_inst_inst_add_3_58 ;
wire Xd_0__inst_inst_inst_add_3_59 ;
wire Xd_0__inst_inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_inst_add_0_58 ;
wire Xd_0__inst_inst_inst_add_0_59 ;
wire Xd_0__inst_inst_inst_add_3_61_sumout ;
wire Xd_0__inst_inst_inst_add_3_62 ;
wire Xd_0__inst_inst_inst_add_3_63 ;
wire Xd_0__inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_add_0_63 ;
wire Xd_0__inst_inst_inst_add_3_65_sumout ;
wire Xd_0__inst_inst_inst_add_3_66 ;
wire Xd_0__inst_inst_inst_add_3_67 ;
wire Xd_0__inst_inst_inst_add_0_65_sumout ;
wire Xd_0__inst_inst_inst_add_0_66 ;
wire Xd_0__inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_add_3_69_sumout ;
wire Xd_0__inst_inst_inst_add_0_69_sumout ;
wire Xd_0__inst_i19_9_sumout ;
wire Xd_0__inst_i19_10 ;
wire Xd_0__inst_i19_11 ;
wire Xd_0__inst_i19_13_sumout ;
wire Xd_0__inst_i19_14 ;
wire Xd_0__inst_i19_15 ;
wire Xd_0__inst_inst_add_8_1_sumout ;
wire Xd_0__inst_inst_add_8_2 ;
wire Xd_0__inst_inst_add_8_3 ;
wire Xd_0__inst_inst_add_6_1_sumout ;
wire Xd_0__inst_inst_add_6_2 ;
wire Xd_0__inst_inst_add_6_3 ;
wire Xd_0__inst_i19_17_sumout ;
wire Xd_0__inst_i19_18 ;
wire Xd_0__inst_i19_19 ;
wire Xd_0__inst_inst_add_4_1_sumout ;
wire Xd_0__inst_inst_add_4_2 ;
wire Xd_0__inst_inst_add_4_3 ;
wire Xd_0__inst_inst_add_2_1_sumout ;
wire Xd_0__inst_inst_add_2_2 ;
wire Xd_0__inst_inst_add_2_3 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_inst_add_0_3 ;
wire Xd_0__inst_inst_add_8_5_sumout ;
wire Xd_0__inst_inst_add_8_6 ;
wire Xd_0__inst_inst_add_8_7 ;
wire Xd_0__inst_inst_add_6_5_sumout ;
wire Xd_0__inst_inst_add_6_6 ;
wire Xd_0__inst_inst_add_6_7 ;
wire Xd_0__inst_inst_add_4_5_sumout ;
wire Xd_0__inst_inst_add_4_6 ;
wire Xd_0__inst_inst_add_4_7 ;
wire Xd_0__inst_inst_add_2_5_sumout ;
wire Xd_0__inst_inst_add_2_6 ;
wire Xd_0__inst_inst_add_2_7 ;
wire Xd_0__inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_add_0_6 ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_8_9_sumout ;
wire Xd_0__inst_inst_add_8_10 ;
wire Xd_0__inst_inst_add_8_11 ;
wire Xd_0__inst_inst_add_6_9_sumout ;
wire Xd_0__inst_inst_add_6_10 ;
wire Xd_0__inst_inst_add_6_11 ;
wire Xd_0__inst_inst_add_4_9_sumout ;
wire Xd_0__inst_inst_add_4_10 ;
wire Xd_0__inst_inst_add_4_11 ;
wire Xd_0__inst_inst_add_2_9_sumout ;
wire Xd_0__inst_inst_add_2_10 ;
wire Xd_0__inst_inst_add_2_11 ;
wire Xd_0__inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_add_0_10 ;
wire Xd_0__inst_inst_add_0_11 ;
wire Xd_0__inst_inst_add_8_13_sumout ;
wire Xd_0__inst_inst_add_8_14 ;
wire Xd_0__inst_inst_add_8_15 ;
wire Xd_0__inst_inst_add_6_13_sumout ;
wire Xd_0__inst_inst_add_6_14 ;
wire Xd_0__inst_inst_add_6_15 ;
wire Xd_0__inst_inst_add_4_13_sumout ;
wire Xd_0__inst_inst_add_4_14 ;
wire Xd_0__inst_inst_add_4_15 ;
wire Xd_0__inst_inst_add_2_13_sumout ;
wire Xd_0__inst_inst_add_2_14 ;
wire Xd_0__inst_inst_add_2_15 ;
wire Xd_0__inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_add_0_14 ;
wire Xd_0__inst_inst_add_0_15 ;
wire Xd_0__inst_inst_add_8_17_sumout ;
wire Xd_0__inst_inst_add_8_18 ;
wire Xd_0__inst_inst_add_8_19 ;
wire Xd_0__inst_inst_add_6_17_sumout ;
wire Xd_0__inst_inst_add_6_18 ;
wire Xd_0__inst_inst_add_6_19 ;
wire Xd_0__inst_inst_add_4_17_sumout ;
wire Xd_0__inst_inst_add_4_18 ;
wire Xd_0__inst_inst_add_4_19 ;
wire Xd_0__inst_inst_add_2_17_sumout ;
wire Xd_0__inst_inst_add_2_18 ;
wire Xd_0__inst_inst_add_2_19 ;
wire Xd_0__inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_add_0_18 ;
wire Xd_0__inst_inst_add_0_19 ;
wire Xd_0__inst_inst_add_8_21_sumout ;
wire Xd_0__inst_inst_add_8_22 ;
wire Xd_0__inst_inst_add_8_23 ;
wire Xd_0__inst_inst_add_6_21_sumout ;
wire Xd_0__inst_inst_add_6_22 ;
wire Xd_0__inst_inst_add_6_23 ;
wire Xd_0__inst_inst_add_4_21_sumout ;
wire Xd_0__inst_inst_add_4_22 ;
wire Xd_0__inst_inst_add_4_23 ;
wire Xd_0__inst_inst_add_2_21_sumout ;
wire Xd_0__inst_inst_add_2_22 ;
wire Xd_0__inst_inst_add_2_23 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_0_23 ;
wire Xd_0__inst_inst_add_8_25_sumout ;
wire Xd_0__inst_inst_add_8_26 ;
wire Xd_0__inst_inst_add_8_27 ;
wire Xd_0__inst_inst_add_6_25_sumout ;
wire Xd_0__inst_inst_add_6_26 ;
wire Xd_0__inst_inst_add_6_27 ;
wire Xd_0__inst_inst_add_4_25_sumout ;
wire Xd_0__inst_inst_add_4_26 ;
wire Xd_0__inst_inst_add_4_27 ;
wire Xd_0__inst_inst_add_2_25_sumout ;
wire Xd_0__inst_inst_add_2_26 ;
wire Xd_0__inst_inst_add_2_27 ;
wire Xd_0__inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_add_0_26 ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_8_29_sumout ;
wire Xd_0__inst_inst_add_8_30 ;
wire Xd_0__inst_inst_add_8_31 ;
wire Xd_0__inst_inst_add_6_29_sumout ;
wire Xd_0__inst_inst_add_6_30 ;
wire Xd_0__inst_inst_add_6_31 ;
wire Xd_0__inst_inst_add_4_29_sumout ;
wire Xd_0__inst_inst_add_4_30 ;
wire Xd_0__inst_inst_add_4_31 ;
wire Xd_0__inst_inst_add_2_29_sumout ;
wire Xd_0__inst_inst_add_2_30 ;
wire Xd_0__inst_inst_add_2_31 ;
wire Xd_0__inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_add_0_30 ;
wire Xd_0__inst_inst_add_0_31 ;
wire Xd_0__inst_inst_add_8_33_sumout ;
wire Xd_0__inst_inst_add_8_34 ;
wire Xd_0__inst_inst_add_8_35 ;
wire Xd_0__inst_inst_add_6_33_sumout ;
wire Xd_0__inst_inst_add_6_34 ;
wire Xd_0__inst_inst_add_6_35 ;
wire Xd_0__inst_inst_add_4_33_sumout ;
wire Xd_0__inst_inst_add_4_34 ;
wire Xd_0__inst_inst_add_4_35 ;
wire Xd_0__inst_inst_add_2_33_sumout ;
wire Xd_0__inst_inst_add_2_34 ;
wire Xd_0__inst_inst_add_2_35 ;
wire Xd_0__inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_add_0_34 ;
wire Xd_0__inst_inst_add_0_35 ;
wire Xd_0__inst_inst_add_8_37_sumout ;
wire Xd_0__inst_inst_add_8_38 ;
wire Xd_0__inst_inst_add_8_39 ;
wire Xd_0__inst_inst_add_6_37_sumout ;
wire Xd_0__inst_inst_add_6_38 ;
wire Xd_0__inst_inst_add_6_39 ;
wire Xd_0__inst_inst_add_4_37_sumout ;
wire Xd_0__inst_inst_add_4_38 ;
wire Xd_0__inst_inst_add_4_39 ;
wire Xd_0__inst_inst_add_2_37_sumout ;
wire Xd_0__inst_inst_add_2_38 ;
wire Xd_0__inst_inst_add_2_39 ;
wire Xd_0__inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_add_0_38 ;
wire Xd_0__inst_inst_add_0_39 ;
wire Xd_0__inst_inst_add_8_41_sumout ;
wire Xd_0__inst_inst_add_8_42 ;
wire Xd_0__inst_inst_add_8_43 ;
wire Xd_0__inst_inst_add_6_41_sumout ;
wire Xd_0__inst_inst_add_6_42 ;
wire Xd_0__inst_inst_add_6_43 ;
wire Xd_0__inst_inst_add_4_41_sumout ;
wire Xd_0__inst_inst_add_4_42 ;
wire Xd_0__inst_inst_add_4_43 ;
wire Xd_0__inst_inst_add_2_41_sumout ;
wire Xd_0__inst_inst_add_2_42 ;
wire Xd_0__inst_inst_add_2_43 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_0_43 ;
wire Xd_0__inst_inst_add_8_45_sumout ;
wire Xd_0__inst_inst_add_8_46 ;
wire Xd_0__inst_inst_add_8_47 ;
wire Xd_0__inst_inst_add_6_45_sumout ;
wire Xd_0__inst_inst_add_6_46 ;
wire Xd_0__inst_inst_add_6_47 ;
wire Xd_0__inst_inst_add_4_45_sumout ;
wire Xd_0__inst_inst_add_4_46 ;
wire Xd_0__inst_inst_add_4_47 ;
wire Xd_0__inst_inst_add_2_45_sumout ;
wire Xd_0__inst_inst_add_2_46 ;
wire Xd_0__inst_inst_add_2_47 ;
wire Xd_0__inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_add_0_46 ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_8_49_sumout ;
wire Xd_0__inst_inst_add_8_50 ;
wire Xd_0__inst_inst_add_8_51 ;
wire Xd_0__inst_inst_add_6_49_sumout ;
wire Xd_0__inst_inst_add_6_50 ;
wire Xd_0__inst_inst_add_6_51 ;
wire Xd_0__inst_inst_add_4_49_sumout ;
wire Xd_0__inst_inst_add_4_50 ;
wire Xd_0__inst_inst_add_4_51 ;
wire Xd_0__inst_inst_add_2_49_sumout ;
wire Xd_0__inst_inst_add_2_50 ;
wire Xd_0__inst_inst_add_2_51 ;
wire Xd_0__inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_add_0_50 ;
wire Xd_0__inst_inst_add_0_51 ;
wire Xd_0__inst_inst_add_8_53_sumout ;
wire Xd_0__inst_inst_add_8_54 ;
wire Xd_0__inst_inst_add_8_55 ;
wire Xd_0__inst_inst_add_6_53_sumout ;
wire Xd_0__inst_inst_add_6_54 ;
wire Xd_0__inst_inst_add_6_55 ;
wire Xd_0__inst_inst_add_4_53_sumout ;
wire Xd_0__inst_inst_add_4_54 ;
wire Xd_0__inst_inst_add_4_55 ;
wire Xd_0__inst_inst_add_2_53_sumout ;
wire Xd_0__inst_inst_add_2_54 ;
wire Xd_0__inst_inst_add_2_55 ;
wire Xd_0__inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_add_0_54 ;
wire Xd_0__inst_inst_add_0_55 ;
wire Xd_0__inst_inst_add_8_57_sumout ;
wire Xd_0__inst_inst_add_8_58 ;
wire Xd_0__inst_inst_add_8_59 ;
wire Xd_0__inst_inst_add_6_57_sumout ;
wire Xd_0__inst_inst_add_6_58 ;
wire Xd_0__inst_inst_add_6_59 ;
wire Xd_0__inst_inst_add_4_57_sumout ;
wire Xd_0__inst_inst_add_4_58 ;
wire Xd_0__inst_inst_add_4_59 ;
wire Xd_0__inst_inst_add_2_57_sumout ;
wire Xd_0__inst_inst_add_2_58 ;
wire Xd_0__inst_inst_add_2_59 ;
wire Xd_0__inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_add_0_58 ;
wire Xd_0__inst_inst_add_0_59 ;
wire Xd_0__inst_inst_add_8_61_sumout ;
wire Xd_0__inst_inst_add_6_61_sumout ;
wire Xd_0__inst_inst_add_4_61_sumout ;
wire Xd_0__inst_inst_add_2_61_sumout ;
wire Xd_0__inst_inst_add_0_61_sumout ;
wire Xd_0__inst_i19_21_sumout ;
wire Xd_0__inst_i19_22 ;
wire Xd_0__inst_i19_23 ;
wire Xd_0__inst_i19_25_sumout ;
wire Xd_0__inst_i19_26 ;
wire Xd_0__inst_i19_27 ;
wire Xd_0__inst_a1_15__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_29_sumout ;
wire Xd_0__inst_i19_30 ;
wire Xd_0__inst_i19_31 ;
wire Xd_0__inst_i19_33_sumout ;
wire Xd_0__inst_i19_34 ;
wire Xd_0__inst_i19_35 ;
wire Xd_0__inst_i19_37_sumout ;
wire Xd_0__inst_i19_38 ;
wire Xd_0__inst_i19_39 ;
wire Xd_0__inst_a1_15__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_41_sumout ;
wire Xd_0__inst_i19_42 ;
wire Xd_0__inst_i19_43 ;
wire Xd_0__inst_a1_11__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_45_sumout ;
wire Xd_0__inst_i19_46 ;
wire Xd_0__inst_i19_47 ;
wire Xd_0__inst_a1_8__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_49_sumout ;
wire Xd_0__inst_i19_50 ;
wire Xd_0__inst_i19_51 ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_53_sumout ;
wire Xd_0__inst_i19_54 ;
wire Xd_0__inst_i19_55 ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_i19_57_sumout ;
wire Xd_0__inst_i19_58 ;
wire Xd_0__inst_i19_59 ;
wire Xd_0__inst_a1_14__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_i19_61_sumout ;
wire Xd_0__inst_i19_62 ;
wire Xd_0__inst_i19_63 ;
wire Xd_0__inst_i19_65_sumout ;
wire Xd_0__inst_i19_66 ;
wire Xd_0__inst_i19_67 ;
wire Xd_0__inst_i19_69_sumout ;
wire Xd_0__inst_i19_70 ;
wire Xd_0__inst_i19_71 ;
wire Xd_0__inst_i19_73_sumout ;
wire Xd_0__inst_i19_74 ;
wire Xd_0__inst_i19_75 ;
wire Xd_0__inst_i19_77_sumout ;
wire Xd_0__inst_i19_78 ;
wire Xd_0__inst_i19_79 ;
wire Xd_0__inst_i19_81_sumout ;
wire Xd_0__inst_i19_82 ;
wire Xd_0__inst_i19_83 ;
wire Xd_0__inst_i19_85_sumout ;
wire Xd_0__inst_i19_86 ;
wire Xd_0__inst_i19_87 ;
wire Xd_0__inst_mult_30_49 ;
wire Xd_0__inst_mult_30_50 ;
wire Xd_0__inst_mult_30_51 ;
wire Xd_0__inst_mult_31_49 ;
wire Xd_0__inst_mult_31_50 ;
wire Xd_0__inst_mult_31_51 ;
wire Xd_0__inst_mult_30_53 ;
wire Xd_0__inst_mult_30_54 ;
wire Xd_0__inst_mult_30_55 ;
wire Xd_0__inst_mult_31_53 ;
wire Xd_0__inst_mult_31_54 ;
wire Xd_0__inst_mult_31_55 ;
wire Xd_0__inst_mult_30_56 ;
wire Xd_0__inst_mult_30_57 ;
wire Xd_0__inst_mult_30_58 ;
wire Xd_0__inst_mult_31_56 ;
wire Xd_0__inst_mult_31_57 ;
wire Xd_0__inst_mult_31_58 ;
wire Xd_0__inst_mult_30_60 ;
wire Xd_0__inst_mult_30_61 ;
wire Xd_0__inst_mult_30_62 ;
wire Xd_0__inst_mult_31_60 ;
wire Xd_0__inst_mult_31_61 ;
wire Xd_0__inst_mult_31_62 ;
wire Xd_0__inst_mult_30_64 ;
wire Xd_0__inst_mult_30_65 ;
wire Xd_0__inst_mult_30_66 ;
wire Xd_0__inst_mult_31_64 ;
wire Xd_0__inst_mult_31_65 ;
wire Xd_0__inst_mult_31_66 ;
wire Xd_0__inst_mult_30_68 ;
wire Xd_0__inst_mult_30_69 ;
wire Xd_0__inst_mult_30_70 ;
wire Xd_0__inst_mult_31_68 ;
wire Xd_0__inst_mult_31_69 ;
wire Xd_0__inst_mult_31_70 ;
wire Xd_0__inst_mult_30_72 ;
wire Xd_0__inst_mult_30_73 ;
wire Xd_0__inst_mult_30_74 ;
wire Xd_0__inst_mult_31_72 ;
wire Xd_0__inst_mult_31_73 ;
wire Xd_0__inst_mult_31_74 ;
wire Xd_0__inst_mult_30_76 ;
wire Xd_0__inst_mult_30_77 ;
wire Xd_0__inst_mult_30_78 ;
wire Xd_0__inst_mult_31_76 ;
wire Xd_0__inst_mult_31_77 ;
wire Xd_0__inst_mult_31_78 ;
wire Xd_0__inst_mult_30_80 ;
wire Xd_0__inst_mult_31_80 ;
wire Xd_0__inst_mult_31_81 ;
wire Xd_0__inst_mult_31_82 ;
wire Xd_0__inst_i19_89_sumout ;
wire Xd_0__inst_i19_90 ;
wire Xd_0__inst_i19_91 ;
wire Xd_0__inst_i19_93_sumout ;
wire Xd_0__inst_i19_94 ;
wire Xd_0__inst_i19_95 ;
wire Xd_0__inst_mult_30_84 ;
wire Xd_0__inst_mult_30_85 ;
wire Xd_0__inst_mult_30_86 ;
wire Xd_0__inst_mult_31_84 ;
wire Xd_0__inst_mult_31_85 ;
wire Xd_0__inst_mult_31_86 ;
wire Xd_0__inst_i19_97_sumout ;
wire Xd_0__inst_i19_98 ;
wire Xd_0__inst_i19_99 ;
wire Xd_0__inst_i19_101_sumout ;
wire Xd_0__inst_i19_102 ;
wire Xd_0__inst_i19_103 ;
wire Xd_0__inst_i19_105_sumout ;
wire Xd_0__inst_i19_106 ;
wire Xd_0__inst_i19_107 ;
wire Xd_0__inst_i19_109_sumout ;
wire Xd_0__inst_i19_110 ;
wire Xd_0__inst_i19_111 ;
wire Xd_0__inst_mult_30_88 ;
wire Xd_0__inst_mult_30_89 ;
wire Xd_0__inst_mult_30_90 ;
wire Xd_0__inst_mult_31_88 ;
wire Xd_0__inst_mult_31_89 ;
wire Xd_0__inst_mult_31_90 ;
wire Xd_0__inst_mult_30_92 ;
wire Xd_0__inst_mult_30_93 ;
wire Xd_0__inst_mult_30_94 ;
wire Xd_0__inst_mult_31_92 ;
wire Xd_0__inst_mult_31_93 ;
wire Xd_0__inst_mult_31_94 ;
wire Xd_0__inst_mult_28_49 ;
wire Xd_0__inst_mult_28_50 ;
wire Xd_0__inst_mult_28_51 ;
wire Xd_0__inst_mult_29_49 ;
wire Xd_0__inst_mult_29_50 ;
wire Xd_0__inst_mult_29_51 ;
wire Xd_0__inst_mult_26_49 ;
wire Xd_0__inst_mult_26_50 ;
wire Xd_0__inst_mult_26_51 ;
wire Xd_0__inst_mult_27_49 ;
wire Xd_0__inst_mult_27_50 ;
wire Xd_0__inst_mult_27_51 ;
wire Xd_0__inst_mult_24_49 ;
wire Xd_0__inst_mult_24_50 ;
wire Xd_0__inst_mult_24_51 ;
wire Xd_0__inst_mult_25_49 ;
wire Xd_0__inst_mult_25_50 ;
wire Xd_0__inst_mult_25_51 ;
wire Xd_0__inst_mult_22_49 ;
wire Xd_0__inst_mult_22_50 ;
wire Xd_0__inst_mult_22_51 ;
wire Xd_0__inst_mult_23_49 ;
wire Xd_0__inst_mult_23_50 ;
wire Xd_0__inst_mult_23_51 ;
wire Xd_0__inst_mult_20_49 ;
wire Xd_0__inst_mult_20_50 ;
wire Xd_0__inst_mult_20_51 ;
wire Xd_0__inst_mult_21_49 ;
wire Xd_0__inst_mult_21_50 ;
wire Xd_0__inst_mult_21_51 ;
wire Xd_0__inst_mult_18_49 ;
wire Xd_0__inst_mult_18_50 ;
wire Xd_0__inst_mult_18_51 ;
wire Xd_0__inst_mult_19_49 ;
wire Xd_0__inst_mult_19_50 ;
wire Xd_0__inst_mult_19_51 ;
wire Xd_0__inst_mult_30_97 ;
wire Xd_0__inst_mult_30_98 ;
wire Xd_0__inst_mult_31_97 ;
wire Xd_0__inst_mult_31_98 ;
wire Xd_0__inst_mult_16_49 ;
wire Xd_0__inst_mult_16_50 ;
wire Xd_0__inst_mult_16_51 ;
wire Xd_0__inst_mult_17_49 ;
wire Xd_0__inst_mult_17_50 ;
wire Xd_0__inst_mult_17_51 ;
wire Xd_0__inst_mult_14_49 ;
wire Xd_0__inst_mult_14_50 ;
wire Xd_0__inst_mult_14_51 ;
wire Xd_0__inst_mult_15_49 ;
wire Xd_0__inst_mult_15_50 ;
wire Xd_0__inst_mult_15_51 ;
wire Xd_0__inst_mult_12_49 ;
wire Xd_0__inst_mult_12_50 ;
wire Xd_0__inst_mult_12_51 ;
wire Xd_0__inst_mult_13_49 ;
wire Xd_0__inst_mult_13_50 ;
wire Xd_0__inst_mult_13_51 ;
wire Xd_0__inst_mult_10_49 ;
wire Xd_0__inst_mult_10_50 ;
wire Xd_0__inst_mult_10_51 ;
wire Xd_0__inst_mult_11_49 ;
wire Xd_0__inst_mult_11_50 ;
wire Xd_0__inst_mult_11_51 ;
wire Xd_0__inst_mult_8_49 ;
wire Xd_0__inst_mult_8_50 ;
wire Xd_0__inst_mult_8_51 ;
wire Xd_0__inst_mult_9_49 ;
wire Xd_0__inst_mult_9_50 ;
wire Xd_0__inst_mult_9_51 ;
wire Xd_0__inst_mult_6_49 ;
wire Xd_0__inst_mult_6_50 ;
wire Xd_0__inst_mult_6_51 ;
wire Xd_0__inst_mult_7_49 ;
wire Xd_0__inst_mult_7_50 ;
wire Xd_0__inst_mult_7_51 ;
wire Xd_0__inst_mult_4_49 ;
wire Xd_0__inst_mult_4_50 ;
wire Xd_0__inst_mult_4_51 ;
wire Xd_0__inst_mult_5_49 ;
wire Xd_0__inst_mult_5_50 ;
wire Xd_0__inst_mult_5_51 ;
wire Xd_0__inst_mult_2_49 ;
wire Xd_0__inst_mult_2_50 ;
wire Xd_0__inst_mult_2_51 ;
wire Xd_0__inst_mult_3_49 ;
wire Xd_0__inst_mult_3_50 ;
wire Xd_0__inst_mult_3_51 ;
wire Xd_0__inst_mult_0_49 ;
wire Xd_0__inst_mult_0_50 ;
wire Xd_0__inst_mult_0_51 ;
wire Xd_0__inst_mult_1_49 ;
wire Xd_0__inst_mult_1_50 ;
wire Xd_0__inst_mult_1_51 ;
wire Xd_0__inst_mult_28_53 ;
wire Xd_0__inst_mult_28_54 ;
wire Xd_0__inst_mult_28_55 ;
wire Xd_0__inst_mult_29_53 ;
wire Xd_0__inst_mult_29_54 ;
wire Xd_0__inst_mult_29_55 ;
wire Xd_0__inst_mult_26_53 ;
wire Xd_0__inst_mult_26_54 ;
wire Xd_0__inst_mult_26_55 ;
wire Xd_0__inst_mult_27_53 ;
wire Xd_0__inst_mult_27_54 ;
wire Xd_0__inst_mult_27_55 ;
wire Xd_0__inst_mult_24_53 ;
wire Xd_0__inst_mult_24_54 ;
wire Xd_0__inst_mult_24_55 ;
wire Xd_0__inst_mult_25_53 ;
wire Xd_0__inst_mult_25_54 ;
wire Xd_0__inst_mult_25_55 ;
wire Xd_0__inst_mult_22_53 ;
wire Xd_0__inst_mult_22_54 ;
wire Xd_0__inst_mult_22_55 ;
wire Xd_0__inst_mult_23_53 ;
wire Xd_0__inst_mult_23_54 ;
wire Xd_0__inst_mult_23_55 ;
wire Xd_0__inst_mult_20_53 ;
wire Xd_0__inst_mult_20_54 ;
wire Xd_0__inst_mult_20_55 ;
wire Xd_0__inst_mult_21_53 ;
wire Xd_0__inst_mult_21_54 ;
wire Xd_0__inst_mult_21_55 ;
wire Xd_0__inst_mult_18_53 ;
wire Xd_0__inst_mult_18_54 ;
wire Xd_0__inst_mult_18_55 ;
wire Xd_0__inst_mult_19_53 ;
wire Xd_0__inst_mult_19_54 ;
wire Xd_0__inst_mult_19_55 ;
wire Xd_0__inst_mult_16_53 ;
wire Xd_0__inst_mult_16_54 ;
wire Xd_0__inst_mult_16_55 ;
wire Xd_0__inst_mult_17_53 ;
wire Xd_0__inst_mult_17_54 ;
wire Xd_0__inst_mult_17_55 ;
wire Xd_0__inst_mult_14_53 ;
wire Xd_0__inst_mult_14_54 ;
wire Xd_0__inst_mult_14_55 ;
wire Xd_0__inst_mult_15_53 ;
wire Xd_0__inst_mult_15_54 ;
wire Xd_0__inst_mult_15_55 ;
wire Xd_0__inst_mult_12_53 ;
wire Xd_0__inst_mult_12_54 ;
wire Xd_0__inst_mult_12_55 ;
wire Xd_0__inst_mult_13_53 ;
wire Xd_0__inst_mult_13_54 ;
wire Xd_0__inst_mult_13_55 ;
wire Xd_0__inst_mult_10_53 ;
wire Xd_0__inst_mult_10_54 ;
wire Xd_0__inst_mult_10_55 ;
wire Xd_0__inst_mult_11_53 ;
wire Xd_0__inst_mult_11_54 ;
wire Xd_0__inst_mult_11_55 ;
wire Xd_0__inst_mult_8_53 ;
wire Xd_0__inst_mult_8_54 ;
wire Xd_0__inst_mult_8_55 ;
wire Xd_0__inst_mult_9_53 ;
wire Xd_0__inst_mult_9_54 ;
wire Xd_0__inst_mult_9_55 ;
wire Xd_0__inst_mult_6_53 ;
wire Xd_0__inst_mult_6_54 ;
wire Xd_0__inst_mult_6_55 ;
wire Xd_0__inst_mult_7_53 ;
wire Xd_0__inst_mult_7_54 ;
wire Xd_0__inst_mult_7_55 ;
wire Xd_0__inst_mult_4_53 ;
wire Xd_0__inst_mult_4_54 ;
wire Xd_0__inst_mult_4_55 ;
wire Xd_0__inst_mult_5_53 ;
wire Xd_0__inst_mult_5_54 ;
wire Xd_0__inst_mult_5_55 ;
wire Xd_0__inst_mult_2_53 ;
wire Xd_0__inst_mult_2_54 ;
wire Xd_0__inst_mult_2_55 ;
wire Xd_0__inst_mult_3_53 ;
wire Xd_0__inst_mult_3_54 ;
wire Xd_0__inst_mult_3_55 ;
wire Xd_0__inst_mult_0_53 ;
wire Xd_0__inst_mult_0_54 ;
wire Xd_0__inst_mult_0_55 ;
wire Xd_0__inst_mult_1_53 ;
wire Xd_0__inst_mult_1_54 ;
wire Xd_0__inst_mult_1_55 ;
wire Xd_0__inst_mult_28_56 ;
wire Xd_0__inst_mult_28_57 ;
wire Xd_0__inst_mult_28_58 ;
wire Xd_0__inst_mult_29_56 ;
wire Xd_0__inst_mult_29_57 ;
wire Xd_0__inst_mult_29_58 ;
wire Xd_0__inst_mult_26_56 ;
wire Xd_0__inst_mult_26_57 ;
wire Xd_0__inst_mult_26_58 ;
wire Xd_0__inst_mult_27_56 ;
wire Xd_0__inst_mult_27_57 ;
wire Xd_0__inst_mult_27_58 ;
wire Xd_0__inst_mult_24_56 ;
wire Xd_0__inst_mult_24_57 ;
wire Xd_0__inst_mult_24_58 ;
wire Xd_0__inst_mult_25_56 ;
wire Xd_0__inst_mult_25_57 ;
wire Xd_0__inst_mult_25_58 ;
wire Xd_0__inst_mult_22_56 ;
wire Xd_0__inst_mult_22_57 ;
wire Xd_0__inst_mult_22_58 ;
wire Xd_0__inst_mult_23_56 ;
wire Xd_0__inst_mult_23_57 ;
wire Xd_0__inst_mult_23_58 ;
wire Xd_0__inst_mult_20_56 ;
wire Xd_0__inst_mult_20_57 ;
wire Xd_0__inst_mult_20_58 ;
wire Xd_0__inst_mult_21_56 ;
wire Xd_0__inst_mult_21_57 ;
wire Xd_0__inst_mult_21_58 ;
wire Xd_0__inst_mult_18_56 ;
wire Xd_0__inst_mult_18_57 ;
wire Xd_0__inst_mult_18_58 ;
wire Xd_0__inst_mult_19_56 ;
wire Xd_0__inst_mult_19_57 ;
wire Xd_0__inst_mult_19_58 ;
wire Xd_0__inst_mult_16_56 ;
wire Xd_0__inst_mult_16_57 ;
wire Xd_0__inst_mult_16_58 ;
wire Xd_0__inst_mult_17_56 ;
wire Xd_0__inst_mult_17_57 ;
wire Xd_0__inst_mult_17_58 ;
wire Xd_0__inst_mult_14_56 ;
wire Xd_0__inst_mult_14_57 ;
wire Xd_0__inst_mult_14_58 ;
wire Xd_0__inst_mult_15_56 ;
wire Xd_0__inst_mult_15_57 ;
wire Xd_0__inst_mult_15_58 ;
wire Xd_0__inst_mult_12_56 ;
wire Xd_0__inst_mult_12_57 ;
wire Xd_0__inst_mult_12_58 ;
wire Xd_0__inst_mult_13_56 ;
wire Xd_0__inst_mult_13_57 ;
wire Xd_0__inst_mult_13_58 ;
wire Xd_0__inst_mult_10_56 ;
wire Xd_0__inst_mult_10_57 ;
wire Xd_0__inst_mult_10_58 ;
wire Xd_0__inst_mult_11_56 ;
wire Xd_0__inst_mult_11_57 ;
wire Xd_0__inst_mult_11_58 ;
wire Xd_0__inst_mult_8_56 ;
wire Xd_0__inst_mult_8_57 ;
wire Xd_0__inst_mult_8_58 ;
wire Xd_0__inst_mult_9_56 ;
wire Xd_0__inst_mult_9_57 ;
wire Xd_0__inst_mult_9_58 ;
wire Xd_0__inst_mult_6_56 ;
wire Xd_0__inst_mult_6_57 ;
wire Xd_0__inst_mult_6_58 ;
wire Xd_0__inst_mult_7_56 ;
wire Xd_0__inst_mult_7_57 ;
wire Xd_0__inst_mult_7_58 ;
wire Xd_0__inst_mult_4_56 ;
wire Xd_0__inst_mult_4_57 ;
wire Xd_0__inst_mult_4_58 ;
wire Xd_0__inst_mult_5_56 ;
wire Xd_0__inst_mult_5_57 ;
wire Xd_0__inst_mult_5_58 ;
wire Xd_0__inst_mult_2_56 ;
wire Xd_0__inst_mult_2_57 ;
wire Xd_0__inst_mult_2_58 ;
wire Xd_0__inst_mult_3_56 ;
wire Xd_0__inst_mult_3_57 ;
wire Xd_0__inst_mult_3_58 ;
wire Xd_0__inst_mult_0_56 ;
wire Xd_0__inst_mult_0_57 ;
wire Xd_0__inst_mult_0_58 ;
wire Xd_0__inst_mult_1_56 ;
wire Xd_0__inst_mult_1_57 ;
wire Xd_0__inst_mult_1_58 ;
wire Xd_0__inst_mult_28_60 ;
wire Xd_0__inst_mult_28_61 ;
wire Xd_0__inst_mult_28_62 ;
wire Xd_0__inst_mult_29_60 ;
wire Xd_0__inst_mult_29_61 ;
wire Xd_0__inst_mult_29_62 ;
wire Xd_0__inst_mult_26_60 ;
wire Xd_0__inst_mult_26_61 ;
wire Xd_0__inst_mult_26_62 ;
wire Xd_0__inst_mult_27_60 ;
wire Xd_0__inst_mult_27_61 ;
wire Xd_0__inst_mult_27_62 ;
wire Xd_0__inst_mult_24_60 ;
wire Xd_0__inst_mult_24_61 ;
wire Xd_0__inst_mult_24_62 ;
wire Xd_0__inst_mult_25_60 ;
wire Xd_0__inst_mult_25_61 ;
wire Xd_0__inst_mult_25_62 ;
wire Xd_0__inst_mult_22_60 ;
wire Xd_0__inst_mult_22_61 ;
wire Xd_0__inst_mult_22_62 ;
wire Xd_0__inst_mult_23_60 ;
wire Xd_0__inst_mult_23_61 ;
wire Xd_0__inst_mult_23_62 ;
wire Xd_0__inst_mult_20_60 ;
wire Xd_0__inst_mult_20_61 ;
wire Xd_0__inst_mult_20_62 ;
wire Xd_0__inst_mult_21_60 ;
wire Xd_0__inst_mult_21_61 ;
wire Xd_0__inst_mult_21_62 ;
wire Xd_0__inst_mult_18_60 ;
wire Xd_0__inst_mult_18_61 ;
wire Xd_0__inst_mult_18_62 ;
wire Xd_0__inst_mult_19_60 ;
wire Xd_0__inst_mult_19_61 ;
wire Xd_0__inst_mult_19_62 ;
wire Xd_0__inst_mult_16_60 ;
wire Xd_0__inst_mult_16_61 ;
wire Xd_0__inst_mult_16_62 ;
wire Xd_0__inst_mult_17_60 ;
wire Xd_0__inst_mult_17_61 ;
wire Xd_0__inst_mult_17_62 ;
wire Xd_0__inst_mult_14_60 ;
wire Xd_0__inst_mult_14_61 ;
wire Xd_0__inst_mult_14_62 ;
wire Xd_0__inst_mult_15_60 ;
wire Xd_0__inst_mult_15_61 ;
wire Xd_0__inst_mult_15_62 ;
wire Xd_0__inst_mult_12_60 ;
wire Xd_0__inst_mult_12_61 ;
wire Xd_0__inst_mult_12_62 ;
wire Xd_0__inst_mult_13_60 ;
wire Xd_0__inst_mult_13_61 ;
wire Xd_0__inst_mult_13_62 ;
wire Xd_0__inst_mult_10_60 ;
wire Xd_0__inst_mult_10_61 ;
wire Xd_0__inst_mult_10_62 ;
wire Xd_0__inst_mult_11_60 ;
wire Xd_0__inst_mult_11_61 ;
wire Xd_0__inst_mult_11_62 ;
wire Xd_0__inst_mult_8_60 ;
wire Xd_0__inst_mult_8_61 ;
wire Xd_0__inst_mult_8_62 ;
wire Xd_0__inst_mult_9_60 ;
wire Xd_0__inst_mult_9_61 ;
wire Xd_0__inst_mult_9_62 ;
wire Xd_0__inst_mult_6_60 ;
wire Xd_0__inst_mult_6_61 ;
wire Xd_0__inst_mult_6_62 ;
wire Xd_0__inst_mult_7_60 ;
wire Xd_0__inst_mult_7_61 ;
wire Xd_0__inst_mult_7_62 ;
wire Xd_0__inst_mult_4_60 ;
wire Xd_0__inst_mult_4_61 ;
wire Xd_0__inst_mult_4_62 ;
wire Xd_0__inst_mult_5_60 ;
wire Xd_0__inst_mult_5_61 ;
wire Xd_0__inst_mult_5_62 ;
wire Xd_0__inst_mult_2_60 ;
wire Xd_0__inst_mult_2_61 ;
wire Xd_0__inst_mult_2_62 ;
wire Xd_0__inst_mult_3_60 ;
wire Xd_0__inst_mult_3_61 ;
wire Xd_0__inst_mult_3_62 ;
wire Xd_0__inst_mult_0_60 ;
wire Xd_0__inst_mult_0_61 ;
wire Xd_0__inst_mult_0_62 ;
wire Xd_0__inst_mult_1_60 ;
wire Xd_0__inst_mult_1_61 ;
wire Xd_0__inst_mult_1_62 ;
wire Xd_0__inst_mult_28_64 ;
wire Xd_0__inst_mult_28_65 ;
wire Xd_0__inst_mult_28_66 ;
wire Xd_0__inst_mult_29_64 ;
wire Xd_0__inst_mult_29_65 ;
wire Xd_0__inst_mult_29_66 ;
wire Xd_0__inst_mult_26_64 ;
wire Xd_0__inst_mult_26_65 ;
wire Xd_0__inst_mult_26_66 ;
wire Xd_0__inst_mult_27_64 ;
wire Xd_0__inst_mult_27_65 ;
wire Xd_0__inst_mult_27_66 ;
wire Xd_0__inst_mult_24_64 ;
wire Xd_0__inst_mult_24_65 ;
wire Xd_0__inst_mult_24_66 ;
wire Xd_0__inst_mult_25_64 ;
wire Xd_0__inst_mult_25_65 ;
wire Xd_0__inst_mult_25_66 ;
wire Xd_0__inst_mult_22_64 ;
wire Xd_0__inst_mult_22_65 ;
wire Xd_0__inst_mult_22_66 ;
wire Xd_0__inst_mult_23_64 ;
wire Xd_0__inst_mult_23_65 ;
wire Xd_0__inst_mult_23_66 ;
wire Xd_0__inst_mult_20_64 ;
wire Xd_0__inst_mult_20_65 ;
wire Xd_0__inst_mult_20_66 ;
wire Xd_0__inst_mult_21_64 ;
wire Xd_0__inst_mult_21_65 ;
wire Xd_0__inst_mult_21_66 ;
wire Xd_0__inst_mult_18_64 ;
wire Xd_0__inst_mult_18_65 ;
wire Xd_0__inst_mult_18_66 ;
wire Xd_0__inst_mult_19_64 ;
wire Xd_0__inst_mult_19_65 ;
wire Xd_0__inst_mult_19_66 ;
wire Xd_0__inst_mult_16_64 ;
wire Xd_0__inst_mult_16_65 ;
wire Xd_0__inst_mult_16_66 ;
wire Xd_0__inst_mult_17_64 ;
wire Xd_0__inst_mult_17_65 ;
wire Xd_0__inst_mult_17_66 ;
wire Xd_0__inst_mult_14_64 ;
wire Xd_0__inst_mult_14_65 ;
wire Xd_0__inst_mult_14_66 ;
wire Xd_0__inst_mult_15_64 ;
wire Xd_0__inst_mult_15_65 ;
wire Xd_0__inst_mult_15_66 ;
wire Xd_0__inst_mult_12_64 ;
wire Xd_0__inst_mult_12_65 ;
wire Xd_0__inst_mult_12_66 ;
wire Xd_0__inst_mult_13_64 ;
wire Xd_0__inst_mult_13_65 ;
wire Xd_0__inst_mult_13_66 ;
wire Xd_0__inst_mult_10_64 ;
wire Xd_0__inst_mult_10_65 ;
wire Xd_0__inst_mult_10_66 ;
wire Xd_0__inst_mult_11_64 ;
wire Xd_0__inst_mult_11_65 ;
wire Xd_0__inst_mult_11_66 ;
wire Xd_0__inst_mult_8_64 ;
wire Xd_0__inst_mult_8_65 ;
wire Xd_0__inst_mult_8_66 ;
wire Xd_0__inst_mult_9_64 ;
wire Xd_0__inst_mult_9_65 ;
wire Xd_0__inst_mult_9_66 ;
wire Xd_0__inst_mult_6_64 ;
wire Xd_0__inst_mult_6_65 ;
wire Xd_0__inst_mult_6_66 ;
wire Xd_0__inst_mult_7_64 ;
wire Xd_0__inst_mult_7_65 ;
wire Xd_0__inst_mult_7_66 ;
wire Xd_0__inst_mult_4_64 ;
wire Xd_0__inst_mult_4_65 ;
wire Xd_0__inst_mult_4_66 ;
wire Xd_0__inst_mult_5_64 ;
wire Xd_0__inst_mult_5_65 ;
wire Xd_0__inst_mult_5_66 ;
wire Xd_0__inst_mult_2_64 ;
wire Xd_0__inst_mult_2_65 ;
wire Xd_0__inst_mult_2_66 ;
wire Xd_0__inst_mult_3_64 ;
wire Xd_0__inst_mult_3_65 ;
wire Xd_0__inst_mult_3_66 ;
wire Xd_0__inst_mult_0_64 ;
wire Xd_0__inst_mult_0_65 ;
wire Xd_0__inst_mult_0_66 ;
wire Xd_0__inst_mult_1_64 ;
wire Xd_0__inst_mult_1_65 ;
wire Xd_0__inst_mult_1_66 ;
wire Xd_0__inst_mult_28_68 ;
wire Xd_0__inst_mult_28_69 ;
wire Xd_0__inst_mult_28_70 ;
wire Xd_0__inst_mult_29_68 ;
wire Xd_0__inst_mult_29_69 ;
wire Xd_0__inst_mult_29_70 ;
wire Xd_0__inst_mult_26_68 ;
wire Xd_0__inst_mult_26_69 ;
wire Xd_0__inst_mult_26_70 ;
wire Xd_0__inst_mult_27_68 ;
wire Xd_0__inst_mult_27_69 ;
wire Xd_0__inst_mult_27_70 ;
wire Xd_0__inst_mult_24_68 ;
wire Xd_0__inst_mult_24_69 ;
wire Xd_0__inst_mult_24_70 ;
wire Xd_0__inst_mult_25_68 ;
wire Xd_0__inst_mult_25_69 ;
wire Xd_0__inst_mult_25_70 ;
wire Xd_0__inst_mult_22_68 ;
wire Xd_0__inst_mult_22_69 ;
wire Xd_0__inst_mult_22_70 ;
wire Xd_0__inst_mult_23_68 ;
wire Xd_0__inst_mult_23_69 ;
wire Xd_0__inst_mult_23_70 ;
wire Xd_0__inst_mult_20_68 ;
wire Xd_0__inst_mult_20_69 ;
wire Xd_0__inst_mult_20_70 ;
wire Xd_0__inst_mult_21_68 ;
wire Xd_0__inst_mult_21_69 ;
wire Xd_0__inst_mult_21_70 ;
wire Xd_0__inst_mult_18_68 ;
wire Xd_0__inst_mult_18_69 ;
wire Xd_0__inst_mult_18_70 ;
wire Xd_0__inst_mult_19_68 ;
wire Xd_0__inst_mult_19_69 ;
wire Xd_0__inst_mult_19_70 ;
wire Xd_0__inst_mult_16_68 ;
wire Xd_0__inst_mult_16_69 ;
wire Xd_0__inst_mult_16_70 ;
wire Xd_0__inst_mult_17_68 ;
wire Xd_0__inst_mult_17_69 ;
wire Xd_0__inst_mult_17_70 ;
wire Xd_0__inst_mult_14_68 ;
wire Xd_0__inst_mult_14_69 ;
wire Xd_0__inst_mult_14_70 ;
wire Xd_0__inst_mult_15_68 ;
wire Xd_0__inst_mult_15_69 ;
wire Xd_0__inst_mult_15_70 ;
wire Xd_0__inst_mult_12_68 ;
wire Xd_0__inst_mult_12_69 ;
wire Xd_0__inst_mult_12_70 ;
wire Xd_0__inst_mult_13_68 ;
wire Xd_0__inst_mult_13_69 ;
wire Xd_0__inst_mult_13_70 ;
wire Xd_0__inst_mult_10_68 ;
wire Xd_0__inst_mult_10_69 ;
wire Xd_0__inst_mult_10_70 ;
wire Xd_0__inst_mult_11_68 ;
wire Xd_0__inst_mult_11_69 ;
wire Xd_0__inst_mult_11_70 ;
wire Xd_0__inst_mult_8_68 ;
wire Xd_0__inst_mult_8_69 ;
wire Xd_0__inst_mult_8_70 ;
wire Xd_0__inst_mult_9_68 ;
wire Xd_0__inst_mult_9_69 ;
wire Xd_0__inst_mult_9_70 ;
wire Xd_0__inst_mult_6_68 ;
wire Xd_0__inst_mult_6_69 ;
wire Xd_0__inst_mult_6_70 ;
wire Xd_0__inst_mult_7_68 ;
wire Xd_0__inst_mult_7_69 ;
wire Xd_0__inst_mult_7_70 ;
wire Xd_0__inst_mult_4_68 ;
wire Xd_0__inst_mult_4_69 ;
wire Xd_0__inst_mult_4_70 ;
wire Xd_0__inst_mult_5_68 ;
wire Xd_0__inst_mult_5_69 ;
wire Xd_0__inst_mult_5_70 ;
wire Xd_0__inst_mult_2_68 ;
wire Xd_0__inst_mult_2_69 ;
wire Xd_0__inst_mult_2_70 ;
wire Xd_0__inst_mult_3_68 ;
wire Xd_0__inst_mult_3_69 ;
wire Xd_0__inst_mult_3_70 ;
wire Xd_0__inst_mult_0_68 ;
wire Xd_0__inst_mult_0_69 ;
wire Xd_0__inst_mult_0_70 ;
wire Xd_0__inst_mult_1_68 ;
wire Xd_0__inst_mult_1_69 ;
wire Xd_0__inst_mult_1_70 ;
wire Xd_0__inst_mult_28_72 ;
wire Xd_0__inst_mult_28_73 ;
wire Xd_0__inst_mult_28_74 ;
wire Xd_0__inst_mult_29_72 ;
wire Xd_0__inst_mult_29_73 ;
wire Xd_0__inst_mult_29_74 ;
wire Xd_0__inst_mult_26_72 ;
wire Xd_0__inst_mult_26_73 ;
wire Xd_0__inst_mult_26_74 ;
wire Xd_0__inst_mult_27_72 ;
wire Xd_0__inst_mult_27_73 ;
wire Xd_0__inst_mult_27_74 ;
wire Xd_0__inst_mult_24_72 ;
wire Xd_0__inst_mult_24_73 ;
wire Xd_0__inst_mult_24_74 ;
wire Xd_0__inst_mult_25_72 ;
wire Xd_0__inst_mult_25_73 ;
wire Xd_0__inst_mult_25_74 ;
wire Xd_0__inst_mult_22_72 ;
wire Xd_0__inst_mult_22_73 ;
wire Xd_0__inst_mult_22_74 ;
wire Xd_0__inst_mult_23_72 ;
wire Xd_0__inst_mult_23_73 ;
wire Xd_0__inst_mult_23_74 ;
wire Xd_0__inst_mult_20_72 ;
wire Xd_0__inst_mult_20_73 ;
wire Xd_0__inst_mult_20_74 ;
wire Xd_0__inst_mult_21_72 ;
wire Xd_0__inst_mult_21_73 ;
wire Xd_0__inst_mult_21_74 ;
wire Xd_0__inst_mult_18_72 ;
wire Xd_0__inst_mult_18_73 ;
wire Xd_0__inst_mult_18_74 ;
wire Xd_0__inst_mult_19_72 ;
wire Xd_0__inst_mult_19_73 ;
wire Xd_0__inst_mult_19_74 ;
wire Xd_0__inst_mult_16_72 ;
wire Xd_0__inst_mult_16_73 ;
wire Xd_0__inst_mult_16_74 ;
wire Xd_0__inst_mult_17_72 ;
wire Xd_0__inst_mult_17_73 ;
wire Xd_0__inst_mult_17_74 ;
wire Xd_0__inst_mult_14_72 ;
wire Xd_0__inst_mult_14_73 ;
wire Xd_0__inst_mult_14_74 ;
wire Xd_0__inst_mult_15_72 ;
wire Xd_0__inst_mult_15_73 ;
wire Xd_0__inst_mult_15_74 ;
wire Xd_0__inst_mult_12_72 ;
wire Xd_0__inst_mult_12_73 ;
wire Xd_0__inst_mult_12_74 ;
wire Xd_0__inst_mult_13_72 ;
wire Xd_0__inst_mult_13_73 ;
wire Xd_0__inst_mult_13_74 ;
wire Xd_0__inst_mult_10_72 ;
wire Xd_0__inst_mult_10_73 ;
wire Xd_0__inst_mult_10_74 ;
wire Xd_0__inst_mult_11_72 ;
wire Xd_0__inst_mult_11_73 ;
wire Xd_0__inst_mult_11_74 ;
wire Xd_0__inst_mult_8_72 ;
wire Xd_0__inst_mult_8_73 ;
wire Xd_0__inst_mult_8_74 ;
wire Xd_0__inst_mult_9_72 ;
wire Xd_0__inst_mult_9_73 ;
wire Xd_0__inst_mult_9_74 ;
wire Xd_0__inst_mult_6_72 ;
wire Xd_0__inst_mult_6_73 ;
wire Xd_0__inst_mult_6_74 ;
wire Xd_0__inst_mult_7_72 ;
wire Xd_0__inst_mult_7_73 ;
wire Xd_0__inst_mult_7_74 ;
wire Xd_0__inst_mult_4_72 ;
wire Xd_0__inst_mult_4_73 ;
wire Xd_0__inst_mult_4_74 ;
wire Xd_0__inst_mult_5_72 ;
wire Xd_0__inst_mult_5_73 ;
wire Xd_0__inst_mult_5_74 ;
wire Xd_0__inst_mult_2_72 ;
wire Xd_0__inst_mult_2_73 ;
wire Xd_0__inst_mult_2_74 ;
wire Xd_0__inst_mult_3_72 ;
wire Xd_0__inst_mult_3_73 ;
wire Xd_0__inst_mult_3_74 ;
wire Xd_0__inst_mult_0_72 ;
wire Xd_0__inst_mult_0_73 ;
wire Xd_0__inst_mult_0_74 ;
wire Xd_0__inst_mult_1_72 ;
wire Xd_0__inst_mult_1_73 ;
wire Xd_0__inst_mult_1_74 ;
wire Xd_0__inst_mult_28_76 ;
wire Xd_0__inst_mult_28_77 ;
wire Xd_0__inst_mult_28_78 ;
wire Xd_0__inst_mult_29_76 ;
wire Xd_0__inst_mult_29_77 ;
wire Xd_0__inst_mult_29_78 ;
wire Xd_0__inst_mult_26_76 ;
wire Xd_0__inst_mult_26_77 ;
wire Xd_0__inst_mult_26_78 ;
wire Xd_0__inst_mult_27_76 ;
wire Xd_0__inst_mult_27_77 ;
wire Xd_0__inst_mult_27_78 ;
wire Xd_0__inst_mult_24_76 ;
wire Xd_0__inst_mult_24_77 ;
wire Xd_0__inst_mult_24_78 ;
wire Xd_0__inst_mult_25_76 ;
wire Xd_0__inst_mult_25_77 ;
wire Xd_0__inst_mult_25_78 ;
wire Xd_0__inst_mult_22_76 ;
wire Xd_0__inst_mult_22_77 ;
wire Xd_0__inst_mult_22_78 ;
wire Xd_0__inst_mult_23_76 ;
wire Xd_0__inst_mult_23_77 ;
wire Xd_0__inst_mult_23_78 ;
wire Xd_0__inst_mult_20_76 ;
wire Xd_0__inst_mult_20_77 ;
wire Xd_0__inst_mult_20_78 ;
wire Xd_0__inst_mult_21_76 ;
wire Xd_0__inst_mult_21_77 ;
wire Xd_0__inst_mult_21_78 ;
wire Xd_0__inst_mult_18_76 ;
wire Xd_0__inst_mult_18_77 ;
wire Xd_0__inst_mult_18_78 ;
wire Xd_0__inst_mult_19_76 ;
wire Xd_0__inst_mult_19_77 ;
wire Xd_0__inst_mult_19_78 ;
wire Xd_0__inst_mult_16_76 ;
wire Xd_0__inst_mult_16_77 ;
wire Xd_0__inst_mult_16_78 ;
wire Xd_0__inst_mult_17_76 ;
wire Xd_0__inst_mult_17_77 ;
wire Xd_0__inst_mult_17_78 ;
wire Xd_0__inst_mult_14_76 ;
wire Xd_0__inst_mult_14_77 ;
wire Xd_0__inst_mult_14_78 ;
wire Xd_0__inst_mult_15_76 ;
wire Xd_0__inst_mult_15_77 ;
wire Xd_0__inst_mult_15_78 ;
wire Xd_0__inst_mult_12_76 ;
wire Xd_0__inst_mult_12_77 ;
wire Xd_0__inst_mult_12_78 ;
wire Xd_0__inst_mult_13_76 ;
wire Xd_0__inst_mult_13_77 ;
wire Xd_0__inst_mult_13_78 ;
wire Xd_0__inst_mult_10_76 ;
wire Xd_0__inst_mult_10_77 ;
wire Xd_0__inst_mult_10_78 ;
wire Xd_0__inst_mult_11_76 ;
wire Xd_0__inst_mult_11_77 ;
wire Xd_0__inst_mult_11_78 ;
wire Xd_0__inst_mult_8_76 ;
wire Xd_0__inst_mult_8_77 ;
wire Xd_0__inst_mult_8_78 ;
wire Xd_0__inst_mult_9_76 ;
wire Xd_0__inst_mult_9_77 ;
wire Xd_0__inst_mult_9_78 ;
wire Xd_0__inst_mult_6_76 ;
wire Xd_0__inst_mult_6_77 ;
wire Xd_0__inst_mult_6_78 ;
wire Xd_0__inst_mult_7_76 ;
wire Xd_0__inst_mult_7_77 ;
wire Xd_0__inst_mult_7_78 ;
wire Xd_0__inst_mult_4_76 ;
wire Xd_0__inst_mult_4_77 ;
wire Xd_0__inst_mult_4_78 ;
wire Xd_0__inst_mult_5_76 ;
wire Xd_0__inst_mult_5_77 ;
wire Xd_0__inst_mult_5_78 ;
wire Xd_0__inst_mult_2_76 ;
wire Xd_0__inst_mult_2_77 ;
wire Xd_0__inst_mult_2_78 ;
wire Xd_0__inst_mult_3_76 ;
wire Xd_0__inst_mult_3_77 ;
wire Xd_0__inst_mult_3_78 ;
wire Xd_0__inst_mult_0_76 ;
wire Xd_0__inst_mult_0_77 ;
wire Xd_0__inst_mult_0_78 ;
wire Xd_0__inst_mult_1_76 ;
wire Xd_0__inst_mult_1_77 ;
wire Xd_0__inst_mult_1_78 ;
wire Xd_0__inst_mult_28_80 ;
wire Xd_0__inst_mult_29_80 ;
wire Xd_0__inst_mult_29_81 ;
wire Xd_0__inst_mult_29_82 ;
wire Xd_0__inst_mult_26_80 ;
wire Xd_0__inst_mult_27_80 ;
wire Xd_0__inst_mult_27_81 ;
wire Xd_0__inst_mult_27_82 ;
wire Xd_0__inst_mult_24_80 ;
wire Xd_0__inst_mult_25_80 ;
wire Xd_0__inst_mult_25_81 ;
wire Xd_0__inst_mult_25_82 ;
wire Xd_0__inst_mult_22_80 ;
wire Xd_0__inst_mult_23_80 ;
wire Xd_0__inst_mult_23_81 ;
wire Xd_0__inst_mult_23_82 ;
wire Xd_0__inst_mult_20_80 ;
wire Xd_0__inst_mult_21_80 ;
wire Xd_0__inst_mult_21_81 ;
wire Xd_0__inst_mult_21_82 ;
wire Xd_0__inst_mult_18_80 ;
wire Xd_0__inst_mult_19_80 ;
wire Xd_0__inst_mult_19_81 ;
wire Xd_0__inst_mult_19_82 ;
wire Xd_0__inst_mult_16_80 ;
wire Xd_0__inst_mult_16_81 ;
wire Xd_0__inst_mult_16_82 ;
wire Xd_0__inst_mult_17_80 ;
wire Xd_0__inst_mult_17_81 ;
wire Xd_0__inst_mult_17_82 ;
wire Xd_0__inst_mult_14_80 ;
wire Xd_0__inst_mult_15_80 ;
wire Xd_0__inst_mult_15_81 ;
wire Xd_0__inst_mult_15_82 ;
wire Xd_0__inst_mult_12_80 ;
wire Xd_0__inst_mult_13_80 ;
wire Xd_0__inst_mult_13_81 ;
wire Xd_0__inst_mult_13_82 ;
wire Xd_0__inst_mult_10_80 ;
wire Xd_0__inst_mult_11_80 ;
wire Xd_0__inst_mult_8_80 ;
wire Xd_0__inst_mult_8_81 ;
wire Xd_0__inst_mult_8_82 ;
wire Xd_0__inst_mult_9_80 ;
wire Xd_0__inst_mult_6_80 ;
wire Xd_0__inst_mult_6_81 ;
wire Xd_0__inst_mult_6_82 ;
wire Xd_0__inst_mult_7_80 ;
wire Xd_0__inst_mult_4_80 ;
wire Xd_0__inst_mult_4_81 ;
wire Xd_0__inst_mult_4_82 ;
wire Xd_0__inst_mult_5_80 ;
wire Xd_0__inst_mult_2_80 ;
wire Xd_0__inst_mult_2_81 ;
wire Xd_0__inst_mult_2_82 ;
wire Xd_0__inst_mult_3_80 ;
wire Xd_0__inst_mult_0_80 ;
wire Xd_0__inst_mult_0_81 ;
wire Xd_0__inst_mult_0_82 ;
wire Xd_0__inst_mult_1_80 ;
wire Xd_0__inst_mult_28_84 ;
wire Xd_0__inst_mult_28_85 ;
wire Xd_0__inst_mult_28_86 ;
wire Xd_0__inst_mult_29_84 ;
wire Xd_0__inst_mult_29_85 ;
wire Xd_0__inst_mult_29_86 ;
wire Xd_0__inst_mult_26_84 ;
wire Xd_0__inst_mult_26_85 ;
wire Xd_0__inst_mult_26_86 ;
wire Xd_0__inst_mult_27_84 ;
wire Xd_0__inst_mult_27_85 ;
wire Xd_0__inst_mult_27_86 ;
wire Xd_0__inst_mult_24_84 ;
wire Xd_0__inst_mult_24_85 ;
wire Xd_0__inst_mult_24_86 ;
wire Xd_0__inst_mult_25_84 ;
wire Xd_0__inst_mult_25_85 ;
wire Xd_0__inst_mult_25_86 ;
wire Xd_0__inst_mult_22_84 ;
wire Xd_0__inst_mult_22_85 ;
wire Xd_0__inst_mult_22_86 ;
wire Xd_0__inst_mult_23_84 ;
wire Xd_0__inst_mult_23_85 ;
wire Xd_0__inst_mult_23_86 ;
wire Xd_0__inst_mult_20_84 ;
wire Xd_0__inst_mult_20_85 ;
wire Xd_0__inst_mult_20_86 ;
wire Xd_0__inst_mult_21_84 ;
wire Xd_0__inst_mult_21_85 ;
wire Xd_0__inst_mult_21_86 ;
wire Xd_0__inst_mult_18_84 ;
wire Xd_0__inst_mult_18_85 ;
wire Xd_0__inst_mult_18_86 ;
wire Xd_0__inst_mult_19_84 ;
wire Xd_0__inst_mult_19_85 ;
wire Xd_0__inst_mult_19_86 ;
wire Xd_0__inst_mult_25_88 ;
wire Xd_0__inst_mult_25_89 ;
wire Xd_0__inst_mult_25_90 ;
wire Xd_0__inst_mult_22_88 ;
wire Xd_0__inst_mult_22_89 ;
wire Xd_0__inst_mult_22_90 ;
wire Xd_0__inst_mult_16_84 ;
wire Xd_0__inst_mult_16_85 ;
wire Xd_0__inst_mult_16_86 ;
wire Xd_0__inst_mult_17_84 ;
wire Xd_0__inst_mult_17_85 ;
wire Xd_0__inst_mult_17_86 ;
wire Xd_0__inst_mult_14_84 ;
wire Xd_0__inst_mult_14_85 ;
wire Xd_0__inst_mult_14_86 ;
wire Xd_0__inst_mult_15_84 ;
wire Xd_0__inst_mult_15_85 ;
wire Xd_0__inst_mult_15_86 ;
wire Xd_0__inst_mult_12_84 ;
wire Xd_0__inst_mult_12_85 ;
wire Xd_0__inst_mult_12_86 ;
wire Xd_0__inst_mult_13_84 ;
wire Xd_0__inst_mult_13_85 ;
wire Xd_0__inst_mult_13_86 ;
wire Xd_0__inst_mult_10_84 ;
wire Xd_0__inst_mult_10_85 ;
wire Xd_0__inst_mult_10_86 ;
wire Xd_0__inst_mult_11_84 ;
wire Xd_0__inst_mult_11_85 ;
wire Xd_0__inst_mult_11_86 ;
wire Xd_0__inst_mult_8_84 ;
wire Xd_0__inst_mult_8_85 ;
wire Xd_0__inst_mult_8_86 ;
wire Xd_0__inst_mult_9_84 ;
wire Xd_0__inst_mult_9_85 ;
wire Xd_0__inst_mult_9_86 ;
wire Xd_0__inst_mult_6_84 ;
wire Xd_0__inst_mult_6_85 ;
wire Xd_0__inst_mult_6_86 ;
wire Xd_0__inst_mult_7_84 ;
wire Xd_0__inst_mult_7_85 ;
wire Xd_0__inst_mult_7_86 ;
wire Xd_0__inst_mult_4_84 ;
wire Xd_0__inst_mult_4_85 ;
wire Xd_0__inst_mult_4_86 ;
wire Xd_0__inst_mult_5_84 ;
wire Xd_0__inst_mult_5_85 ;
wire Xd_0__inst_mult_5_86 ;
wire Xd_0__inst_i19_113_sumout ;
wire Xd_0__inst_i19_114 ;
wire Xd_0__inst_i19_115 ;
wire Xd_0__inst_i19_117_sumout ;
wire Xd_0__inst_i19_118 ;
wire Xd_0__inst_i19_119 ;
wire Xd_0__inst_mult_2_84 ;
wire Xd_0__inst_mult_2_85 ;
wire Xd_0__inst_mult_2_86 ;
wire Xd_0__inst_mult_3_84 ;
wire Xd_0__inst_mult_3_85 ;
wire Xd_0__inst_mult_3_86 ;
wire Xd_0__inst_i19_121_sumout ;
wire Xd_0__inst_i19_122 ;
wire Xd_0__inst_i19_123 ;
wire Xd_0__inst_i19_125_sumout ;
wire Xd_0__inst_i19_126 ;
wire Xd_0__inst_i19_127 ;
wire Xd_0__inst_mult_0_84 ;
wire Xd_0__inst_mult_0_85 ;
wire Xd_0__inst_mult_0_86 ;
wire Xd_0__inst_mult_1_84 ;
wire Xd_0__inst_mult_1_85 ;
wire Xd_0__inst_mult_1_86 ;
wire Xd_0__inst_mult_28_88 ;
wire Xd_0__inst_mult_28_89 ;
wire Xd_0__inst_mult_28_90 ;
wire Xd_0__inst_mult_29_88 ;
wire Xd_0__inst_mult_29_89 ;
wire Xd_0__inst_mult_29_90 ;
wire Xd_0__inst_mult_26_88 ;
wire Xd_0__inst_mult_26_89 ;
wire Xd_0__inst_mult_26_90 ;
wire Xd_0__inst_mult_27_88 ;
wire Xd_0__inst_mult_27_89 ;
wire Xd_0__inst_mult_27_90 ;
wire Xd_0__inst_mult_24_88 ;
wire Xd_0__inst_mult_24_89 ;
wire Xd_0__inst_mult_24_90 ;
wire Xd_0__inst_mult_25_92 ;
wire Xd_0__inst_mult_25_93 ;
wire Xd_0__inst_mult_25_94 ;
wire Xd_0__inst_mult_22_92 ;
wire Xd_0__inst_mult_22_93 ;
wire Xd_0__inst_mult_22_94 ;
wire Xd_0__inst_mult_23_88 ;
wire Xd_0__inst_mult_23_89 ;
wire Xd_0__inst_mult_23_90 ;
wire Xd_0__inst_mult_20_88 ;
wire Xd_0__inst_mult_20_89 ;
wire Xd_0__inst_mult_20_90 ;
wire Xd_0__inst_mult_21_88 ;
wire Xd_0__inst_mult_21_89 ;
wire Xd_0__inst_mult_21_90 ;
wire Xd_0__inst_mult_18_88 ;
wire Xd_0__inst_mult_18_89 ;
wire Xd_0__inst_mult_18_90 ;
wire Xd_0__inst_mult_19_88 ;
wire Xd_0__inst_mult_19_89 ;
wire Xd_0__inst_mult_19_90 ;
wire Xd_0__inst_mult_16_88 ;
wire Xd_0__inst_mult_16_89 ;
wire Xd_0__inst_mult_16_90 ;
wire Xd_0__inst_mult_17_88 ;
wire Xd_0__inst_mult_17_89 ;
wire Xd_0__inst_mult_17_90 ;
wire Xd_0__inst_mult_14_88 ;
wire Xd_0__inst_mult_14_89 ;
wire Xd_0__inst_mult_14_90 ;
wire Xd_0__inst_mult_15_88 ;
wire Xd_0__inst_mult_15_89 ;
wire Xd_0__inst_mult_15_90 ;
wire Xd_0__inst_mult_12_88 ;
wire Xd_0__inst_mult_12_89 ;
wire Xd_0__inst_mult_12_90 ;
wire Xd_0__inst_mult_13_88 ;
wire Xd_0__inst_mult_13_89 ;
wire Xd_0__inst_mult_13_90 ;
wire Xd_0__inst_mult_10_88 ;
wire Xd_0__inst_mult_10_89 ;
wire Xd_0__inst_mult_10_90 ;
wire Xd_0__inst_mult_11_88 ;
wire Xd_0__inst_mult_11_89 ;
wire Xd_0__inst_mult_11_90 ;
wire Xd_0__inst_mult_8_88 ;
wire Xd_0__inst_mult_8_89 ;
wire Xd_0__inst_mult_8_90 ;
wire Xd_0__inst_mult_9_88 ;
wire Xd_0__inst_mult_9_89 ;
wire Xd_0__inst_mult_9_90 ;
wire Xd_0__inst_mult_6_88 ;
wire Xd_0__inst_mult_6_89 ;
wire Xd_0__inst_mult_6_90 ;
wire Xd_0__inst_mult_7_88 ;
wire Xd_0__inst_mult_7_89 ;
wire Xd_0__inst_mult_7_90 ;
wire Xd_0__inst_mult_4_88 ;
wire Xd_0__inst_mult_4_89 ;
wire Xd_0__inst_mult_4_90 ;
wire Xd_0__inst_mult_5_88 ;
wire Xd_0__inst_mult_5_89 ;
wire Xd_0__inst_mult_5_90 ;
wire Xd_0__inst_mult_2_88 ;
wire Xd_0__inst_mult_2_89 ;
wire Xd_0__inst_mult_2_90 ;
wire Xd_0__inst_mult_3_88 ;
wire Xd_0__inst_mult_3_89 ;
wire Xd_0__inst_mult_3_90 ;
wire Xd_0__inst_mult_0_88 ;
wire Xd_0__inst_mult_0_89 ;
wire Xd_0__inst_mult_0_90 ;
wire Xd_0__inst_mult_1_88 ;
wire Xd_0__inst_mult_1_89 ;
wire Xd_0__inst_mult_1_90 ;
wire Xd_0__inst_mult_28_92 ;
wire Xd_0__inst_mult_28_93 ;
wire Xd_0__inst_mult_28_94 ;
wire Xd_0__inst_mult_29_92 ;
wire Xd_0__inst_mult_29_93 ;
wire Xd_0__inst_mult_29_94 ;
wire Xd_0__inst_mult_26_92 ;
wire Xd_0__inst_mult_26_93 ;
wire Xd_0__inst_mult_26_94 ;
wire Xd_0__inst_mult_27_92 ;
wire Xd_0__inst_mult_27_93 ;
wire Xd_0__inst_mult_27_94 ;
wire Xd_0__inst_mult_24_92 ;
wire Xd_0__inst_mult_24_93 ;
wire Xd_0__inst_mult_24_94 ;
wire Xd_0__inst_mult_25_96 ;
wire Xd_0__inst_mult_25_97 ;
wire Xd_0__inst_mult_25_98 ;
wire Xd_0__inst_mult_22_96 ;
wire Xd_0__inst_mult_22_97 ;
wire Xd_0__inst_mult_22_98 ;
wire Xd_0__inst_mult_23_92 ;
wire Xd_0__inst_mult_23_93 ;
wire Xd_0__inst_mult_23_94 ;
wire Xd_0__inst_mult_20_92 ;
wire Xd_0__inst_mult_20_93 ;
wire Xd_0__inst_mult_20_94 ;
wire Xd_0__inst_mult_21_92 ;
wire Xd_0__inst_mult_21_93 ;
wire Xd_0__inst_mult_21_94 ;
wire Xd_0__inst_mult_18_92 ;
wire Xd_0__inst_mult_18_93 ;
wire Xd_0__inst_mult_18_94 ;
wire Xd_0__inst_mult_19_92 ;
wire Xd_0__inst_mult_19_93 ;
wire Xd_0__inst_mult_19_94 ;
wire Xd_0__inst_mult_16_92 ;
wire Xd_0__inst_mult_16_93 ;
wire Xd_0__inst_mult_16_94 ;
wire Xd_0__inst_mult_17_92 ;
wire Xd_0__inst_mult_17_93 ;
wire Xd_0__inst_mult_17_94 ;
wire Xd_0__inst_mult_14_92 ;
wire Xd_0__inst_mult_14_93 ;
wire Xd_0__inst_mult_14_94 ;
wire Xd_0__inst_mult_15_92 ;
wire Xd_0__inst_mult_15_93 ;
wire Xd_0__inst_mult_15_94 ;
wire Xd_0__inst_mult_12_92 ;
wire Xd_0__inst_mult_12_93 ;
wire Xd_0__inst_mult_12_94 ;
wire Xd_0__inst_mult_13_92 ;
wire Xd_0__inst_mult_13_93 ;
wire Xd_0__inst_mult_13_94 ;
wire Xd_0__inst_mult_10_92 ;
wire Xd_0__inst_mult_10_93 ;
wire Xd_0__inst_mult_10_94 ;
wire Xd_0__inst_mult_11_92 ;
wire Xd_0__inst_mult_11_93 ;
wire Xd_0__inst_mult_11_94 ;
wire Xd_0__inst_mult_8_92 ;
wire Xd_0__inst_mult_8_93 ;
wire Xd_0__inst_mult_8_94 ;
wire Xd_0__inst_mult_9_92 ;
wire Xd_0__inst_mult_9_93 ;
wire Xd_0__inst_mult_9_94 ;
wire Xd_0__inst_mult_6_92 ;
wire Xd_0__inst_mult_6_93 ;
wire Xd_0__inst_mult_6_94 ;
wire Xd_0__inst_mult_7_92 ;
wire Xd_0__inst_mult_7_93 ;
wire Xd_0__inst_mult_7_94 ;
wire Xd_0__inst_mult_4_92 ;
wire Xd_0__inst_mult_4_93 ;
wire Xd_0__inst_mult_4_94 ;
wire Xd_0__inst_mult_5_92 ;
wire Xd_0__inst_mult_5_93 ;
wire Xd_0__inst_mult_5_94 ;
wire Xd_0__inst_mult_2_92 ;
wire Xd_0__inst_mult_2_93 ;
wire Xd_0__inst_mult_2_94 ;
wire Xd_0__inst_mult_3_92 ;
wire Xd_0__inst_mult_3_93 ;
wire Xd_0__inst_mult_3_94 ;
wire Xd_0__inst_mult_0_92 ;
wire Xd_0__inst_mult_0_93 ;
wire Xd_0__inst_mult_0_94 ;
wire Xd_0__inst_mult_1_92 ;
wire Xd_0__inst_mult_1_93 ;
wire Xd_0__inst_mult_1_94 ;
wire Xd_0__inst_mult_28_97 ;
wire Xd_0__inst_mult_28_98 ;
wire Xd_0__inst_mult_29_97 ;
wire Xd_0__inst_mult_29_98 ;
wire Xd_0__inst_mult_26_97 ;
wire Xd_0__inst_mult_26_98 ;
wire Xd_0__inst_mult_27_97 ;
wire Xd_0__inst_mult_27_98 ;
wire Xd_0__inst_mult_24_97 ;
wire Xd_0__inst_mult_24_98 ;
wire Xd_0__inst_mult_25_101 ;
wire Xd_0__inst_mult_25_102 ;
wire Xd_0__inst_mult_22_101 ;
wire Xd_0__inst_mult_22_102 ;
wire Xd_0__inst_mult_23_97 ;
wire Xd_0__inst_mult_23_98 ;
wire Xd_0__inst_mult_20_97 ;
wire Xd_0__inst_mult_20_98 ;
wire Xd_0__inst_mult_21_97 ;
wire Xd_0__inst_mult_21_98 ;
wire Xd_0__inst_mult_18_97 ;
wire Xd_0__inst_mult_18_98 ;
wire Xd_0__inst_mult_19_97 ;
wire Xd_0__inst_mult_19_98 ;
wire Xd_0__inst_mult_30_100 ;
wire Xd_0__inst_mult_30_101 ;
wire Xd_0__inst_mult_30_102 ;
wire Xd_0__inst_mult_31_100 ;
wire Xd_0__inst_mult_31_101 ;
wire Xd_0__inst_mult_31_102 ;
wire Xd_0__inst_mult_16_97 ;
wire Xd_0__inst_mult_16_98 ;
wire Xd_0__inst_mult_17_97 ;
wire Xd_0__inst_mult_17_98 ;
wire Xd_0__inst_mult_14_97 ;
wire Xd_0__inst_mult_14_98 ;
wire Xd_0__inst_mult_15_97 ;
wire Xd_0__inst_mult_15_98 ;
wire Xd_0__inst_mult_12_97 ;
wire Xd_0__inst_mult_12_98 ;
wire Xd_0__inst_mult_13_97 ;
wire Xd_0__inst_mult_13_98 ;
wire Xd_0__inst_mult_10_97 ;
wire Xd_0__inst_mult_10_98 ;
wire Xd_0__inst_mult_11_97 ;
wire Xd_0__inst_mult_11_98 ;
wire Xd_0__inst_mult_8_97 ;
wire Xd_0__inst_mult_8_98 ;
wire Xd_0__inst_mult_9_97 ;
wire Xd_0__inst_mult_9_98 ;
wire Xd_0__inst_mult_6_97 ;
wire Xd_0__inst_mult_6_98 ;
wire Xd_0__inst_mult_7_97 ;
wire Xd_0__inst_mult_7_98 ;
wire Xd_0__inst_mult_4_97 ;
wire Xd_0__inst_mult_4_98 ;
wire Xd_0__inst_mult_5_97 ;
wire Xd_0__inst_mult_5_98 ;
wire Xd_0__inst_mult_2_97 ;
wire Xd_0__inst_mult_2_98 ;
wire Xd_0__inst_mult_3_97 ;
wire Xd_0__inst_mult_3_98 ;
wire Xd_0__inst_mult_0_97 ;
wire Xd_0__inst_mult_0_98 ;
wire Xd_0__inst_mult_1_97 ;
wire Xd_0__inst_mult_1_98 ;
wire Xd_0__inst_mult_30_104 ;
wire Xd_0__inst_mult_30_105 ;
wire Xd_0__inst_mult_30_106 ;
wire Xd_0__inst_mult_30_108 ;
wire Xd_0__inst_mult_30_109 ;
wire Xd_0__inst_mult_30_110 ;
wire Xd_0__inst_mult_31_104 ;
wire Xd_0__inst_mult_31_105 ;
wire Xd_0__inst_mult_31_106 ;
wire Xd_0__inst_mult_31_108 ;
wire Xd_0__inst_mult_31_109 ;
wire Xd_0__inst_mult_31_110 ;
wire Xd_0__inst_mult_30_112 ;
wire Xd_0__inst_mult_30_113 ;
wire Xd_0__inst_mult_30_114 ;
wire Xd_0__inst_mult_30_116 ;
wire Xd_0__inst_mult_30_117 ;
wire Xd_0__inst_mult_30_118 ;
wire Xd_0__inst_mult_31_112 ;
wire Xd_0__inst_mult_31_113 ;
wire Xd_0__inst_mult_31_114 ;
wire Xd_0__inst_mult_31_116 ;
wire Xd_0__inst_mult_31_117 ;
wire Xd_0__inst_mult_31_118 ;
wire Xd_0__inst_mult_30_120 ;
wire Xd_0__inst_mult_30_121 ;
wire Xd_0__inst_mult_30_122 ;
wire Xd_0__inst_mult_30_124 ;
wire Xd_0__inst_mult_30_125 ;
wire Xd_0__inst_mult_30_126 ;
wire Xd_0__inst_mult_31_120 ;
wire Xd_0__inst_mult_31_121 ;
wire Xd_0__inst_mult_31_122 ;
wire Xd_0__inst_mult_31_124 ;
wire Xd_0__inst_mult_31_125 ;
wire Xd_0__inst_mult_31_126 ;
wire Xd_0__inst_mult_30_128 ;
wire Xd_0__inst_mult_30_129 ;
wire Xd_0__inst_mult_30_130 ;
wire Xd_0__inst_mult_30_132 ;
wire Xd_0__inst_mult_30_133 ;
wire Xd_0__inst_mult_30_134 ;
wire Xd_0__inst_mult_31_128 ;
wire Xd_0__inst_mult_31_129 ;
wire Xd_0__inst_mult_31_130 ;
wire Xd_0__inst_mult_31_132 ;
wire Xd_0__inst_mult_31_133 ;
wire Xd_0__inst_mult_31_134 ;
wire Xd_0__inst_mult_30_136 ;
wire Xd_0__inst_mult_30_137 ;
wire Xd_0__inst_mult_30_138 ;
wire Xd_0__inst_mult_30_140 ;
wire Xd_0__inst_mult_30_141 ;
wire Xd_0__inst_mult_30_142 ;
wire Xd_0__inst_mult_31_136 ;
wire Xd_0__inst_mult_31_137 ;
wire Xd_0__inst_mult_31_138 ;
wire Xd_0__inst_mult_31_140 ;
wire Xd_0__inst_mult_31_141 ;
wire Xd_0__inst_mult_31_142 ;
wire Xd_0__inst_mult_30_144 ;
wire Xd_0__inst_mult_30_145 ;
wire Xd_0__inst_mult_30_146 ;
wire Xd_0__inst_mult_30_148 ;
wire Xd_0__inst_mult_30_149 ;
wire Xd_0__inst_mult_30_150 ;
wire Xd_0__inst_mult_31_144 ;
wire Xd_0__inst_mult_31_145 ;
wire Xd_0__inst_mult_31_146 ;
wire Xd_0__inst_mult_31_148 ;
wire Xd_0__inst_mult_31_149 ;
wire Xd_0__inst_mult_31_150 ;
wire Xd_0__inst_mult_30_152 ;
wire Xd_0__inst_mult_31_152 ;
wire Xd_0__inst_mult_14_100 ;
wire Xd_0__inst_mult_14_101 ;
wire Xd_0__inst_mult_14_102 ;
wire Xd_0__inst_mult_19_100 ;
wire Xd_0__inst_mult_19_101 ;
wire Xd_0__inst_mult_19_102 ;
wire Xd_0__inst_mult_21_100 ;
wire Xd_0__inst_mult_21_101 ;
wire Xd_0__inst_mult_21_102 ;
wire Xd_0__inst_mult_18_100 ;
wire Xd_0__inst_mult_18_101 ;
wire Xd_0__inst_mult_18_102 ;
wire Xd_0__inst_mult_17_100 ;
wire Xd_0__inst_mult_17_101 ;
wire Xd_0__inst_mult_17_102 ;
wire Xd_0__inst_mult_16_100 ;
wire Xd_0__inst_mult_16_101 ;
wire Xd_0__inst_mult_16_102 ;
wire Xd_0__inst_mult_20_100 ;
wire Xd_0__inst_mult_20_101 ;
wire Xd_0__inst_mult_20_102 ;
wire Xd_0__inst_mult_28_100 ;
wire Xd_0__inst_mult_28_101 ;
wire Xd_0__inst_mult_28_102 ;
wire Xd_0__inst_mult_12_100 ;
wire Xd_0__inst_mult_12_101 ;
wire Xd_0__inst_mult_12_102 ;
wire Xd_0__inst_mult_5_100 ;
wire Xd_0__inst_mult_5_101 ;
wire Xd_0__inst_mult_5_102 ;
wire Xd_0__inst_mult_15_100 ;
wire Xd_0__inst_mult_15_101 ;
wire Xd_0__inst_mult_15_102 ;
wire Xd_0__inst_mult_7_100 ;
wire Xd_0__inst_mult_7_101 ;
wire Xd_0__inst_mult_7_102 ;
wire Xd_0__inst_mult_25_104 ;
wire Xd_0__inst_mult_25_105 ;
wire Xd_0__inst_mult_25_106 ;
wire Xd_0__inst_mult_22_104 ;
wire Xd_0__inst_mult_22_105 ;
wire Xd_0__inst_mult_22_106 ;
wire Xd_0__inst_mult_6_100 ;
wire Xd_0__inst_mult_6_101 ;
wire Xd_0__inst_mult_6_102 ;
wire Xd_0__inst_mult_9_100 ;
wire Xd_0__inst_mult_9_101 ;
wire Xd_0__inst_mult_9_102 ;
wire Xd_0__inst_mult_8_100 ;
wire Xd_0__inst_mult_8_101 ;
wire Xd_0__inst_mult_8_102 ;
wire Xd_0__inst_mult_11_100 ;
wire Xd_0__inst_mult_11_101 ;
wire Xd_0__inst_mult_11_102 ;
wire Xd_0__inst_mult_10_100 ;
wire Xd_0__inst_mult_10_101 ;
wire Xd_0__inst_mult_10_102 ;
wire Xd_0__inst_mult_13_100 ;
wire Xd_0__inst_mult_13_101 ;
wire Xd_0__inst_mult_13_102 ;
wire Xd_0__inst_mult_4_100 ;
wire Xd_0__inst_mult_4_101 ;
wire Xd_0__inst_mult_4_102 ;
wire Xd_0__inst_mult_2_100 ;
wire Xd_0__inst_mult_2_101 ;
wire Xd_0__inst_mult_2_102 ;
wire Xd_0__inst_mult_3_100 ;
wire Xd_0__inst_mult_3_101 ;
wire Xd_0__inst_mult_3_102 ;
wire Xd_0__inst_mult_0_100 ;
wire Xd_0__inst_mult_0_101 ;
wire Xd_0__inst_mult_0_102 ;
wire Xd_0__inst_mult_1_100 ;
wire Xd_0__inst_mult_1_101 ;
wire Xd_0__inst_mult_1_102 ;
wire Xd_0__inst_mult_23_100 ;
wire Xd_0__inst_mult_23_101 ;
wire Xd_0__inst_mult_23_102 ;
wire Xd_0__inst_mult_29_100 ;
wire Xd_0__inst_mult_29_101 ;
wire Xd_0__inst_mult_29_102 ;
wire Xd_0__inst_mult_26_100 ;
wire Xd_0__inst_mult_26_101 ;
wire Xd_0__inst_mult_26_102 ;
wire Xd_0__inst_mult_24_100 ;
wire Xd_0__inst_mult_24_101 ;
wire Xd_0__inst_mult_24_102 ;
wire Xd_0__inst_mult_27_100 ;
wire Xd_0__inst_mult_27_101 ;
wire Xd_0__inst_mult_27_102 ;
wire Xd_0__inst_mult_28_104 ;
wire Xd_0__inst_mult_28_105 ;
wire Xd_0__inst_mult_28_106 ;
wire Xd_0__inst_mult_29_104 ;
wire Xd_0__inst_mult_29_105 ;
wire Xd_0__inst_mult_29_106 ;
wire Xd_0__inst_mult_26_104 ;
wire Xd_0__inst_mult_26_105 ;
wire Xd_0__inst_mult_26_106 ;
wire Xd_0__inst_mult_27_104 ;
wire Xd_0__inst_mult_27_105 ;
wire Xd_0__inst_mult_27_106 ;
wire Xd_0__inst_mult_24_104 ;
wire Xd_0__inst_mult_24_105 ;
wire Xd_0__inst_mult_24_106 ;
wire Xd_0__inst_mult_25_108 ;
wire Xd_0__inst_mult_25_109 ;
wire Xd_0__inst_mult_25_110 ;
wire Xd_0__inst_mult_22_108 ;
wire Xd_0__inst_mult_22_109 ;
wire Xd_0__inst_mult_22_110 ;
wire Xd_0__inst_mult_23_104 ;
wire Xd_0__inst_mult_23_105 ;
wire Xd_0__inst_mult_23_106 ;
wire Xd_0__inst_mult_20_104 ;
wire Xd_0__inst_mult_20_105 ;
wire Xd_0__inst_mult_20_106 ;
wire Xd_0__inst_mult_21_104 ;
wire Xd_0__inst_mult_21_105 ;
wire Xd_0__inst_mult_21_106 ;
wire Xd_0__inst_mult_18_104 ;
wire Xd_0__inst_mult_18_105 ;
wire Xd_0__inst_mult_18_106 ;
wire Xd_0__inst_mult_19_104 ;
wire Xd_0__inst_mult_19_105 ;
wire Xd_0__inst_mult_19_106 ;
wire Xd_0__inst_mult_16_104 ;
wire Xd_0__inst_mult_16_105 ;
wire Xd_0__inst_mult_16_106 ;
wire Xd_0__inst_mult_17_104 ;
wire Xd_0__inst_mult_17_105 ;
wire Xd_0__inst_mult_17_106 ;
wire Xd_0__inst_mult_14_104 ;
wire Xd_0__inst_mult_14_105 ;
wire Xd_0__inst_mult_14_106 ;
wire Xd_0__inst_mult_15_104 ;
wire Xd_0__inst_mult_15_105 ;
wire Xd_0__inst_mult_15_106 ;
wire Xd_0__inst_mult_12_104 ;
wire Xd_0__inst_mult_12_105 ;
wire Xd_0__inst_mult_12_106 ;
wire Xd_0__inst_mult_13_104 ;
wire Xd_0__inst_mult_13_105 ;
wire Xd_0__inst_mult_13_106 ;
wire Xd_0__inst_mult_10_104 ;
wire Xd_0__inst_mult_10_105 ;
wire Xd_0__inst_mult_10_106 ;
wire Xd_0__inst_mult_11_104 ;
wire Xd_0__inst_mult_11_105 ;
wire Xd_0__inst_mult_11_106 ;
wire Xd_0__inst_mult_8_104 ;
wire Xd_0__inst_mult_8_105 ;
wire Xd_0__inst_mult_8_106 ;
wire Xd_0__inst_mult_9_104 ;
wire Xd_0__inst_mult_9_105 ;
wire Xd_0__inst_mult_9_106 ;
wire Xd_0__inst_mult_6_104 ;
wire Xd_0__inst_mult_6_105 ;
wire Xd_0__inst_mult_6_106 ;
wire Xd_0__inst_mult_7_104 ;
wire Xd_0__inst_mult_7_105 ;
wire Xd_0__inst_mult_7_106 ;
wire Xd_0__inst_mult_4_104 ;
wire Xd_0__inst_mult_4_105 ;
wire Xd_0__inst_mult_4_106 ;
wire Xd_0__inst_mult_5_104 ;
wire Xd_0__inst_mult_5_105 ;
wire Xd_0__inst_mult_5_106 ;
wire Xd_0__inst_mult_2_104 ;
wire Xd_0__inst_mult_2_105 ;
wire Xd_0__inst_mult_2_106 ;
wire Xd_0__inst_mult_3_104 ;
wire Xd_0__inst_mult_3_105 ;
wire Xd_0__inst_mult_3_106 ;
wire Xd_0__inst_mult_0_104 ;
wire Xd_0__inst_mult_0_105 ;
wire Xd_0__inst_mult_0_106 ;
wire Xd_0__inst_mult_1_104 ;
wire Xd_0__inst_mult_1_105 ;
wire Xd_0__inst_mult_1_106 ;
wire Xd_0__inst_mult_28_108 ;
wire Xd_0__inst_mult_28_109 ;
wire Xd_0__inst_mult_28_110 ;
wire Xd_0__inst_mult_28_112 ;
wire Xd_0__inst_mult_28_113 ;
wire Xd_0__inst_mult_28_114 ;
wire Xd_0__inst_mult_29_108 ;
wire Xd_0__inst_mult_29_109 ;
wire Xd_0__inst_mult_29_110 ;
wire Xd_0__inst_mult_29_112 ;
wire Xd_0__inst_mult_29_113 ;
wire Xd_0__inst_mult_29_114 ;
wire Xd_0__inst_mult_26_108 ;
wire Xd_0__inst_mult_26_109 ;
wire Xd_0__inst_mult_26_110 ;
wire Xd_0__inst_mult_26_112 ;
wire Xd_0__inst_mult_26_113 ;
wire Xd_0__inst_mult_26_114 ;
wire Xd_0__inst_mult_27_108 ;
wire Xd_0__inst_mult_27_109 ;
wire Xd_0__inst_mult_27_110 ;
wire Xd_0__inst_mult_27_112 ;
wire Xd_0__inst_mult_27_113 ;
wire Xd_0__inst_mult_27_114 ;
wire Xd_0__inst_mult_24_108 ;
wire Xd_0__inst_mult_24_109 ;
wire Xd_0__inst_mult_24_110 ;
wire Xd_0__inst_mult_24_112 ;
wire Xd_0__inst_mult_24_113 ;
wire Xd_0__inst_mult_24_114 ;
wire Xd_0__inst_mult_25_112 ;
wire Xd_0__inst_mult_25_113 ;
wire Xd_0__inst_mult_25_114 ;
wire Xd_0__inst_mult_25_116 ;
wire Xd_0__inst_mult_25_117 ;
wire Xd_0__inst_mult_25_118 ;
wire Xd_0__inst_mult_22_112 ;
wire Xd_0__inst_mult_22_113 ;
wire Xd_0__inst_mult_22_114 ;
wire Xd_0__inst_mult_22_116 ;
wire Xd_0__inst_mult_22_117 ;
wire Xd_0__inst_mult_22_118 ;
wire Xd_0__inst_mult_23_108 ;
wire Xd_0__inst_mult_23_109 ;
wire Xd_0__inst_mult_23_110 ;
wire Xd_0__inst_mult_23_112 ;
wire Xd_0__inst_mult_23_113 ;
wire Xd_0__inst_mult_23_114 ;
wire Xd_0__inst_mult_20_108 ;
wire Xd_0__inst_mult_20_109 ;
wire Xd_0__inst_mult_20_110 ;
wire Xd_0__inst_mult_20_112 ;
wire Xd_0__inst_mult_20_113 ;
wire Xd_0__inst_mult_20_114 ;
wire Xd_0__inst_mult_21_108 ;
wire Xd_0__inst_mult_21_109 ;
wire Xd_0__inst_mult_21_110 ;
wire Xd_0__inst_mult_21_112 ;
wire Xd_0__inst_mult_21_113 ;
wire Xd_0__inst_mult_21_114 ;
wire Xd_0__inst_mult_18_108 ;
wire Xd_0__inst_mult_18_109 ;
wire Xd_0__inst_mult_18_110 ;
wire Xd_0__inst_mult_18_112 ;
wire Xd_0__inst_mult_18_113 ;
wire Xd_0__inst_mult_18_114 ;
wire Xd_0__inst_mult_19_108 ;
wire Xd_0__inst_mult_19_109 ;
wire Xd_0__inst_mult_19_110 ;
wire Xd_0__inst_mult_19_112 ;
wire Xd_0__inst_mult_19_113 ;
wire Xd_0__inst_mult_19_114 ;
wire Xd_0__inst_mult_30_157 ;
wire Xd_0__inst_mult_30_158 ;
wire Xd_0__inst_mult_31_157 ;
wire Xd_0__inst_mult_31_158 ;
wire Xd_0__inst_mult_16_108 ;
wire Xd_0__inst_mult_16_109 ;
wire Xd_0__inst_mult_16_110 ;
wire Xd_0__inst_mult_16_112 ;
wire Xd_0__inst_mult_16_113 ;
wire Xd_0__inst_mult_16_114 ;
wire Xd_0__inst_mult_17_108 ;
wire Xd_0__inst_mult_17_109 ;
wire Xd_0__inst_mult_17_110 ;
wire Xd_0__inst_mult_17_112 ;
wire Xd_0__inst_mult_17_113 ;
wire Xd_0__inst_mult_17_114 ;
wire Xd_0__inst_mult_14_108 ;
wire Xd_0__inst_mult_14_109 ;
wire Xd_0__inst_mult_14_110 ;
wire Xd_0__inst_mult_14_112 ;
wire Xd_0__inst_mult_14_113 ;
wire Xd_0__inst_mult_14_114 ;
wire Xd_0__inst_mult_15_108 ;
wire Xd_0__inst_mult_15_109 ;
wire Xd_0__inst_mult_15_110 ;
wire Xd_0__inst_mult_15_112 ;
wire Xd_0__inst_mult_15_113 ;
wire Xd_0__inst_mult_15_114 ;
wire Xd_0__inst_mult_12_108 ;
wire Xd_0__inst_mult_12_109 ;
wire Xd_0__inst_mult_12_110 ;
wire Xd_0__inst_mult_12_112 ;
wire Xd_0__inst_mult_12_113 ;
wire Xd_0__inst_mult_12_114 ;
wire Xd_0__inst_mult_13_108 ;
wire Xd_0__inst_mult_13_109 ;
wire Xd_0__inst_mult_13_110 ;
wire Xd_0__inst_mult_13_112 ;
wire Xd_0__inst_mult_13_113 ;
wire Xd_0__inst_mult_13_114 ;
wire Xd_0__inst_mult_10_108 ;
wire Xd_0__inst_mult_10_109 ;
wire Xd_0__inst_mult_10_110 ;
wire Xd_0__inst_mult_10_112 ;
wire Xd_0__inst_mult_10_113 ;
wire Xd_0__inst_mult_10_114 ;
wire Xd_0__inst_mult_11_108 ;
wire Xd_0__inst_mult_11_109 ;
wire Xd_0__inst_mult_11_110 ;
wire Xd_0__inst_mult_11_112 ;
wire Xd_0__inst_mult_11_113 ;
wire Xd_0__inst_mult_11_114 ;
wire Xd_0__inst_mult_8_108 ;
wire Xd_0__inst_mult_8_109 ;
wire Xd_0__inst_mult_8_110 ;
wire Xd_0__inst_mult_8_112 ;
wire Xd_0__inst_mult_8_113 ;
wire Xd_0__inst_mult_8_114 ;
wire Xd_0__inst_mult_9_108 ;
wire Xd_0__inst_mult_9_109 ;
wire Xd_0__inst_mult_9_110 ;
wire Xd_0__inst_mult_9_112 ;
wire Xd_0__inst_mult_9_113 ;
wire Xd_0__inst_mult_9_114 ;
wire Xd_0__inst_mult_6_108 ;
wire Xd_0__inst_mult_6_109 ;
wire Xd_0__inst_mult_6_110 ;
wire Xd_0__inst_mult_6_112 ;
wire Xd_0__inst_mult_6_113 ;
wire Xd_0__inst_mult_6_114 ;
wire Xd_0__inst_mult_7_108 ;
wire Xd_0__inst_mult_7_109 ;
wire Xd_0__inst_mult_7_110 ;
wire Xd_0__inst_mult_7_112 ;
wire Xd_0__inst_mult_7_113 ;
wire Xd_0__inst_mult_7_114 ;
wire Xd_0__inst_mult_4_108 ;
wire Xd_0__inst_mult_4_109 ;
wire Xd_0__inst_mult_4_110 ;
wire Xd_0__inst_mult_4_112 ;
wire Xd_0__inst_mult_4_113 ;
wire Xd_0__inst_mult_4_114 ;
wire Xd_0__inst_mult_5_108 ;
wire Xd_0__inst_mult_5_109 ;
wire Xd_0__inst_mult_5_110 ;
wire Xd_0__inst_mult_5_112 ;
wire Xd_0__inst_mult_5_113 ;
wire Xd_0__inst_mult_5_114 ;
wire Xd_0__inst_mult_2_108 ;
wire Xd_0__inst_mult_2_109 ;
wire Xd_0__inst_mult_2_110 ;
wire Xd_0__inst_mult_2_112 ;
wire Xd_0__inst_mult_2_113 ;
wire Xd_0__inst_mult_2_114 ;
wire Xd_0__inst_mult_3_108 ;
wire Xd_0__inst_mult_3_109 ;
wire Xd_0__inst_mult_3_110 ;
wire Xd_0__inst_mult_3_112 ;
wire Xd_0__inst_mult_3_113 ;
wire Xd_0__inst_mult_3_114 ;
wire Xd_0__inst_mult_0_108 ;
wire Xd_0__inst_mult_0_109 ;
wire Xd_0__inst_mult_0_110 ;
wire Xd_0__inst_mult_0_112 ;
wire Xd_0__inst_mult_0_113 ;
wire Xd_0__inst_mult_0_114 ;
wire Xd_0__inst_mult_1_108 ;
wire Xd_0__inst_mult_1_109 ;
wire Xd_0__inst_mult_1_110 ;
wire Xd_0__inst_mult_1_112 ;
wire Xd_0__inst_mult_1_113 ;
wire Xd_0__inst_mult_1_114 ;
wire Xd_0__inst_mult_28_116 ;
wire Xd_0__inst_mult_28_117 ;
wire Xd_0__inst_mult_28_118 ;
wire Xd_0__inst_mult_28_120 ;
wire Xd_0__inst_mult_28_121 ;
wire Xd_0__inst_mult_28_122 ;
wire Xd_0__inst_mult_29_116 ;
wire Xd_0__inst_mult_29_117 ;
wire Xd_0__inst_mult_29_118 ;
wire Xd_0__inst_mult_29_120 ;
wire Xd_0__inst_mult_29_121 ;
wire Xd_0__inst_mult_29_122 ;
wire Xd_0__inst_mult_26_116 ;
wire Xd_0__inst_mult_26_117 ;
wire Xd_0__inst_mult_26_118 ;
wire Xd_0__inst_mult_26_120 ;
wire Xd_0__inst_mult_26_121 ;
wire Xd_0__inst_mult_26_122 ;
wire Xd_0__inst_mult_27_116 ;
wire Xd_0__inst_mult_27_117 ;
wire Xd_0__inst_mult_27_118 ;
wire Xd_0__inst_mult_27_120 ;
wire Xd_0__inst_mult_27_121 ;
wire Xd_0__inst_mult_27_122 ;
wire Xd_0__inst_mult_24_116 ;
wire Xd_0__inst_mult_24_117 ;
wire Xd_0__inst_mult_24_118 ;
wire Xd_0__inst_mult_24_120 ;
wire Xd_0__inst_mult_24_121 ;
wire Xd_0__inst_mult_24_122 ;
wire Xd_0__inst_mult_25_120 ;
wire Xd_0__inst_mult_25_121 ;
wire Xd_0__inst_mult_25_122 ;
wire Xd_0__inst_mult_25_124 ;
wire Xd_0__inst_mult_25_125 ;
wire Xd_0__inst_mult_25_126 ;
wire Xd_0__inst_mult_22_120 ;
wire Xd_0__inst_mult_22_121 ;
wire Xd_0__inst_mult_22_122 ;
wire Xd_0__inst_mult_22_124 ;
wire Xd_0__inst_mult_22_125 ;
wire Xd_0__inst_mult_22_126 ;
wire Xd_0__inst_mult_23_116 ;
wire Xd_0__inst_mult_23_117 ;
wire Xd_0__inst_mult_23_118 ;
wire Xd_0__inst_mult_23_120 ;
wire Xd_0__inst_mult_23_121 ;
wire Xd_0__inst_mult_23_122 ;
wire Xd_0__inst_mult_20_116 ;
wire Xd_0__inst_mult_20_117 ;
wire Xd_0__inst_mult_20_118 ;
wire Xd_0__inst_mult_20_120 ;
wire Xd_0__inst_mult_20_121 ;
wire Xd_0__inst_mult_20_122 ;
wire Xd_0__inst_mult_21_116 ;
wire Xd_0__inst_mult_21_117 ;
wire Xd_0__inst_mult_21_118 ;
wire Xd_0__inst_mult_21_120 ;
wire Xd_0__inst_mult_21_121 ;
wire Xd_0__inst_mult_21_122 ;
wire Xd_0__inst_mult_18_116 ;
wire Xd_0__inst_mult_18_117 ;
wire Xd_0__inst_mult_18_118 ;
wire Xd_0__inst_mult_18_120 ;
wire Xd_0__inst_mult_18_121 ;
wire Xd_0__inst_mult_18_122 ;
wire Xd_0__inst_mult_19_116 ;
wire Xd_0__inst_mult_19_117 ;
wire Xd_0__inst_mult_19_118 ;
wire Xd_0__inst_mult_19_120 ;
wire Xd_0__inst_mult_19_121 ;
wire Xd_0__inst_mult_19_122 ;
wire Xd_0__inst_mult_16_116 ;
wire Xd_0__inst_mult_16_117 ;
wire Xd_0__inst_mult_16_118 ;
wire Xd_0__inst_mult_16_120 ;
wire Xd_0__inst_mult_16_121 ;
wire Xd_0__inst_mult_16_122 ;
wire Xd_0__inst_mult_17_116 ;
wire Xd_0__inst_mult_17_117 ;
wire Xd_0__inst_mult_17_118 ;
wire Xd_0__inst_mult_17_120 ;
wire Xd_0__inst_mult_17_121 ;
wire Xd_0__inst_mult_17_122 ;
wire Xd_0__inst_mult_14_116 ;
wire Xd_0__inst_mult_14_117 ;
wire Xd_0__inst_mult_14_118 ;
wire Xd_0__inst_mult_14_120 ;
wire Xd_0__inst_mult_14_121 ;
wire Xd_0__inst_mult_14_122 ;
wire Xd_0__inst_mult_15_116 ;
wire Xd_0__inst_mult_15_117 ;
wire Xd_0__inst_mult_15_118 ;
wire Xd_0__inst_mult_15_120 ;
wire Xd_0__inst_mult_15_121 ;
wire Xd_0__inst_mult_15_122 ;
wire Xd_0__inst_mult_12_116 ;
wire Xd_0__inst_mult_12_117 ;
wire Xd_0__inst_mult_12_118 ;
wire Xd_0__inst_mult_12_120 ;
wire Xd_0__inst_mult_12_121 ;
wire Xd_0__inst_mult_12_122 ;
wire Xd_0__inst_mult_13_116 ;
wire Xd_0__inst_mult_13_117 ;
wire Xd_0__inst_mult_13_118 ;
wire Xd_0__inst_mult_13_120 ;
wire Xd_0__inst_mult_13_121 ;
wire Xd_0__inst_mult_13_122 ;
wire Xd_0__inst_mult_10_116 ;
wire Xd_0__inst_mult_10_117 ;
wire Xd_0__inst_mult_10_118 ;
wire Xd_0__inst_mult_10_120 ;
wire Xd_0__inst_mult_10_121 ;
wire Xd_0__inst_mult_10_122 ;
wire Xd_0__inst_mult_11_116 ;
wire Xd_0__inst_mult_11_117 ;
wire Xd_0__inst_mult_11_118 ;
wire Xd_0__inst_mult_11_120 ;
wire Xd_0__inst_mult_11_121 ;
wire Xd_0__inst_mult_11_122 ;
wire Xd_0__inst_mult_8_116 ;
wire Xd_0__inst_mult_8_117 ;
wire Xd_0__inst_mult_8_118 ;
wire Xd_0__inst_mult_8_120 ;
wire Xd_0__inst_mult_8_121 ;
wire Xd_0__inst_mult_8_122 ;
wire Xd_0__inst_mult_9_116 ;
wire Xd_0__inst_mult_9_117 ;
wire Xd_0__inst_mult_9_118 ;
wire Xd_0__inst_mult_9_120 ;
wire Xd_0__inst_mult_9_121 ;
wire Xd_0__inst_mult_9_122 ;
wire Xd_0__inst_mult_6_116 ;
wire Xd_0__inst_mult_6_117 ;
wire Xd_0__inst_mult_6_118 ;
wire Xd_0__inst_mult_6_120 ;
wire Xd_0__inst_mult_6_121 ;
wire Xd_0__inst_mult_6_122 ;
wire Xd_0__inst_mult_7_116 ;
wire Xd_0__inst_mult_7_117 ;
wire Xd_0__inst_mult_7_118 ;
wire Xd_0__inst_mult_7_120 ;
wire Xd_0__inst_mult_7_121 ;
wire Xd_0__inst_mult_7_122 ;
wire Xd_0__inst_mult_4_116 ;
wire Xd_0__inst_mult_4_117 ;
wire Xd_0__inst_mult_4_118 ;
wire Xd_0__inst_mult_4_120 ;
wire Xd_0__inst_mult_4_121 ;
wire Xd_0__inst_mult_4_122 ;
wire Xd_0__inst_mult_5_116 ;
wire Xd_0__inst_mult_5_117 ;
wire Xd_0__inst_mult_5_118 ;
wire Xd_0__inst_mult_5_120 ;
wire Xd_0__inst_mult_5_121 ;
wire Xd_0__inst_mult_5_122 ;
wire Xd_0__inst_mult_2_116 ;
wire Xd_0__inst_mult_2_117 ;
wire Xd_0__inst_mult_2_118 ;
wire Xd_0__inst_mult_2_120 ;
wire Xd_0__inst_mult_2_121 ;
wire Xd_0__inst_mult_2_122 ;
wire Xd_0__inst_mult_3_116 ;
wire Xd_0__inst_mult_3_117 ;
wire Xd_0__inst_mult_3_118 ;
wire Xd_0__inst_mult_3_120 ;
wire Xd_0__inst_mult_3_121 ;
wire Xd_0__inst_mult_3_122 ;
wire Xd_0__inst_mult_0_116 ;
wire Xd_0__inst_mult_0_117 ;
wire Xd_0__inst_mult_0_118 ;
wire Xd_0__inst_mult_0_120 ;
wire Xd_0__inst_mult_0_121 ;
wire Xd_0__inst_mult_0_122 ;
wire Xd_0__inst_mult_1_116 ;
wire Xd_0__inst_mult_1_117 ;
wire Xd_0__inst_mult_1_118 ;
wire Xd_0__inst_mult_1_120 ;
wire Xd_0__inst_mult_1_121 ;
wire Xd_0__inst_mult_1_122 ;
wire Xd_0__inst_mult_28_124 ;
wire Xd_0__inst_mult_28_125 ;
wire Xd_0__inst_mult_28_126 ;
wire Xd_0__inst_mult_28_128 ;
wire Xd_0__inst_mult_28_129 ;
wire Xd_0__inst_mult_28_130 ;
wire Xd_0__inst_mult_29_124 ;
wire Xd_0__inst_mult_29_125 ;
wire Xd_0__inst_mult_29_126 ;
wire Xd_0__inst_mult_29_128 ;
wire Xd_0__inst_mult_29_129 ;
wire Xd_0__inst_mult_29_130 ;
wire Xd_0__inst_mult_26_124 ;
wire Xd_0__inst_mult_26_125 ;
wire Xd_0__inst_mult_26_126 ;
wire Xd_0__inst_mult_26_128 ;
wire Xd_0__inst_mult_26_129 ;
wire Xd_0__inst_mult_26_130 ;
wire Xd_0__inst_mult_27_124 ;
wire Xd_0__inst_mult_27_125 ;
wire Xd_0__inst_mult_27_126 ;
wire Xd_0__inst_mult_27_128 ;
wire Xd_0__inst_mult_27_129 ;
wire Xd_0__inst_mult_27_130 ;
wire Xd_0__inst_mult_24_124 ;
wire Xd_0__inst_mult_24_125 ;
wire Xd_0__inst_mult_24_126 ;
wire Xd_0__inst_mult_24_128 ;
wire Xd_0__inst_mult_24_129 ;
wire Xd_0__inst_mult_24_130 ;
wire Xd_0__inst_mult_25_128 ;
wire Xd_0__inst_mult_25_129 ;
wire Xd_0__inst_mult_25_130 ;
wire Xd_0__inst_mult_25_132 ;
wire Xd_0__inst_mult_25_133 ;
wire Xd_0__inst_mult_25_134 ;
wire Xd_0__inst_mult_22_128 ;
wire Xd_0__inst_mult_22_129 ;
wire Xd_0__inst_mult_22_130 ;
wire Xd_0__inst_mult_22_132 ;
wire Xd_0__inst_mult_22_133 ;
wire Xd_0__inst_mult_22_134 ;
wire Xd_0__inst_mult_23_124 ;
wire Xd_0__inst_mult_23_125 ;
wire Xd_0__inst_mult_23_126 ;
wire Xd_0__inst_mult_23_128 ;
wire Xd_0__inst_mult_23_129 ;
wire Xd_0__inst_mult_23_130 ;
wire Xd_0__inst_mult_20_124 ;
wire Xd_0__inst_mult_20_125 ;
wire Xd_0__inst_mult_20_126 ;
wire Xd_0__inst_mult_20_128 ;
wire Xd_0__inst_mult_20_129 ;
wire Xd_0__inst_mult_20_130 ;
wire Xd_0__inst_mult_21_124 ;
wire Xd_0__inst_mult_21_125 ;
wire Xd_0__inst_mult_21_126 ;
wire Xd_0__inst_mult_21_128 ;
wire Xd_0__inst_mult_21_129 ;
wire Xd_0__inst_mult_21_130 ;
wire Xd_0__inst_mult_18_124 ;
wire Xd_0__inst_mult_18_125 ;
wire Xd_0__inst_mult_18_126 ;
wire Xd_0__inst_mult_18_128 ;
wire Xd_0__inst_mult_18_129 ;
wire Xd_0__inst_mult_18_130 ;
wire Xd_0__inst_mult_19_124 ;
wire Xd_0__inst_mult_19_125 ;
wire Xd_0__inst_mult_19_126 ;
wire Xd_0__inst_mult_19_128 ;
wire Xd_0__inst_mult_19_129 ;
wire Xd_0__inst_mult_19_130 ;
wire Xd_0__inst_mult_16_124 ;
wire Xd_0__inst_mult_16_125 ;
wire Xd_0__inst_mult_16_126 ;
wire Xd_0__inst_mult_16_128 ;
wire Xd_0__inst_mult_16_129 ;
wire Xd_0__inst_mult_16_130 ;
wire Xd_0__inst_mult_17_124 ;
wire Xd_0__inst_mult_17_125 ;
wire Xd_0__inst_mult_17_126 ;
wire Xd_0__inst_mult_17_128 ;
wire Xd_0__inst_mult_17_129 ;
wire Xd_0__inst_mult_17_130 ;
wire Xd_0__inst_mult_14_124 ;
wire Xd_0__inst_mult_14_125 ;
wire Xd_0__inst_mult_14_126 ;
wire Xd_0__inst_mult_14_128 ;
wire Xd_0__inst_mult_14_129 ;
wire Xd_0__inst_mult_14_130 ;
wire Xd_0__inst_mult_15_124 ;
wire Xd_0__inst_mult_15_125 ;
wire Xd_0__inst_mult_15_126 ;
wire Xd_0__inst_mult_15_128 ;
wire Xd_0__inst_mult_15_129 ;
wire Xd_0__inst_mult_15_130 ;
wire Xd_0__inst_mult_12_124 ;
wire Xd_0__inst_mult_12_125 ;
wire Xd_0__inst_mult_12_126 ;
wire Xd_0__inst_mult_12_128 ;
wire Xd_0__inst_mult_12_129 ;
wire Xd_0__inst_mult_12_130 ;
wire Xd_0__inst_mult_13_124 ;
wire Xd_0__inst_mult_13_125 ;
wire Xd_0__inst_mult_13_126 ;
wire Xd_0__inst_mult_13_128 ;
wire Xd_0__inst_mult_13_129 ;
wire Xd_0__inst_mult_13_130 ;
wire Xd_0__inst_mult_10_124 ;
wire Xd_0__inst_mult_10_125 ;
wire Xd_0__inst_mult_10_126 ;
wire Xd_0__inst_mult_10_128 ;
wire Xd_0__inst_mult_10_129 ;
wire Xd_0__inst_mult_10_130 ;
wire Xd_0__inst_mult_11_124 ;
wire Xd_0__inst_mult_11_125 ;
wire Xd_0__inst_mult_11_126 ;
wire Xd_0__inst_mult_11_128 ;
wire Xd_0__inst_mult_11_129 ;
wire Xd_0__inst_mult_11_130 ;
wire Xd_0__inst_mult_8_124 ;
wire Xd_0__inst_mult_8_125 ;
wire Xd_0__inst_mult_8_126 ;
wire Xd_0__inst_mult_8_128 ;
wire Xd_0__inst_mult_8_129 ;
wire Xd_0__inst_mult_8_130 ;
wire Xd_0__inst_mult_9_124 ;
wire Xd_0__inst_mult_9_125 ;
wire Xd_0__inst_mult_9_126 ;
wire Xd_0__inst_mult_9_128 ;
wire Xd_0__inst_mult_9_129 ;
wire Xd_0__inst_mult_9_130 ;
wire Xd_0__inst_mult_6_124 ;
wire Xd_0__inst_mult_6_125 ;
wire Xd_0__inst_mult_6_126 ;
wire Xd_0__inst_mult_6_128 ;
wire Xd_0__inst_mult_6_129 ;
wire Xd_0__inst_mult_6_130 ;
wire Xd_0__inst_mult_7_124 ;
wire Xd_0__inst_mult_7_125 ;
wire Xd_0__inst_mult_7_126 ;
wire Xd_0__inst_mult_7_128 ;
wire Xd_0__inst_mult_7_129 ;
wire Xd_0__inst_mult_7_130 ;
wire Xd_0__inst_mult_4_124 ;
wire Xd_0__inst_mult_4_125 ;
wire Xd_0__inst_mult_4_126 ;
wire Xd_0__inst_mult_4_128 ;
wire Xd_0__inst_mult_4_129 ;
wire Xd_0__inst_mult_4_130 ;
wire Xd_0__inst_mult_5_124 ;
wire Xd_0__inst_mult_5_125 ;
wire Xd_0__inst_mult_5_126 ;
wire Xd_0__inst_mult_5_128 ;
wire Xd_0__inst_mult_5_129 ;
wire Xd_0__inst_mult_5_130 ;
wire Xd_0__inst_mult_2_124 ;
wire Xd_0__inst_mult_2_125 ;
wire Xd_0__inst_mult_2_126 ;
wire Xd_0__inst_mult_2_128 ;
wire Xd_0__inst_mult_2_129 ;
wire Xd_0__inst_mult_2_130 ;
wire Xd_0__inst_mult_3_124 ;
wire Xd_0__inst_mult_3_125 ;
wire Xd_0__inst_mult_3_126 ;
wire Xd_0__inst_mult_3_128 ;
wire Xd_0__inst_mult_3_129 ;
wire Xd_0__inst_mult_3_130 ;
wire Xd_0__inst_mult_0_124 ;
wire Xd_0__inst_mult_0_125 ;
wire Xd_0__inst_mult_0_126 ;
wire Xd_0__inst_mult_0_128 ;
wire Xd_0__inst_mult_0_129 ;
wire Xd_0__inst_mult_0_130 ;
wire Xd_0__inst_mult_1_124 ;
wire Xd_0__inst_mult_1_125 ;
wire Xd_0__inst_mult_1_126 ;
wire Xd_0__inst_mult_1_128 ;
wire Xd_0__inst_mult_1_129 ;
wire Xd_0__inst_mult_1_130 ;
wire Xd_0__inst_mult_28_132 ;
wire Xd_0__inst_mult_28_133 ;
wire Xd_0__inst_mult_28_134 ;
wire Xd_0__inst_mult_28_136 ;
wire Xd_0__inst_mult_28_137 ;
wire Xd_0__inst_mult_28_138 ;
wire Xd_0__inst_mult_29_132 ;
wire Xd_0__inst_mult_29_133 ;
wire Xd_0__inst_mult_29_134 ;
wire Xd_0__inst_mult_29_136 ;
wire Xd_0__inst_mult_29_137 ;
wire Xd_0__inst_mult_29_138 ;
wire Xd_0__inst_mult_26_132 ;
wire Xd_0__inst_mult_26_133 ;
wire Xd_0__inst_mult_26_134 ;
wire Xd_0__inst_mult_26_136 ;
wire Xd_0__inst_mult_26_137 ;
wire Xd_0__inst_mult_26_138 ;
wire Xd_0__inst_mult_27_132 ;
wire Xd_0__inst_mult_27_133 ;
wire Xd_0__inst_mult_27_134 ;
wire Xd_0__inst_mult_27_136 ;
wire Xd_0__inst_mult_27_137 ;
wire Xd_0__inst_mult_27_138 ;
wire Xd_0__inst_mult_24_132 ;
wire Xd_0__inst_mult_24_133 ;
wire Xd_0__inst_mult_24_134 ;
wire Xd_0__inst_mult_24_136 ;
wire Xd_0__inst_mult_24_137 ;
wire Xd_0__inst_mult_24_138 ;
wire Xd_0__inst_mult_25_136 ;
wire Xd_0__inst_mult_25_137 ;
wire Xd_0__inst_mult_25_138 ;
wire Xd_0__inst_mult_25_140 ;
wire Xd_0__inst_mult_25_141 ;
wire Xd_0__inst_mult_25_142 ;
wire Xd_0__inst_mult_22_136 ;
wire Xd_0__inst_mult_22_137 ;
wire Xd_0__inst_mult_22_138 ;
wire Xd_0__inst_mult_22_140 ;
wire Xd_0__inst_mult_22_141 ;
wire Xd_0__inst_mult_22_142 ;
wire Xd_0__inst_mult_23_132 ;
wire Xd_0__inst_mult_23_133 ;
wire Xd_0__inst_mult_23_134 ;
wire Xd_0__inst_mult_23_136 ;
wire Xd_0__inst_mult_23_137 ;
wire Xd_0__inst_mult_23_138 ;
wire Xd_0__inst_mult_20_132 ;
wire Xd_0__inst_mult_20_133 ;
wire Xd_0__inst_mult_20_134 ;
wire Xd_0__inst_mult_20_136 ;
wire Xd_0__inst_mult_20_137 ;
wire Xd_0__inst_mult_20_138 ;
wire Xd_0__inst_mult_21_132 ;
wire Xd_0__inst_mult_21_133 ;
wire Xd_0__inst_mult_21_134 ;
wire Xd_0__inst_mult_21_136 ;
wire Xd_0__inst_mult_21_137 ;
wire Xd_0__inst_mult_21_138 ;
wire Xd_0__inst_mult_18_132 ;
wire Xd_0__inst_mult_18_133 ;
wire Xd_0__inst_mult_18_134 ;
wire Xd_0__inst_mult_18_136 ;
wire Xd_0__inst_mult_18_137 ;
wire Xd_0__inst_mult_18_138 ;
wire Xd_0__inst_mult_19_132 ;
wire Xd_0__inst_mult_19_133 ;
wire Xd_0__inst_mult_19_134 ;
wire Xd_0__inst_mult_19_136 ;
wire Xd_0__inst_mult_19_137 ;
wire Xd_0__inst_mult_19_138 ;
wire Xd_0__inst_mult_16_132 ;
wire Xd_0__inst_mult_16_133 ;
wire Xd_0__inst_mult_16_134 ;
wire Xd_0__inst_mult_16_136 ;
wire Xd_0__inst_mult_16_137 ;
wire Xd_0__inst_mult_16_138 ;
wire Xd_0__inst_mult_17_132 ;
wire Xd_0__inst_mult_17_133 ;
wire Xd_0__inst_mult_17_134 ;
wire Xd_0__inst_mult_17_136 ;
wire Xd_0__inst_mult_17_137 ;
wire Xd_0__inst_mult_17_138 ;
wire Xd_0__inst_mult_14_132 ;
wire Xd_0__inst_mult_14_133 ;
wire Xd_0__inst_mult_14_134 ;
wire Xd_0__inst_mult_14_136 ;
wire Xd_0__inst_mult_14_137 ;
wire Xd_0__inst_mult_14_138 ;
wire Xd_0__inst_mult_15_132 ;
wire Xd_0__inst_mult_15_133 ;
wire Xd_0__inst_mult_15_134 ;
wire Xd_0__inst_mult_15_136 ;
wire Xd_0__inst_mult_15_137 ;
wire Xd_0__inst_mult_15_138 ;
wire Xd_0__inst_mult_12_132 ;
wire Xd_0__inst_mult_12_133 ;
wire Xd_0__inst_mult_12_134 ;
wire Xd_0__inst_mult_12_136 ;
wire Xd_0__inst_mult_12_137 ;
wire Xd_0__inst_mult_12_138 ;
wire Xd_0__inst_mult_13_132 ;
wire Xd_0__inst_mult_13_133 ;
wire Xd_0__inst_mult_13_134 ;
wire Xd_0__inst_mult_13_136 ;
wire Xd_0__inst_mult_13_137 ;
wire Xd_0__inst_mult_13_138 ;
wire Xd_0__inst_mult_10_132 ;
wire Xd_0__inst_mult_10_133 ;
wire Xd_0__inst_mult_10_134 ;
wire Xd_0__inst_mult_10_136 ;
wire Xd_0__inst_mult_10_137 ;
wire Xd_0__inst_mult_10_138 ;
wire Xd_0__inst_mult_11_132 ;
wire Xd_0__inst_mult_11_133 ;
wire Xd_0__inst_mult_11_134 ;
wire Xd_0__inst_mult_11_136 ;
wire Xd_0__inst_mult_11_137 ;
wire Xd_0__inst_mult_11_138 ;
wire Xd_0__inst_mult_8_132 ;
wire Xd_0__inst_mult_8_133 ;
wire Xd_0__inst_mult_8_134 ;
wire Xd_0__inst_mult_8_136 ;
wire Xd_0__inst_mult_8_137 ;
wire Xd_0__inst_mult_8_138 ;
wire Xd_0__inst_mult_9_132 ;
wire Xd_0__inst_mult_9_133 ;
wire Xd_0__inst_mult_9_134 ;
wire Xd_0__inst_mult_9_136 ;
wire Xd_0__inst_mult_9_137 ;
wire Xd_0__inst_mult_9_138 ;
wire Xd_0__inst_mult_6_132 ;
wire Xd_0__inst_mult_6_133 ;
wire Xd_0__inst_mult_6_134 ;
wire Xd_0__inst_mult_6_136 ;
wire Xd_0__inst_mult_6_137 ;
wire Xd_0__inst_mult_6_138 ;
wire Xd_0__inst_mult_7_132 ;
wire Xd_0__inst_mult_7_133 ;
wire Xd_0__inst_mult_7_134 ;
wire Xd_0__inst_mult_7_136 ;
wire Xd_0__inst_mult_7_137 ;
wire Xd_0__inst_mult_7_138 ;
wire Xd_0__inst_mult_4_132 ;
wire Xd_0__inst_mult_4_133 ;
wire Xd_0__inst_mult_4_134 ;
wire Xd_0__inst_mult_4_136 ;
wire Xd_0__inst_mult_4_137 ;
wire Xd_0__inst_mult_4_138 ;
wire Xd_0__inst_mult_5_132 ;
wire Xd_0__inst_mult_5_133 ;
wire Xd_0__inst_mult_5_134 ;
wire Xd_0__inst_mult_5_136 ;
wire Xd_0__inst_mult_5_137 ;
wire Xd_0__inst_mult_5_138 ;
wire Xd_0__inst_mult_2_132 ;
wire Xd_0__inst_mult_2_133 ;
wire Xd_0__inst_mult_2_134 ;
wire Xd_0__inst_mult_2_136 ;
wire Xd_0__inst_mult_2_137 ;
wire Xd_0__inst_mult_2_138 ;
wire Xd_0__inst_mult_3_132 ;
wire Xd_0__inst_mult_3_133 ;
wire Xd_0__inst_mult_3_134 ;
wire Xd_0__inst_mult_3_136 ;
wire Xd_0__inst_mult_3_137 ;
wire Xd_0__inst_mult_3_138 ;
wire Xd_0__inst_mult_0_132 ;
wire Xd_0__inst_mult_0_133 ;
wire Xd_0__inst_mult_0_134 ;
wire Xd_0__inst_mult_0_136 ;
wire Xd_0__inst_mult_0_137 ;
wire Xd_0__inst_mult_0_138 ;
wire Xd_0__inst_mult_1_132 ;
wire Xd_0__inst_mult_1_133 ;
wire Xd_0__inst_mult_1_134 ;
wire Xd_0__inst_mult_1_136 ;
wire Xd_0__inst_mult_1_137 ;
wire Xd_0__inst_mult_1_138 ;
wire Xd_0__inst_mult_28_140 ;
wire Xd_0__inst_mult_28_141 ;
wire Xd_0__inst_mult_28_142 ;
wire Xd_0__inst_mult_28_144 ;
wire Xd_0__inst_mult_28_145 ;
wire Xd_0__inst_mult_28_146 ;
wire Xd_0__inst_mult_29_140 ;
wire Xd_0__inst_mult_29_141 ;
wire Xd_0__inst_mult_29_142 ;
wire Xd_0__inst_mult_29_144 ;
wire Xd_0__inst_mult_29_145 ;
wire Xd_0__inst_mult_29_146 ;
wire Xd_0__inst_mult_26_140 ;
wire Xd_0__inst_mult_26_141 ;
wire Xd_0__inst_mult_26_142 ;
wire Xd_0__inst_mult_26_144 ;
wire Xd_0__inst_mult_26_145 ;
wire Xd_0__inst_mult_26_146 ;
wire Xd_0__inst_mult_27_140 ;
wire Xd_0__inst_mult_27_141 ;
wire Xd_0__inst_mult_27_142 ;
wire Xd_0__inst_mult_27_144 ;
wire Xd_0__inst_mult_27_145 ;
wire Xd_0__inst_mult_27_146 ;
wire Xd_0__inst_mult_24_140 ;
wire Xd_0__inst_mult_24_141 ;
wire Xd_0__inst_mult_24_142 ;
wire Xd_0__inst_mult_24_144 ;
wire Xd_0__inst_mult_24_145 ;
wire Xd_0__inst_mult_24_146 ;
wire Xd_0__inst_mult_25_144 ;
wire Xd_0__inst_mult_25_145 ;
wire Xd_0__inst_mult_25_146 ;
wire Xd_0__inst_mult_22_144 ;
wire Xd_0__inst_mult_22_145 ;
wire Xd_0__inst_mult_22_146 ;
wire Xd_0__inst_mult_23_140 ;
wire Xd_0__inst_mult_23_141 ;
wire Xd_0__inst_mult_23_142 ;
wire Xd_0__inst_mult_23_144 ;
wire Xd_0__inst_mult_23_145 ;
wire Xd_0__inst_mult_23_146 ;
wire Xd_0__inst_mult_20_140 ;
wire Xd_0__inst_mult_20_141 ;
wire Xd_0__inst_mult_20_142 ;
wire Xd_0__inst_mult_20_144 ;
wire Xd_0__inst_mult_20_145 ;
wire Xd_0__inst_mult_20_146 ;
wire Xd_0__inst_mult_21_140 ;
wire Xd_0__inst_mult_21_141 ;
wire Xd_0__inst_mult_21_142 ;
wire Xd_0__inst_mult_21_144 ;
wire Xd_0__inst_mult_21_145 ;
wire Xd_0__inst_mult_21_146 ;
wire Xd_0__inst_mult_18_140 ;
wire Xd_0__inst_mult_18_141 ;
wire Xd_0__inst_mult_18_142 ;
wire Xd_0__inst_mult_18_144 ;
wire Xd_0__inst_mult_18_145 ;
wire Xd_0__inst_mult_18_146 ;
wire Xd_0__inst_mult_19_140 ;
wire Xd_0__inst_mult_19_141 ;
wire Xd_0__inst_mult_19_142 ;
wire Xd_0__inst_mult_19_144 ;
wire Xd_0__inst_mult_19_145 ;
wire Xd_0__inst_mult_19_146 ;
wire Xd_0__inst_mult_16_140 ;
wire Xd_0__inst_mult_16_141 ;
wire Xd_0__inst_mult_16_142 ;
wire Xd_0__inst_mult_16_144 ;
wire Xd_0__inst_mult_16_145 ;
wire Xd_0__inst_mult_16_146 ;
wire Xd_0__inst_mult_17_140 ;
wire Xd_0__inst_mult_17_141 ;
wire Xd_0__inst_mult_17_142 ;
wire Xd_0__inst_mult_17_144 ;
wire Xd_0__inst_mult_17_145 ;
wire Xd_0__inst_mult_17_146 ;
wire Xd_0__inst_mult_14_140 ;
wire Xd_0__inst_mult_14_141 ;
wire Xd_0__inst_mult_14_142 ;
wire Xd_0__inst_mult_14_144 ;
wire Xd_0__inst_mult_14_145 ;
wire Xd_0__inst_mult_14_146 ;
wire Xd_0__inst_mult_15_140 ;
wire Xd_0__inst_mult_15_141 ;
wire Xd_0__inst_mult_15_142 ;
wire Xd_0__inst_mult_15_144 ;
wire Xd_0__inst_mult_15_145 ;
wire Xd_0__inst_mult_15_146 ;
wire Xd_0__inst_mult_12_140 ;
wire Xd_0__inst_mult_12_141 ;
wire Xd_0__inst_mult_12_142 ;
wire Xd_0__inst_mult_12_144 ;
wire Xd_0__inst_mult_12_145 ;
wire Xd_0__inst_mult_12_146 ;
wire Xd_0__inst_mult_13_140 ;
wire Xd_0__inst_mult_13_141 ;
wire Xd_0__inst_mult_13_142 ;
wire Xd_0__inst_mult_13_144 ;
wire Xd_0__inst_mult_13_145 ;
wire Xd_0__inst_mult_13_146 ;
wire Xd_0__inst_mult_10_140 ;
wire Xd_0__inst_mult_10_141 ;
wire Xd_0__inst_mult_10_142 ;
wire Xd_0__inst_mult_10_144 ;
wire Xd_0__inst_mult_10_145 ;
wire Xd_0__inst_mult_10_146 ;
wire Xd_0__inst_mult_11_140 ;
wire Xd_0__inst_mult_11_141 ;
wire Xd_0__inst_mult_11_142 ;
wire Xd_0__inst_mult_11_144 ;
wire Xd_0__inst_mult_11_145 ;
wire Xd_0__inst_mult_11_146 ;
wire Xd_0__inst_mult_8_140 ;
wire Xd_0__inst_mult_8_141 ;
wire Xd_0__inst_mult_8_142 ;
wire Xd_0__inst_mult_8_144 ;
wire Xd_0__inst_mult_8_145 ;
wire Xd_0__inst_mult_8_146 ;
wire Xd_0__inst_mult_9_140 ;
wire Xd_0__inst_mult_9_141 ;
wire Xd_0__inst_mult_9_142 ;
wire Xd_0__inst_mult_9_144 ;
wire Xd_0__inst_mult_9_145 ;
wire Xd_0__inst_mult_9_146 ;
wire Xd_0__inst_mult_6_140 ;
wire Xd_0__inst_mult_6_141 ;
wire Xd_0__inst_mult_6_142 ;
wire Xd_0__inst_mult_6_144 ;
wire Xd_0__inst_mult_6_145 ;
wire Xd_0__inst_mult_6_146 ;
wire Xd_0__inst_mult_7_140 ;
wire Xd_0__inst_mult_7_141 ;
wire Xd_0__inst_mult_7_142 ;
wire Xd_0__inst_mult_7_144 ;
wire Xd_0__inst_mult_7_145 ;
wire Xd_0__inst_mult_7_146 ;
wire Xd_0__inst_mult_4_140 ;
wire Xd_0__inst_mult_4_141 ;
wire Xd_0__inst_mult_4_142 ;
wire Xd_0__inst_mult_4_144 ;
wire Xd_0__inst_mult_4_145 ;
wire Xd_0__inst_mult_4_146 ;
wire Xd_0__inst_mult_5_140 ;
wire Xd_0__inst_mult_5_141 ;
wire Xd_0__inst_mult_5_142 ;
wire Xd_0__inst_mult_5_144 ;
wire Xd_0__inst_mult_5_145 ;
wire Xd_0__inst_mult_5_146 ;
wire Xd_0__inst_mult_2_140 ;
wire Xd_0__inst_mult_2_141 ;
wire Xd_0__inst_mult_2_142 ;
wire Xd_0__inst_mult_2_144 ;
wire Xd_0__inst_mult_2_145 ;
wire Xd_0__inst_mult_2_146 ;
wire Xd_0__inst_mult_3_140 ;
wire Xd_0__inst_mult_3_141 ;
wire Xd_0__inst_mult_3_142 ;
wire Xd_0__inst_mult_3_144 ;
wire Xd_0__inst_mult_3_145 ;
wire Xd_0__inst_mult_3_146 ;
wire Xd_0__inst_mult_0_140 ;
wire Xd_0__inst_mult_0_141 ;
wire Xd_0__inst_mult_0_142 ;
wire Xd_0__inst_mult_0_144 ;
wire Xd_0__inst_mult_0_145 ;
wire Xd_0__inst_mult_0_146 ;
wire Xd_0__inst_mult_1_140 ;
wire Xd_0__inst_mult_1_141 ;
wire Xd_0__inst_mult_1_142 ;
wire Xd_0__inst_mult_1_144 ;
wire Xd_0__inst_mult_1_145 ;
wire Xd_0__inst_mult_1_146 ;
wire Xd_0__inst_mult_28_148 ;
wire Xd_0__inst_mult_28_149 ;
wire Xd_0__inst_mult_28_150 ;
wire Xd_0__inst_mult_29_148 ;
wire Xd_0__inst_mult_29_149 ;
wire Xd_0__inst_mult_29_150 ;
wire Xd_0__inst_mult_26_148 ;
wire Xd_0__inst_mult_26_149 ;
wire Xd_0__inst_mult_26_150 ;
wire Xd_0__inst_mult_27_148 ;
wire Xd_0__inst_mult_27_149 ;
wire Xd_0__inst_mult_27_150 ;
wire Xd_0__inst_mult_24_148 ;
wire Xd_0__inst_mult_24_149 ;
wire Xd_0__inst_mult_24_150 ;
wire Xd_0__inst_mult_25_148 ;
wire Xd_0__inst_mult_25_149 ;
wire Xd_0__inst_mult_25_150 ;
wire Xd_0__inst_mult_22_148 ;
wire Xd_0__inst_mult_22_149 ;
wire Xd_0__inst_mult_22_150 ;
wire Xd_0__inst_mult_23_148 ;
wire Xd_0__inst_mult_23_149 ;
wire Xd_0__inst_mult_23_150 ;
wire Xd_0__inst_mult_20_148 ;
wire Xd_0__inst_mult_20_149 ;
wire Xd_0__inst_mult_20_150 ;
wire Xd_0__inst_mult_21_148 ;
wire Xd_0__inst_mult_21_149 ;
wire Xd_0__inst_mult_21_150 ;
wire Xd_0__inst_mult_18_148 ;
wire Xd_0__inst_mult_18_149 ;
wire Xd_0__inst_mult_18_150 ;
wire Xd_0__inst_mult_19_148 ;
wire Xd_0__inst_mult_19_149 ;
wire Xd_0__inst_mult_19_150 ;
wire Xd_0__inst_mult_16_148 ;
wire Xd_0__inst_mult_16_149 ;
wire Xd_0__inst_mult_16_150 ;
wire Xd_0__inst_mult_17_148 ;
wire Xd_0__inst_mult_17_149 ;
wire Xd_0__inst_mult_17_150 ;
wire Xd_0__inst_mult_14_148 ;
wire Xd_0__inst_mult_14_149 ;
wire Xd_0__inst_mult_14_150 ;
wire Xd_0__inst_mult_15_148 ;
wire Xd_0__inst_mult_15_149 ;
wire Xd_0__inst_mult_15_150 ;
wire Xd_0__inst_mult_12_148 ;
wire Xd_0__inst_mult_12_149 ;
wire Xd_0__inst_mult_12_150 ;
wire Xd_0__inst_mult_13_148 ;
wire Xd_0__inst_mult_13_149 ;
wire Xd_0__inst_mult_13_150 ;
wire Xd_0__inst_mult_10_148 ;
wire Xd_0__inst_mult_10_149 ;
wire Xd_0__inst_mult_10_150 ;
wire Xd_0__inst_mult_11_148 ;
wire Xd_0__inst_mult_11_149 ;
wire Xd_0__inst_mult_11_150 ;
wire Xd_0__inst_mult_8_148 ;
wire Xd_0__inst_mult_8_149 ;
wire Xd_0__inst_mult_8_150 ;
wire Xd_0__inst_mult_9_148 ;
wire Xd_0__inst_mult_9_149 ;
wire Xd_0__inst_mult_9_150 ;
wire Xd_0__inst_mult_6_148 ;
wire Xd_0__inst_mult_6_149 ;
wire Xd_0__inst_mult_6_150 ;
wire Xd_0__inst_mult_7_148 ;
wire Xd_0__inst_mult_7_149 ;
wire Xd_0__inst_mult_7_150 ;
wire Xd_0__inst_mult_4_148 ;
wire Xd_0__inst_mult_4_149 ;
wire Xd_0__inst_mult_4_150 ;
wire Xd_0__inst_mult_5_148 ;
wire Xd_0__inst_mult_5_149 ;
wire Xd_0__inst_mult_5_150 ;
wire Xd_0__inst_mult_2_148 ;
wire Xd_0__inst_mult_2_149 ;
wire Xd_0__inst_mult_2_150 ;
wire Xd_0__inst_mult_3_148 ;
wire Xd_0__inst_mult_3_149 ;
wire Xd_0__inst_mult_3_150 ;
wire Xd_0__inst_mult_0_148 ;
wire Xd_0__inst_mult_0_149 ;
wire Xd_0__inst_mult_0_150 ;
wire Xd_0__inst_mult_1_148 ;
wire Xd_0__inst_mult_1_149 ;
wire Xd_0__inst_mult_1_150 ;
wire Xd_0__inst_mult_28_152 ;
wire Xd_0__inst_mult_29_152 ;
wire Xd_0__inst_mult_26_152 ;
wire Xd_0__inst_mult_27_152 ;
wire Xd_0__inst_mult_24_152 ;
wire Xd_0__inst_mult_25_152 ;
wire Xd_0__inst_mult_22_152 ;
wire Xd_0__inst_mult_23_152 ;
wire Xd_0__inst_mult_20_152 ;
wire Xd_0__inst_mult_21_152 ;
wire Xd_0__inst_mult_18_152 ;
wire Xd_0__inst_mult_19_152 ;
wire Xd_0__inst_mult_16_152 ;
wire Xd_0__inst_mult_17_152 ;
wire Xd_0__inst_mult_14_152 ;
wire Xd_0__inst_mult_15_152 ;
wire Xd_0__inst_mult_12_152 ;
wire Xd_0__inst_mult_13_152 ;
wire Xd_0__inst_mult_10_152 ;
wire Xd_0__inst_mult_11_152 ;
wire Xd_0__inst_mult_8_152 ;
wire Xd_0__inst_mult_9_152 ;
wire Xd_0__inst_mult_6_152 ;
wire Xd_0__inst_mult_7_152 ;
wire Xd_0__inst_mult_4_152 ;
wire Xd_0__inst_mult_5_152 ;
wire Xd_0__inst_mult_2_152 ;
wire Xd_0__inst_mult_3_152 ;
wire Xd_0__inst_mult_0_152 ;
wire Xd_0__inst_mult_1_152 ;
wire Xd_0__inst_mult_28_157 ;
wire Xd_0__inst_mult_28_158 ;
wire Xd_0__inst_mult_29_157 ;
wire Xd_0__inst_mult_29_158 ;
wire Xd_0__inst_mult_26_157 ;
wire Xd_0__inst_mult_26_158 ;
wire Xd_0__inst_mult_27_157 ;
wire Xd_0__inst_mult_27_158 ;
wire Xd_0__inst_mult_24_157 ;
wire Xd_0__inst_mult_24_158 ;
wire Xd_0__inst_mult_25_157 ;
wire Xd_0__inst_mult_25_158 ;
wire Xd_0__inst_mult_22_157 ;
wire Xd_0__inst_mult_22_158 ;
wire Xd_0__inst_mult_23_157 ;
wire Xd_0__inst_mult_23_158 ;
wire Xd_0__inst_mult_20_157 ;
wire Xd_0__inst_mult_20_158 ;
wire Xd_0__inst_mult_21_157 ;
wire Xd_0__inst_mult_21_158 ;
wire Xd_0__inst_mult_18_157 ;
wire Xd_0__inst_mult_18_158 ;
wire Xd_0__inst_mult_19_157 ;
wire Xd_0__inst_mult_19_158 ;
wire Xd_0__inst_mult_30_161 ;
wire Xd_0__inst_mult_30_162 ;
wire Xd_0__inst_mult_31_161 ;
wire Xd_0__inst_mult_31_162 ;
wire Xd_0__inst_mult_16_157 ;
wire Xd_0__inst_mult_16_158 ;
wire Xd_0__inst_mult_17_157 ;
wire Xd_0__inst_mult_17_158 ;
wire Xd_0__inst_mult_14_157 ;
wire Xd_0__inst_mult_14_158 ;
wire Xd_0__inst_mult_15_157 ;
wire Xd_0__inst_mult_15_158 ;
wire Xd_0__inst_mult_12_157 ;
wire Xd_0__inst_mult_12_158 ;
wire Xd_0__inst_mult_13_157 ;
wire Xd_0__inst_mult_13_158 ;
wire Xd_0__inst_mult_10_157 ;
wire Xd_0__inst_mult_10_158 ;
wire Xd_0__inst_mult_11_157 ;
wire Xd_0__inst_mult_11_158 ;
wire Xd_0__inst_mult_8_157 ;
wire Xd_0__inst_mult_8_158 ;
wire Xd_0__inst_mult_9_157 ;
wire Xd_0__inst_mult_9_158 ;
wire Xd_0__inst_mult_6_157 ;
wire Xd_0__inst_mult_6_158 ;
wire Xd_0__inst_mult_7_157 ;
wire Xd_0__inst_mult_7_158 ;
wire Xd_0__inst_mult_4_157 ;
wire Xd_0__inst_mult_4_158 ;
wire Xd_0__inst_mult_5_157 ;
wire Xd_0__inst_mult_5_158 ;
wire Xd_0__inst_mult_2_157 ;
wire Xd_0__inst_mult_2_158 ;
wire Xd_0__inst_mult_3_157 ;
wire Xd_0__inst_mult_3_158 ;
wire Xd_0__inst_mult_0_157 ;
wire Xd_0__inst_mult_0_158 ;
wire Xd_0__inst_mult_1_157 ;
wire Xd_0__inst_mult_1_158 ;
wire Xd_0__inst_mult_28_161 ;
wire Xd_0__inst_mult_28_162 ;
wire Xd_0__inst_mult_29_161 ;
wire Xd_0__inst_mult_29_162 ;
wire Xd_0__inst_mult_26_161 ;
wire Xd_0__inst_mult_26_162 ;
wire Xd_0__inst_mult_27_161 ;
wire Xd_0__inst_mult_27_162 ;
wire Xd_0__inst_mult_24_161 ;
wire Xd_0__inst_mult_24_162 ;
wire Xd_0__inst_mult_25_161 ;
wire Xd_0__inst_mult_25_162 ;
wire Xd_0__inst_mult_22_161 ;
wire Xd_0__inst_mult_22_162 ;
wire Xd_0__inst_mult_23_161 ;
wire Xd_0__inst_mult_23_162 ;
wire Xd_0__inst_mult_20_161 ;
wire Xd_0__inst_mult_20_162 ;
wire Xd_0__inst_mult_21_161 ;
wire Xd_0__inst_mult_21_162 ;
wire Xd_0__inst_mult_18_161 ;
wire Xd_0__inst_mult_18_162 ;
wire Xd_0__inst_mult_19_161 ;
wire Xd_0__inst_mult_19_162 ;
wire Xd_0__inst_mult_16_161 ;
wire Xd_0__inst_mult_16_162 ;
wire Xd_0__inst_mult_17_161 ;
wire Xd_0__inst_mult_17_162 ;
wire Xd_0__inst_mult_14_161 ;
wire Xd_0__inst_mult_14_162 ;
wire Xd_0__inst_mult_15_161 ;
wire Xd_0__inst_mult_15_162 ;
wire Xd_0__inst_mult_12_161 ;
wire Xd_0__inst_mult_12_162 ;
wire Xd_0__inst_mult_13_161 ;
wire Xd_0__inst_mult_13_162 ;
wire Xd_0__inst_mult_10_161 ;
wire Xd_0__inst_mult_10_162 ;
wire Xd_0__inst_mult_11_161 ;
wire Xd_0__inst_mult_11_162 ;
wire Xd_0__inst_mult_8_161 ;
wire Xd_0__inst_mult_8_162 ;
wire Xd_0__inst_mult_9_161 ;
wire Xd_0__inst_mult_9_162 ;
wire Xd_0__inst_mult_6_161 ;
wire Xd_0__inst_mult_6_162 ;
wire Xd_0__inst_mult_7_161 ;
wire Xd_0__inst_mult_7_162 ;
wire Xd_0__inst_mult_4_161 ;
wire Xd_0__inst_mult_4_162 ;
wire Xd_0__inst_mult_5_161 ;
wire Xd_0__inst_mult_5_162 ;
wire Xd_0__inst_mult_2_161 ;
wire Xd_0__inst_mult_2_162 ;
wire Xd_0__inst_mult_3_161 ;
wire Xd_0__inst_mult_3_162 ;
wire Xd_0__inst_mult_0_161 ;
wire Xd_0__inst_mult_0_162 ;
wire Xd_0__inst_mult_1_161 ;
wire Xd_0__inst_mult_1_162 ;
wire Xd_0__inst_inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_first_level_4__0__q ;
wire Xd_0__inst_inst_first_level_3__0__q ;
wire Xd_0__inst_inst_first_level_5__0__q ;
wire Xd_0__inst_inst_first_level_2__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_4__1__q ;
wire Xd_0__inst_inst_first_level_3__1__q ;
wire Xd_0__inst_inst_first_level_5__1__q ;
wire Xd_0__inst_inst_first_level_2__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_4__2__q ;
wire Xd_0__inst_inst_first_level_3__2__q ;
wire Xd_0__inst_inst_first_level_5__2__q ;
wire Xd_0__inst_inst_first_level_2__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_4__3__q ;
wire Xd_0__inst_inst_first_level_3__3__q ;
wire Xd_0__inst_inst_first_level_5__3__q ;
wire Xd_0__inst_inst_first_level_2__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_4__4__q ;
wire Xd_0__inst_inst_first_level_3__4__q ;
wire Xd_0__inst_inst_first_level_5__4__q ;
wire Xd_0__inst_inst_first_level_2__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_4__5__q ;
wire Xd_0__inst_inst_first_level_3__5__q ;
wire Xd_0__inst_inst_first_level_5__5__q ;
wire Xd_0__inst_inst_first_level_2__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_4__6__q ;
wire Xd_0__inst_inst_first_level_3__6__q ;
wire Xd_0__inst_inst_first_level_5__6__q ;
wire Xd_0__inst_inst_first_level_2__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_4__7__q ;
wire Xd_0__inst_inst_first_level_3__7__q ;
wire Xd_0__inst_inst_first_level_5__7__q ;
wire Xd_0__inst_inst_first_level_2__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_4__8__q ;
wire Xd_0__inst_inst_first_level_3__8__q ;
wire Xd_0__inst_inst_first_level_5__8__q ;
wire Xd_0__inst_inst_first_level_2__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_4__9__q ;
wire Xd_0__inst_inst_first_level_3__9__q ;
wire Xd_0__inst_inst_first_level_5__9__q ;
wire Xd_0__inst_inst_first_level_2__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_4__10__q ;
wire Xd_0__inst_inst_first_level_3__10__q ;
wire Xd_0__inst_inst_first_level_5__10__q ;
wire Xd_0__inst_inst_first_level_2__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_4__11__q ;
wire Xd_0__inst_inst_first_level_3__11__q ;
wire Xd_0__inst_inst_first_level_5__11__q ;
wire Xd_0__inst_inst_first_level_2__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_4__12__q ;
wire Xd_0__inst_inst_first_level_3__12__q ;
wire Xd_0__inst_inst_first_level_5__12__q ;
wire Xd_0__inst_inst_first_level_2__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_4__13__q ;
wire Xd_0__inst_inst_first_level_3__13__q ;
wire Xd_0__inst_inst_first_level_5__15__q ;
wire Xd_0__inst_inst_first_level_2__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_4__14__q ;
wire Xd_0__inst_inst_first_level_3__14__q ;
wire Xd_0__inst_inst_first_level_2__14__q ;
wire Xd_0__inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_first_level_4__15__q ;
wire Xd_0__inst_inst_first_level_3__15__q ;
wire Xd_0__inst_inst_first_level_2__15__q ;
wire Xd_0__inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_0__15__q ;
wire Xd_0__inst_r_sum1_15__0__q ;
wire Xd_0__inst_r_sum1_15__1__q ;
wire Xd_0__inst_r_sum1_15__2__q ;
wire Xd_0__inst_r_sum1_15__3__q ;
wire Xd_0__inst_r_sum1_15__4__q ;
wire Xd_0__inst_r_sum1_15__5__q ;
wire Xd_0__inst_r_sum1_15__6__q ;
wire Xd_0__inst_r_sum1_15__7__q ;
wire Xd_0__inst_r_sum1_15__8__q ;
wire Xd_0__inst_r_sum1_15__9__q ;
wire Xd_0__inst_r_sum1_15__10__q ;
wire Xd_0__inst_r_sum1_15__11__q ;
wire Xd_0__inst_r_sum1_15__12__q ;
wire Xd_0__inst_r_sum1_15__13__q ;
wire Xd_0__inst_r_sum1_14__0__q ;
wire Xd_0__inst_r_sum1_13__0__q ;
wire Xd_0__inst_r_sum1_12__0__q ;
wire Xd_0__inst_r_sum1_11__0__q ;
wire Xd_0__inst_r_sum1_10__0__q ;
wire Xd_0__inst_r_sum1_9__0__q ;
wire Xd_0__inst_r_sum1_8__0__q ;
wire Xd_0__inst_r_sum1_7__0__q ;
wire Xd_0__inst_r_sum1_6__0__q ;
wire Xd_0__inst_r_sum1_5__0__q ;
wire Xd_0__inst_r_sum1_4__0__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_14__1__q ;
wire Xd_0__inst_r_sum1_13__1__q ;
wire Xd_0__inst_r_sum1_12__1__q ;
wire Xd_0__inst_r_sum1_11__1__q ;
wire Xd_0__inst_r_sum1_10__1__q ;
wire Xd_0__inst_r_sum1_9__1__q ;
wire Xd_0__inst_r_sum1_8__1__q ;
wire Xd_0__inst_r_sum1_7__1__q ;
wire Xd_0__inst_r_sum1_6__1__q ;
wire Xd_0__inst_r_sum1_5__1__q ;
wire Xd_0__inst_r_sum1_4__1__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_14__2__q ;
wire Xd_0__inst_r_sum1_13__2__q ;
wire Xd_0__inst_r_sum1_12__2__q ;
wire Xd_0__inst_r_sum1_11__2__q ;
wire Xd_0__inst_r_sum1_10__2__q ;
wire Xd_0__inst_r_sum1_9__2__q ;
wire Xd_0__inst_r_sum1_8__2__q ;
wire Xd_0__inst_r_sum1_7__2__q ;
wire Xd_0__inst_r_sum1_6__2__q ;
wire Xd_0__inst_r_sum1_5__2__q ;
wire Xd_0__inst_r_sum1_4__2__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_14__3__q ;
wire Xd_0__inst_r_sum1_13__3__q ;
wire Xd_0__inst_r_sum1_12__3__q ;
wire Xd_0__inst_r_sum1_11__3__q ;
wire Xd_0__inst_r_sum1_10__3__q ;
wire Xd_0__inst_r_sum1_9__3__q ;
wire Xd_0__inst_r_sum1_8__3__q ;
wire Xd_0__inst_r_sum1_7__3__q ;
wire Xd_0__inst_r_sum1_6__3__q ;
wire Xd_0__inst_r_sum1_5__3__q ;
wire Xd_0__inst_r_sum1_4__3__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_14__4__q ;
wire Xd_0__inst_r_sum1_13__4__q ;
wire Xd_0__inst_r_sum1_12__4__q ;
wire Xd_0__inst_r_sum1_11__4__q ;
wire Xd_0__inst_r_sum1_10__4__q ;
wire Xd_0__inst_r_sum1_9__4__q ;
wire Xd_0__inst_r_sum1_8__4__q ;
wire Xd_0__inst_r_sum1_7__4__q ;
wire Xd_0__inst_r_sum1_6__4__q ;
wire Xd_0__inst_r_sum1_5__4__q ;
wire Xd_0__inst_r_sum1_4__4__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_14__5__q ;
wire Xd_0__inst_r_sum1_13__5__q ;
wire Xd_0__inst_r_sum1_12__5__q ;
wire Xd_0__inst_r_sum1_11__5__q ;
wire Xd_0__inst_r_sum1_10__5__q ;
wire Xd_0__inst_r_sum1_9__5__q ;
wire Xd_0__inst_r_sum1_8__5__q ;
wire Xd_0__inst_r_sum1_7__5__q ;
wire Xd_0__inst_r_sum1_6__5__q ;
wire Xd_0__inst_r_sum1_5__5__q ;
wire Xd_0__inst_r_sum1_4__5__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_14__6__q ;
wire Xd_0__inst_r_sum1_13__6__q ;
wire Xd_0__inst_r_sum1_12__6__q ;
wire Xd_0__inst_r_sum1_11__6__q ;
wire Xd_0__inst_r_sum1_10__6__q ;
wire Xd_0__inst_r_sum1_9__6__q ;
wire Xd_0__inst_r_sum1_8__6__q ;
wire Xd_0__inst_r_sum1_7__6__q ;
wire Xd_0__inst_r_sum1_6__6__q ;
wire Xd_0__inst_r_sum1_5__6__q ;
wire Xd_0__inst_r_sum1_4__6__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_14__7__q ;
wire Xd_0__inst_r_sum1_13__7__q ;
wire Xd_0__inst_r_sum1_12__7__q ;
wire Xd_0__inst_r_sum1_11__7__q ;
wire Xd_0__inst_r_sum1_10__7__q ;
wire Xd_0__inst_r_sum1_9__7__q ;
wire Xd_0__inst_r_sum1_8__7__q ;
wire Xd_0__inst_r_sum1_7__7__q ;
wire Xd_0__inst_r_sum1_6__7__q ;
wire Xd_0__inst_r_sum1_5__7__q ;
wire Xd_0__inst_r_sum1_4__7__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_14__8__q ;
wire Xd_0__inst_r_sum1_13__8__q ;
wire Xd_0__inst_r_sum1_12__8__q ;
wire Xd_0__inst_r_sum1_11__8__q ;
wire Xd_0__inst_r_sum1_10__8__q ;
wire Xd_0__inst_r_sum1_9__8__q ;
wire Xd_0__inst_r_sum1_8__8__q ;
wire Xd_0__inst_r_sum1_7__8__q ;
wire Xd_0__inst_r_sum1_6__8__q ;
wire Xd_0__inst_r_sum1_5__8__q ;
wire Xd_0__inst_r_sum1_4__8__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_14__9__q ;
wire Xd_0__inst_r_sum1_13__9__q ;
wire Xd_0__inst_r_sum1_12__9__q ;
wire Xd_0__inst_r_sum1_11__9__q ;
wire Xd_0__inst_r_sum1_10__9__q ;
wire Xd_0__inst_r_sum1_9__9__q ;
wire Xd_0__inst_r_sum1_8__9__q ;
wire Xd_0__inst_r_sum1_7__9__q ;
wire Xd_0__inst_r_sum1_6__9__q ;
wire Xd_0__inst_r_sum1_5__9__q ;
wire Xd_0__inst_r_sum1_4__9__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_14__10__q ;
wire Xd_0__inst_r_sum1_13__10__q ;
wire Xd_0__inst_r_sum1_12__10__q ;
wire Xd_0__inst_r_sum1_11__10__q ;
wire Xd_0__inst_r_sum1_10__10__q ;
wire Xd_0__inst_r_sum1_9__10__q ;
wire Xd_0__inst_r_sum1_8__10__q ;
wire Xd_0__inst_r_sum1_7__10__q ;
wire Xd_0__inst_r_sum1_6__10__q ;
wire Xd_0__inst_r_sum1_5__10__q ;
wire Xd_0__inst_r_sum1_4__10__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_14__11__q ;
wire Xd_0__inst_r_sum1_13__11__q ;
wire Xd_0__inst_r_sum1_12__11__q ;
wire Xd_0__inst_r_sum1_11__11__q ;
wire Xd_0__inst_r_sum1_10__11__q ;
wire Xd_0__inst_r_sum1_9__11__q ;
wire Xd_0__inst_r_sum1_8__11__q ;
wire Xd_0__inst_r_sum1_7__11__q ;
wire Xd_0__inst_r_sum1_6__11__q ;
wire Xd_0__inst_r_sum1_5__11__q ;
wire Xd_0__inst_r_sum1_4__11__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_14__12__q ;
wire Xd_0__inst_r_sum1_13__12__q ;
wire Xd_0__inst_r_sum1_12__12__q ;
wire Xd_0__inst_r_sum1_11__12__q ;
wire Xd_0__inst_r_sum1_10__12__q ;
wire Xd_0__inst_r_sum1_9__12__q ;
wire Xd_0__inst_r_sum1_8__12__q ;
wire Xd_0__inst_r_sum1_7__12__q ;
wire Xd_0__inst_r_sum1_6__12__q ;
wire Xd_0__inst_r_sum1_5__12__q ;
wire Xd_0__inst_r_sum1_4__12__q ;
wire Xd_0__inst_r_sum1_3__12__q ;
wire Xd_0__inst_r_sum1_2__12__q ;
wire Xd_0__inst_r_sum1_1__12__q ;
wire Xd_0__inst_r_sum1_0__12__q ;
wire Xd_0__inst_r_sum1_14__13__q ;
wire Xd_0__inst_r_sum1_13__13__q ;
wire Xd_0__inst_r_sum1_12__13__q ;
wire Xd_0__inst_r_sum1_11__13__q ;
wire Xd_0__inst_r_sum1_10__13__q ;
wire Xd_0__inst_r_sum1_9__13__q ;
wire Xd_0__inst_r_sum1_8__13__q ;
wire Xd_0__inst_r_sum1_7__13__q ;
wire Xd_0__inst_r_sum1_6__13__q ;
wire Xd_0__inst_r_sum1_5__13__q ;
wire Xd_0__inst_r_sum1_4__13__q ;
wire Xd_0__inst_r_sum1_3__13__q ;
wire Xd_0__inst_r_sum1_2__13__q ;
wire Xd_0__inst_r_sum1_1__13__q ;
wire Xd_0__inst_r_sum1_0__13__q ;
wire Xd_0__inst_product_30__0__q ;
wire Xd_0__inst_product_31__0__q ;
wire Xd_0__inst_product_30__1__q ;
wire Xd_0__inst_product_31__1__q ;
wire Xd_0__inst_product_30__2__q ;
wire Xd_0__inst_product_31__2__q ;
wire Xd_0__inst_product_30__3__q ;
wire Xd_0__inst_product_31__3__q ;
wire Xd_0__inst_product_30__4__q ;
wire Xd_0__inst_product_31__4__q ;
wire Xd_0__inst_product_30__5__q ;
wire Xd_0__inst_product_31__5__q ;
wire Xd_0__inst_product_30__6__q ;
wire Xd_0__inst_product_31__6__q ;
wire Xd_0__inst_product_30__7__q ;
wire Xd_0__inst_product_31__7__q ;
wire Xd_0__inst_product_30__8__q ;
wire Xd_0__inst_product_31__8__q ;
wire Xd_0__inst_product_30__9__q ;
wire Xd_0__inst_product_31__9__q ;
wire Xd_0__inst_product_30__10__q ;
wire Xd_0__inst_product_31__10__q ;
wire Xd_0__inst_product_30__11__q ;
wire Xd_0__inst_product_31__11__q ;
wire Xd_0__inst_product_28__0__q ;
wire Xd_0__inst_product_29__0__q ;
wire Xd_0__inst_product_26__0__q ;
wire Xd_0__inst_product_27__0__q ;
wire Xd_0__inst_product_24__0__q ;
wire Xd_0__inst_product_25__0__q ;
wire Xd_0__inst_product_22__0__q ;
wire Xd_0__inst_product_23__0__q ;
wire Xd_0__inst_product_20__0__q ;
wire Xd_0__inst_product_21__0__q ;
wire Xd_0__inst_product_18__0__q ;
wire Xd_0__inst_product_19__0__q ;
wire Xd_0__inst_product1_30__0__q ;
wire Xd_0__inst_product1_31__0__q ;
wire Xd_0__inst_product_16__0__q ;
wire Xd_0__inst_product_17__0__q ;
wire Xd_0__inst_product_14__0__q ;
wire Xd_0__inst_product_15__0__q ;
wire Xd_0__inst_product_12__0__q ;
wire Xd_0__inst_product_13__0__q ;
wire Xd_0__inst_product_10__0__q ;
wire Xd_0__inst_product_11__0__q ;
wire Xd_0__inst_product_8__0__q ;
wire Xd_0__inst_product_9__0__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product_28__1__q ;
wire Xd_0__inst_product_29__1__q ;
wire Xd_0__inst_product_26__1__q ;
wire Xd_0__inst_product_27__1__q ;
wire Xd_0__inst_product_24__1__q ;
wire Xd_0__inst_product_25__1__q ;
wire Xd_0__inst_product_22__1__q ;
wire Xd_0__inst_product_23__1__q ;
wire Xd_0__inst_product_20__1__q ;
wire Xd_0__inst_product_21__1__q ;
wire Xd_0__inst_product_18__1__q ;
wire Xd_0__inst_product_19__1__q ;
wire Xd_0__inst_product1_30__1__q ;
wire Xd_0__inst_product1_31__1__q ;
wire Xd_0__inst_product_16__1__q ;
wire Xd_0__inst_product_17__1__q ;
wire Xd_0__inst_product_14__1__q ;
wire Xd_0__inst_product_15__1__q ;
wire Xd_0__inst_product_12__1__q ;
wire Xd_0__inst_product_13__1__q ;
wire Xd_0__inst_product_10__1__q ;
wire Xd_0__inst_product_11__1__q ;
wire Xd_0__inst_product_8__1__q ;
wire Xd_0__inst_product_9__1__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product_28__2__q ;
wire Xd_0__inst_product_29__2__q ;
wire Xd_0__inst_product_26__2__q ;
wire Xd_0__inst_product_27__2__q ;
wire Xd_0__inst_product_24__2__q ;
wire Xd_0__inst_product_25__2__q ;
wire Xd_0__inst_product_22__2__q ;
wire Xd_0__inst_product_23__2__q ;
wire Xd_0__inst_product_20__2__q ;
wire Xd_0__inst_product_21__2__q ;
wire Xd_0__inst_product_18__2__q ;
wire Xd_0__inst_product_19__2__q ;
wire Xd_0__inst_product1_30__2__q ;
wire Xd_0__inst_product1_31__2__q ;
wire Xd_0__inst_product_16__2__q ;
wire Xd_0__inst_product_17__2__q ;
wire Xd_0__inst_product_14__2__q ;
wire Xd_0__inst_product_15__2__q ;
wire Xd_0__inst_product_12__2__q ;
wire Xd_0__inst_product_13__2__q ;
wire Xd_0__inst_product_10__2__q ;
wire Xd_0__inst_product_11__2__q ;
wire Xd_0__inst_product_8__2__q ;
wire Xd_0__inst_product_9__2__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product_28__3__q ;
wire Xd_0__inst_product_29__3__q ;
wire Xd_0__inst_product_26__3__q ;
wire Xd_0__inst_product_27__3__q ;
wire Xd_0__inst_product_24__3__q ;
wire Xd_0__inst_product_25__3__q ;
wire Xd_0__inst_product_22__3__q ;
wire Xd_0__inst_product_23__3__q ;
wire Xd_0__inst_product_20__3__q ;
wire Xd_0__inst_product_21__3__q ;
wire Xd_0__inst_product_18__3__q ;
wire Xd_0__inst_product_19__3__q ;
wire Xd_0__inst_product_16__3__q ;
wire Xd_0__inst_product_17__3__q ;
wire Xd_0__inst_product_14__3__q ;
wire Xd_0__inst_product_15__3__q ;
wire Xd_0__inst_product_12__3__q ;
wire Xd_0__inst_product_13__3__q ;
wire Xd_0__inst_product_10__3__q ;
wire Xd_0__inst_product_11__3__q ;
wire Xd_0__inst_product_8__3__q ;
wire Xd_0__inst_product_9__3__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product_28__4__q ;
wire Xd_0__inst_product_29__4__q ;
wire Xd_0__inst_product_26__4__q ;
wire Xd_0__inst_product_27__4__q ;
wire Xd_0__inst_product_24__4__q ;
wire Xd_0__inst_product_25__4__q ;
wire Xd_0__inst_product_22__4__q ;
wire Xd_0__inst_product_23__4__q ;
wire Xd_0__inst_product_20__4__q ;
wire Xd_0__inst_product_21__4__q ;
wire Xd_0__inst_product_18__4__q ;
wire Xd_0__inst_product_19__4__q ;
wire Xd_0__inst_product_16__4__q ;
wire Xd_0__inst_product_17__4__q ;
wire Xd_0__inst_product_14__4__q ;
wire Xd_0__inst_product_15__4__q ;
wire Xd_0__inst_product_12__4__q ;
wire Xd_0__inst_product_13__4__q ;
wire Xd_0__inst_product_10__4__q ;
wire Xd_0__inst_product_11__4__q ;
wire Xd_0__inst_product_8__4__q ;
wire Xd_0__inst_product_9__4__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product_28__5__q ;
wire Xd_0__inst_product_29__5__q ;
wire Xd_0__inst_product_26__5__q ;
wire Xd_0__inst_product_27__5__q ;
wire Xd_0__inst_product_24__5__q ;
wire Xd_0__inst_product_25__5__q ;
wire Xd_0__inst_product_22__5__q ;
wire Xd_0__inst_product_23__5__q ;
wire Xd_0__inst_product_20__5__q ;
wire Xd_0__inst_product_21__5__q ;
wire Xd_0__inst_product_18__5__q ;
wire Xd_0__inst_product_19__5__q ;
wire Xd_0__inst_product_16__5__q ;
wire Xd_0__inst_product_17__5__q ;
wire Xd_0__inst_product_14__5__q ;
wire Xd_0__inst_product_15__5__q ;
wire Xd_0__inst_product_12__5__q ;
wire Xd_0__inst_product_13__5__q ;
wire Xd_0__inst_product_10__5__q ;
wire Xd_0__inst_product_11__5__q ;
wire Xd_0__inst_product_8__5__q ;
wire Xd_0__inst_product_9__5__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_28__6__q ;
wire Xd_0__inst_product_29__6__q ;
wire Xd_0__inst_product_26__6__q ;
wire Xd_0__inst_product_27__6__q ;
wire Xd_0__inst_product_24__6__q ;
wire Xd_0__inst_product_25__6__q ;
wire Xd_0__inst_product_22__6__q ;
wire Xd_0__inst_product_23__6__q ;
wire Xd_0__inst_product_20__6__q ;
wire Xd_0__inst_product_21__6__q ;
wire Xd_0__inst_product_18__6__q ;
wire Xd_0__inst_product_19__6__q ;
wire Xd_0__inst_product_16__6__q ;
wire Xd_0__inst_product_17__6__q ;
wire Xd_0__inst_product_14__6__q ;
wire Xd_0__inst_product_15__6__q ;
wire Xd_0__inst_product_12__6__q ;
wire Xd_0__inst_product_13__6__q ;
wire Xd_0__inst_product_10__6__q ;
wire Xd_0__inst_product_11__6__q ;
wire Xd_0__inst_product_8__6__q ;
wire Xd_0__inst_product_9__6__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_28__7__q ;
wire Xd_0__inst_product_29__7__q ;
wire Xd_0__inst_product_26__7__q ;
wire Xd_0__inst_product_27__7__q ;
wire Xd_0__inst_product_24__7__q ;
wire Xd_0__inst_product_25__7__q ;
wire Xd_0__inst_product_22__7__q ;
wire Xd_0__inst_product_23__7__q ;
wire Xd_0__inst_product_20__7__q ;
wire Xd_0__inst_product_21__7__q ;
wire Xd_0__inst_product_18__7__q ;
wire Xd_0__inst_product_19__7__q ;
wire Xd_0__inst_product_16__7__q ;
wire Xd_0__inst_product_17__7__q ;
wire Xd_0__inst_product_14__7__q ;
wire Xd_0__inst_product_15__7__q ;
wire Xd_0__inst_product_12__7__q ;
wire Xd_0__inst_product_13__7__q ;
wire Xd_0__inst_product_10__7__q ;
wire Xd_0__inst_product_11__7__q ;
wire Xd_0__inst_product_8__7__q ;
wire Xd_0__inst_product_9__7__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_28__8__q ;
wire Xd_0__inst_product_29__8__q ;
wire Xd_0__inst_product_26__8__q ;
wire Xd_0__inst_product_27__8__q ;
wire Xd_0__inst_product_24__8__q ;
wire Xd_0__inst_product_25__8__q ;
wire Xd_0__inst_product_22__8__q ;
wire Xd_0__inst_product_23__8__q ;
wire Xd_0__inst_product_20__8__q ;
wire Xd_0__inst_product_21__8__q ;
wire Xd_0__inst_product_18__8__q ;
wire Xd_0__inst_product_19__8__q ;
wire Xd_0__inst_product_16__8__q ;
wire Xd_0__inst_product_17__8__q ;
wire Xd_0__inst_product_14__8__q ;
wire Xd_0__inst_product_15__8__q ;
wire Xd_0__inst_product_12__8__q ;
wire Xd_0__inst_product_13__8__q ;
wire Xd_0__inst_product_10__8__q ;
wire Xd_0__inst_product_11__8__q ;
wire Xd_0__inst_product_8__8__q ;
wire Xd_0__inst_product_9__8__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_28__9__q ;
wire Xd_0__inst_product_29__9__q ;
wire Xd_0__inst_product_26__9__q ;
wire Xd_0__inst_product_27__9__q ;
wire Xd_0__inst_product_24__9__q ;
wire Xd_0__inst_product_25__9__q ;
wire Xd_0__inst_product_22__9__q ;
wire Xd_0__inst_product_23__9__q ;
wire Xd_0__inst_product_20__9__q ;
wire Xd_0__inst_product_21__9__q ;
wire Xd_0__inst_product_18__9__q ;
wire Xd_0__inst_product_19__9__q ;
wire Xd_0__inst_product_16__9__q ;
wire Xd_0__inst_product_17__9__q ;
wire Xd_0__inst_product_14__9__q ;
wire Xd_0__inst_product_15__9__q ;
wire Xd_0__inst_product_12__9__q ;
wire Xd_0__inst_product_13__9__q ;
wire Xd_0__inst_product_10__9__q ;
wire Xd_0__inst_product_11__9__q ;
wire Xd_0__inst_product_8__9__q ;
wire Xd_0__inst_product_9__9__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_28__10__q ;
wire Xd_0__inst_product_29__10__q ;
wire Xd_0__inst_product_26__10__q ;
wire Xd_0__inst_product_27__10__q ;
wire Xd_0__inst_product_24__10__q ;
wire Xd_0__inst_product_25__10__q ;
wire Xd_0__inst_product_22__10__q ;
wire Xd_0__inst_product_23__10__q ;
wire Xd_0__inst_product_20__10__q ;
wire Xd_0__inst_product_21__10__q ;
wire Xd_0__inst_product_18__10__q ;
wire Xd_0__inst_product_19__10__q ;
wire Xd_0__inst_product_16__10__q ;
wire Xd_0__inst_product_17__10__q ;
wire Xd_0__inst_product_14__10__q ;
wire Xd_0__inst_product_15__10__q ;
wire Xd_0__inst_product_12__10__q ;
wire Xd_0__inst_product_13__10__q ;
wire Xd_0__inst_product_10__10__q ;
wire Xd_0__inst_product_11__10__q ;
wire Xd_0__inst_product_8__10__q ;
wire Xd_0__inst_product_9__10__q ;
wire Xd_0__inst_product_6__10__q ;
wire Xd_0__inst_product_7__10__q ;
wire Xd_0__inst_product_4__10__q ;
wire Xd_0__inst_product_5__10__q ;
wire Xd_0__inst_product_2__10__q ;
wire Xd_0__inst_product_3__10__q ;
wire Xd_0__inst_product_0__10__q ;
wire Xd_0__inst_product_1__10__q ;
wire Xd_0__inst_product_28__11__q ;
wire Xd_0__inst_product_29__11__q ;
wire Xd_0__inst_product_26__11__q ;
wire Xd_0__inst_product_27__11__q ;
wire Xd_0__inst_product_24__11__q ;
wire Xd_0__inst_product_25__11__q ;
wire Xd_0__inst_product_22__11__q ;
wire Xd_0__inst_product_23__11__q ;
wire Xd_0__inst_product_20__11__q ;
wire Xd_0__inst_product_21__11__q ;
wire Xd_0__inst_product_18__11__q ;
wire Xd_0__inst_product_19__11__q ;
wire Xd_0__inst_product_16__11__q ;
wire Xd_0__inst_product_17__11__q ;
wire Xd_0__inst_product_14__11__q ;
wire Xd_0__inst_product_15__11__q ;
wire Xd_0__inst_product_12__11__q ;
wire Xd_0__inst_product_13__11__q ;
wire Xd_0__inst_product_10__11__q ;
wire Xd_0__inst_product_11__11__q ;
wire Xd_0__inst_product_8__11__q ;
wire Xd_0__inst_product_9__11__q ;
wire Xd_0__inst_product_6__11__q ;
wire Xd_0__inst_product_7__11__q ;
wire Xd_0__inst_product_4__11__q ;
wire Xd_0__inst_product_5__11__q ;
wire Xd_0__inst_product_2__11__q ;
wire Xd_0__inst_product_3__11__q ;
wire Xd_0__inst_product_0__11__q ;
wire Xd_0__inst_product_1__11__q ;
wire Xd_0__inst_product1_28__0__q ;
wire Xd_0__inst_product1_29__0__q ;
wire Xd_0__inst_product1_26__0__q ;
wire Xd_0__inst_product1_27__0__q ;
wire Xd_0__inst_product1_24__0__q ;
wire Xd_0__inst_product1_25__0__q ;
wire Xd_0__inst_product1_22__0__q ;
wire Xd_0__inst_product1_23__0__q ;
wire Xd_0__inst_product1_20__0__q ;
wire Xd_0__inst_product1_21__0__q ;
wire Xd_0__inst_product1_18__0__q ;
wire Xd_0__inst_product1_19__0__q ;
wire Xd_0__inst_product1_16__0__q ;
wire Xd_0__inst_product1_17__0__q ;
wire Xd_0__inst_product1_14__0__q ;
wire Xd_0__inst_product1_15__0__q ;
wire Xd_0__inst_product1_12__0__q ;
wire Xd_0__inst_product1_13__0__q ;
wire Xd_0__inst_product1_10__0__q ;
wire Xd_0__inst_product1_11__0__q ;
wire Xd_0__inst_product1_8__0__q ;
wire Xd_0__inst_product1_9__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_28__1__q ;
wire Xd_0__inst_product1_29__1__q ;
wire Xd_0__inst_product1_26__1__q ;
wire Xd_0__inst_product1_27__1__q ;
wire Xd_0__inst_product1_24__1__q ;
wire Xd_0__inst_product1_25__1__q ;
wire Xd_0__inst_product1_22__1__q ;
wire Xd_0__inst_product1_23__1__q ;
wire Xd_0__inst_product1_20__1__q ;
wire Xd_0__inst_product1_21__1__q ;
wire Xd_0__inst_product1_18__1__q ;
wire Xd_0__inst_product1_19__1__q ;
wire Xd_0__inst_product1_16__1__q ;
wire Xd_0__inst_product1_17__1__q ;
wire Xd_0__inst_product1_14__1__q ;
wire Xd_0__inst_product1_15__1__q ;
wire Xd_0__inst_product1_12__1__q ;
wire Xd_0__inst_product1_13__1__q ;
wire Xd_0__inst_product1_10__1__q ;
wire Xd_0__inst_product1_11__1__q ;
wire Xd_0__inst_product1_8__1__q ;
wire Xd_0__inst_product1_9__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_28__2__q ;
wire Xd_0__inst_product1_29__2__q ;
wire Xd_0__inst_product1_26__2__q ;
wire Xd_0__inst_product1_27__2__q ;
wire Xd_0__inst_product1_24__2__q ;
wire Xd_0__inst_product1_25__2__q ;
wire Xd_0__inst_product1_22__2__q ;
wire Xd_0__inst_product1_23__2__q ;
wire Xd_0__inst_product1_20__2__q ;
wire Xd_0__inst_product1_21__2__q ;
wire Xd_0__inst_product1_18__2__q ;
wire Xd_0__inst_product1_19__2__q ;
wire Xd_0__inst_product1_16__2__q ;
wire Xd_0__inst_product1_17__2__q ;
wire Xd_0__inst_product1_14__2__q ;
wire Xd_0__inst_product1_15__2__q ;
wire Xd_0__inst_product1_12__2__q ;
wire Xd_0__inst_product1_13__2__q ;
wire Xd_0__inst_product1_10__2__q ;
wire Xd_0__inst_product1_11__2__q ;
wire Xd_0__inst_product1_8__2__q ;
wire Xd_0__inst_product1_9__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_mult_30_2_q ;
wire Xd_0__inst_mult_30_3_q ;
wire Xd_0__inst_mult_30_4_q ;
wire Xd_0__inst_mult_31_2_q ;
wire Xd_0__inst_mult_31_3_q ;
wire Xd_0__inst_mult_31_4_q ;
wire Xd_0__inst_mult_30_5_q ;
wire Xd_0__inst_mult_30_6_q ;
wire Xd_0__inst_mult_30_7_q ;
wire Xd_0__inst_mult_31_5_q ;
wire Xd_0__inst_mult_31_6_q ;
wire Xd_0__inst_mult_31_7_q ;
wire Xd_0__inst_mult_30_8_q ;
wire Xd_0__inst_mult_30_9_q ;
wire Xd_0__inst_mult_31_8_q ;
wire Xd_0__inst_mult_31_9_q ;
wire Xd_0__inst_mult_30_10_q ;
wire Xd_0__inst_mult_30_11_q ;
wire Xd_0__inst_mult_30_1_q ;
wire Xd_0__inst_mult_31_10_q ;
wire Xd_0__inst_mult_31_11_q ;
wire Xd_0__inst_mult_31_1_q ;
wire Xd_0__inst_mult_30_12_q ;
wire Xd_0__inst_mult_30_13_q ;
wire Xd_0__inst_mult_31_12_q ;
wire Xd_0__inst_mult_31_13_q ;
wire Xd_0__inst_mult_30_14_q ;
wire Xd_0__inst_mult_30_15_q ;
wire Xd_0__inst_mult_31_14_q ;
wire Xd_0__inst_mult_31_15_q ;
wire Xd_0__inst_mult_30_16_q ;
wire Xd_0__inst_mult_30_17_q ;
wire Xd_0__inst_mult_30_18_q ;
wire Xd_0__inst_mult_31_16_q ;
wire Xd_0__inst_mult_31_17_q ;
wire Xd_0__inst_mult_31_18_q ;
wire Xd_0__inst_mult_30_19_q ;
wire Xd_0__inst_mult_30_20_q ;
wire Xd_0__inst_mult_31_19_q ;
wire Xd_0__inst_mult_31_20_q ;
wire Xd_0__inst_mult_28_2_q ;
wire Xd_0__inst_mult_28_3_q ;
wire Xd_0__inst_mult_28_4_q ;
wire Xd_0__inst_mult_29_2_q ;
wire Xd_0__inst_mult_29_3_q ;
wire Xd_0__inst_mult_29_4_q ;
wire Xd_0__inst_mult_26_2_q ;
wire Xd_0__inst_mult_26_3_q ;
wire Xd_0__inst_mult_26_4_q ;
wire Xd_0__inst_mult_27_2_q ;
wire Xd_0__inst_mult_27_3_q ;
wire Xd_0__inst_mult_27_4_q ;
wire Xd_0__inst_mult_24_2_q ;
wire Xd_0__inst_mult_24_3_q ;
wire Xd_0__inst_mult_24_4_q ;
wire Xd_0__inst_mult_25_2_q ;
wire Xd_0__inst_mult_25_3_q ;
wire Xd_0__inst_mult_25_4_q ;
wire Xd_0__inst_mult_22_2_q ;
wire Xd_0__inst_mult_22_3_q ;
wire Xd_0__inst_mult_22_4_q ;
wire Xd_0__inst_mult_23_2_q ;
wire Xd_0__inst_mult_23_3_q ;
wire Xd_0__inst_mult_23_4_q ;
wire Xd_0__inst_mult_20_2_q ;
wire Xd_0__inst_mult_20_3_q ;
wire Xd_0__inst_mult_20_4_q ;
wire Xd_0__inst_mult_21_2_q ;
wire Xd_0__inst_mult_21_3_q ;
wire Xd_0__inst_mult_21_4_q ;
wire Xd_0__inst_mult_18_2_q ;
wire Xd_0__inst_mult_18_3_q ;
wire Xd_0__inst_mult_18_4_q ;
wire Xd_0__inst_mult_19_2_q ;
wire Xd_0__inst_mult_19_3_q ;
wire Xd_0__inst_mult_19_4_q ;
wire Xd_0__inst_mult_30_0_q ;
wire Xd_0__inst_mult_31_0_q ;
wire Xd_0__inst_mult_16_2_q ;
wire Xd_0__inst_mult_16_3_q ;
wire Xd_0__inst_mult_16_4_q ;
wire Xd_0__inst_mult_17_2_q ;
wire Xd_0__inst_mult_17_3_q ;
wire Xd_0__inst_mult_17_4_q ;
wire Xd_0__inst_mult_14_2_q ;
wire Xd_0__inst_mult_14_3_q ;
wire Xd_0__inst_mult_14_4_q ;
wire Xd_0__inst_mult_15_2_q ;
wire Xd_0__inst_mult_15_3_q ;
wire Xd_0__inst_mult_15_4_q ;
wire Xd_0__inst_mult_12_2_q ;
wire Xd_0__inst_mult_12_3_q ;
wire Xd_0__inst_mult_12_4_q ;
wire Xd_0__inst_mult_13_2_q ;
wire Xd_0__inst_mult_13_3_q ;
wire Xd_0__inst_mult_13_4_q ;
wire Xd_0__inst_mult_10_2_q ;
wire Xd_0__inst_mult_10_3_q ;
wire Xd_0__inst_mult_10_4_q ;
wire Xd_0__inst_mult_11_2_q ;
wire Xd_0__inst_mult_11_3_q ;
wire Xd_0__inst_mult_11_4_q ;
wire Xd_0__inst_mult_8_2_q ;
wire Xd_0__inst_mult_8_3_q ;
wire Xd_0__inst_mult_8_4_q ;
wire Xd_0__inst_mult_9_2_q ;
wire Xd_0__inst_mult_9_3_q ;
wire Xd_0__inst_mult_9_4_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_28_5_q ;
wire Xd_0__inst_mult_28_6_q ;
wire Xd_0__inst_mult_28_7_q ;
wire Xd_0__inst_mult_29_5_q ;
wire Xd_0__inst_mult_29_6_q ;
wire Xd_0__inst_mult_29_7_q ;
wire Xd_0__inst_mult_26_5_q ;
wire Xd_0__inst_mult_26_6_q ;
wire Xd_0__inst_mult_26_7_q ;
wire Xd_0__inst_mult_27_5_q ;
wire Xd_0__inst_mult_27_6_q ;
wire Xd_0__inst_mult_27_7_q ;
wire Xd_0__inst_mult_24_5_q ;
wire Xd_0__inst_mult_24_6_q ;
wire Xd_0__inst_mult_24_7_q ;
wire Xd_0__inst_mult_25_5_q ;
wire Xd_0__inst_mult_25_6_q ;
wire Xd_0__inst_mult_25_7_q ;
wire Xd_0__inst_mult_22_5_q ;
wire Xd_0__inst_mult_22_6_q ;
wire Xd_0__inst_mult_22_7_q ;
wire Xd_0__inst_mult_23_5_q ;
wire Xd_0__inst_mult_23_6_q ;
wire Xd_0__inst_mult_23_7_q ;
wire Xd_0__inst_mult_20_5_q ;
wire Xd_0__inst_mult_20_6_q ;
wire Xd_0__inst_mult_20_7_q ;
wire Xd_0__inst_mult_21_5_q ;
wire Xd_0__inst_mult_21_6_q ;
wire Xd_0__inst_mult_21_7_q ;
wire Xd_0__inst_mult_18_5_q ;
wire Xd_0__inst_mult_18_6_q ;
wire Xd_0__inst_mult_18_7_q ;
wire Xd_0__inst_mult_19_5_q ;
wire Xd_0__inst_mult_19_6_q ;
wire Xd_0__inst_mult_19_7_q ;
wire Xd_0__inst_mult_16_5_q ;
wire Xd_0__inst_mult_16_6_q ;
wire Xd_0__inst_mult_16_7_q ;
wire Xd_0__inst_mult_17_5_q ;
wire Xd_0__inst_mult_17_6_q ;
wire Xd_0__inst_mult_17_7_q ;
wire Xd_0__inst_mult_14_5_q ;
wire Xd_0__inst_mult_14_6_q ;
wire Xd_0__inst_mult_14_7_q ;
wire Xd_0__inst_mult_15_5_q ;
wire Xd_0__inst_mult_15_6_q ;
wire Xd_0__inst_mult_15_7_q ;
wire Xd_0__inst_mult_12_5_q ;
wire Xd_0__inst_mult_12_6_q ;
wire Xd_0__inst_mult_12_7_q ;
wire Xd_0__inst_mult_13_5_q ;
wire Xd_0__inst_mult_13_6_q ;
wire Xd_0__inst_mult_13_7_q ;
wire Xd_0__inst_mult_10_5_q ;
wire Xd_0__inst_mult_10_6_q ;
wire Xd_0__inst_mult_10_7_q ;
wire Xd_0__inst_mult_11_5_q ;
wire Xd_0__inst_mult_11_6_q ;
wire Xd_0__inst_mult_11_7_q ;
wire Xd_0__inst_mult_8_5_q ;
wire Xd_0__inst_mult_8_6_q ;
wire Xd_0__inst_mult_8_7_q ;
wire Xd_0__inst_mult_9_5_q ;
wire Xd_0__inst_mult_9_6_q ;
wire Xd_0__inst_mult_9_7_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_28_8_q ;
wire Xd_0__inst_mult_28_9_q ;
wire Xd_0__inst_mult_29_8_q ;
wire Xd_0__inst_mult_29_9_q ;
wire Xd_0__inst_mult_26_8_q ;
wire Xd_0__inst_mult_26_9_q ;
wire Xd_0__inst_mult_27_8_q ;
wire Xd_0__inst_mult_27_9_q ;
wire Xd_0__inst_mult_24_8_q ;
wire Xd_0__inst_mult_24_9_q ;
wire Xd_0__inst_mult_25_8_q ;
wire Xd_0__inst_mult_25_9_q ;
wire Xd_0__inst_mult_22_8_q ;
wire Xd_0__inst_mult_22_9_q ;
wire Xd_0__inst_mult_23_8_q ;
wire Xd_0__inst_mult_23_9_q ;
wire Xd_0__inst_mult_20_8_q ;
wire Xd_0__inst_mult_20_9_q ;
wire Xd_0__inst_mult_21_8_q ;
wire Xd_0__inst_mult_21_9_q ;
wire Xd_0__inst_mult_18_8_q ;
wire Xd_0__inst_mult_18_9_q ;
wire Xd_0__inst_mult_19_8_q ;
wire Xd_0__inst_mult_19_9_q ;
wire Xd_0__inst_mult_16_8_q ;
wire Xd_0__inst_mult_16_9_q ;
wire Xd_0__inst_mult_17_8_q ;
wire Xd_0__inst_mult_17_9_q ;
wire Xd_0__inst_mult_14_8_q ;
wire Xd_0__inst_mult_14_9_q ;
wire Xd_0__inst_mult_15_8_q ;
wire Xd_0__inst_mult_15_9_q ;
wire Xd_0__inst_mult_12_8_q ;
wire Xd_0__inst_mult_12_9_q ;
wire Xd_0__inst_mult_13_8_q ;
wire Xd_0__inst_mult_13_9_q ;
wire Xd_0__inst_mult_10_8_q ;
wire Xd_0__inst_mult_10_9_q ;
wire Xd_0__inst_mult_11_8_q ;
wire Xd_0__inst_mult_11_9_q ;
wire Xd_0__inst_mult_8_8_q ;
wire Xd_0__inst_mult_8_9_q ;
wire Xd_0__inst_mult_9_8_q ;
wire Xd_0__inst_mult_9_9_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_28_10_q ;
wire Xd_0__inst_mult_28_11_q ;
wire Xd_0__inst_mult_28_1_q ;
wire Xd_0__inst_mult_29_10_q ;
wire Xd_0__inst_mult_29_11_q ;
wire Xd_0__inst_mult_29_1_q ;
wire Xd_0__inst_mult_26_10_q ;
wire Xd_0__inst_mult_26_11_q ;
wire Xd_0__inst_mult_26_1_q ;
wire Xd_0__inst_mult_27_10_q ;
wire Xd_0__inst_mult_27_11_q ;
wire Xd_0__inst_mult_27_1_q ;
wire Xd_0__inst_mult_24_10_q ;
wire Xd_0__inst_mult_24_11_q ;
wire Xd_0__inst_mult_24_1_q ;
wire Xd_0__inst_mult_25_10_q ;
wire Xd_0__inst_mult_25_11_q ;
wire Xd_0__inst_mult_25_1_q ;
wire Xd_0__inst_mult_22_10_q ;
wire Xd_0__inst_mult_22_11_q ;
wire Xd_0__inst_mult_22_1_q ;
wire Xd_0__inst_mult_23_10_q ;
wire Xd_0__inst_mult_23_11_q ;
wire Xd_0__inst_mult_23_1_q ;
wire Xd_0__inst_mult_20_10_q ;
wire Xd_0__inst_mult_20_11_q ;
wire Xd_0__inst_mult_20_1_q ;
wire Xd_0__inst_mult_21_10_q ;
wire Xd_0__inst_mult_21_11_q ;
wire Xd_0__inst_mult_21_1_q ;
wire Xd_0__inst_mult_18_10_q ;
wire Xd_0__inst_mult_18_11_q ;
wire Xd_0__inst_mult_18_1_q ;
wire Xd_0__inst_mult_19_10_q ;
wire Xd_0__inst_mult_19_11_q ;
wire Xd_0__inst_mult_19_1_q ;
wire Xd_0__inst_mult_16_10_q ;
wire Xd_0__inst_mult_16_11_q ;
wire Xd_0__inst_mult_16_1_q ;
wire Xd_0__inst_mult_17_10_q ;
wire Xd_0__inst_mult_17_11_q ;
wire Xd_0__inst_mult_17_1_q ;
wire Xd_0__inst_mult_14_10_q ;
wire Xd_0__inst_mult_14_11_q ;
wire Xd_0__inst_mult_14_1_q ;
wire Xd_0__inst_mult_15_10_q ;
wire Xd_0__inst_mult_15_11_q ;
wire Xd_0__inst_mult_15_1_q ;
wire Xd_0__inst_mult_12_10_q ;
wire Xd_0__inst_mult_12_11_q ;
wire Xd_0__inst_mult_12_1_q ;
wire Xd_0__inst_mult_13_10_q ;
wire Xd_0__inst_mult_13_11_q ;
wire Xd_0__inst_mult_13_1_q ;
wire Xd_0__inst_mult_10_10_q ;
wire Xd_0__inst_mult_10_11_q ;
wire Xd_0__inst_mult_10_1_q ;
wire Xd_0__inst_mult_11_10_q ;
wire Xd_0__inst_mult_11_11_q ;
wire Xd_0__inst_mult_11_1_q ;
wire Xd_0__inst_mult_8_10_q ;
wire Xd_0__inst_mult_8_11_q ;
wire Xd_0__inst_mult_8_1_q ;
wire Xd_0__inst_mult_9_10_q ;
wire Xd_0__inst_mult_9_11_q ;
wire Xd_0__inst_mult_9_1_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_28_12_q ;
wire Xd_0__inst_mult_28_13_q ;
wire Xd_0__inst_mult_29_12_q ;
wire Xd_0__inst_mult_29_13_q ;
wire Xd_0__inst_mult_26_12_q ;
wire Xd_0__inst_mult_26_13_q ;
wire Xd_0__inst_mult_27_12_q ;
wire Xd_0__inst_mult_27_13_q ;
wire Xd_0__inst_mult_24_12_q ;
wire Xd_0__inst_mult_24_13_q ;
wire Xd_0__inst_mult_25_12_q ;
wire Xd_0__inst_mult_25_13_q ;
wire Xd_0__inst_mult_22_12_q ;
wire Xd_0__inst_mult_22_13_q ;
wire Xd_0__inst_mult_23_12_q ;
wire Xd_0__inst_mult_23_13_q ;
wire Xd_0__inst_mult_20_12_q ;
wire Xd_0__inst_mult_20_13_q ;
wire Xd_0__inst_mult_21_12_q ;
wire Xd_0__inst_mult_21_13_q ;
wire Xd_0__inst_mult_18_12_q ;
wire Xd_0__inst_mult_18_13_q ;
wire Xd_0__inst_mult_19_12_q ;
wire Xd_0__inst_mult_19_13_q ;
wire Xd_0__inst_mult_16_12_q ;
wire Xd_0__inst_mult_16_13_q ;
wire Xd_0__inst_mult_17_12_q ;
wire Xd_0__inst_mult_17_13_q ;
wire Xd_0__inst_mult_14_12_q ;
wire Xd_0__inst_mult_14_13_q ;
wire Xd_0__inst_mult_15_12_q ;
wire Xd_0__inst_mult_15_13_q ;
wire Xd_0__inst_mult_12_12_q ;
wire Xd_0__inst_mult_12_13_q ;
wire Xd_0__inst_mult_13_12_q ;
wire Xd_0__inst_mult_13_13_q ;
wire Xd_0__inst_mult_10_12_q ;
wire Xd_0__inst_mult_10_13_q ;
wire Xd_0__inst_mult_11_12_q ;
wire Xd_0__inst_mult_11_13_q ;
wire Xd_0__inst_mult_8_12_q ;
wire Xd_0__inst_mult_8_13_q ;
wire Xd_0__inst_mult_9_12_q ;
wire Xd_0__inst_mult_9_13_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_28_14_q ;
wire Xd_0__inst_mult_28_15_q ;
wire Xd_0__inst_mult_29_14_q ;
wire Xd_0__inst_mult_29_15_q ;
wire Xd_0__inst_mult_26_14_q ;
wire Xd_0__inst_mult_26_15_q ;
wire Xd_0__inst_mult_27_14_q ;
wire Xd_0__inst_mult_27_15_q ;
wire Xd_0__inst_mult_24_14_q ;
wire Xd_0__inst_mult_24_15_q ;
wire Xd_0__inst_mult_25_14_q ;
wire Xd_0__inst_mult_25_15_q ;
wire Xd_0__inst_mult_22_14_q ;
wire Xd_0__inst_mult_22_15_q ;
wire Xd_0__inst_mult_23_14_q ;
wire Xd_0__inst_mult_23_15_q ;
wire Xd_0__inst_mult_20_14_q ;
wire Xd_0__inst_mult_20_15_q ;
wire Xd_0__inst_mult_21_14_q ;
wire Xd_0__inst_mult_21_15_q ;
wire Xd_0__inst_mult_18_14_q ;
wire Xd_0__inst_mult_18_15_q ;
wire Xd_0__inst_mult_19_14_q ;
wire Xd_0__inst_mult_19_15_q ;
wire Xd_0__inst_mult_16_14_q ;
wire Xd_0__inst_mult_16_15_q ;
wire Xd_0__inst_mult_17_14_q ;
wire Xd_0__inst_mult_17_15_q ;
wire Xd_0__inst_mult_14_14_q ;
wire Xd_0__inst_mult_14_15_q ;
wire Xd_0__inst_mult_15_14_q ;
wire Xd_0__inst_mult_15_15_q ;
wire Xd_0__inst_mult_12_14_q ;
wire Xd_0__inst_mult_12_15_q ;
wire Xd_0__inst_mult_13_14_q ;
wire Xd_0__inst_mult_13_15_q ;
wire Xd_0__inst_mult_10_14_q ;
wire Xd_0__inst_mult_10_15_q ;
wire Xd_0__inst_mult_11_14_q ;
wire Xd_0__inst_mult_11_15_q ;
wire Xd_0__inst_mult_8_14_q ;
wire Xd_0__inst_mult_8_15_q ;
wire Xd_0__inst_mult_9_14_q ;
wire Xd_0__inst_mult_9_15_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_28_16_q ;
wire Xd_0__inst_mult_28_17_q ;
wire Xd_0__inst_mult_28_18_q ;
wire Xd_0__inst_mult_29_16_q ;
wire Xd_0__inst_mult_29_17_q ;
wire Xd_0__inst_mult_29_18_q ;
wire Xd_0__inst_mult_26_16_q ;
wire Xd_0__inst_mult_26_17_q ;
wire Xd_0__inst_mult_26_18_q ;
wire Xd_0__inst_mult_27_16_q ;
wire Xd_0__inst_mult_27_17_q ;
wire Xd_0__inst_mult_27_18_q ;
wire Xd_0__inst_mult_24_16_q ;
wire Xd_0__inst_mult_24_17_q ;
wire Xd_0__inst_mult_24_18_q ;
wire Xd_0__inst_mult_25_16_q ;
wire Xd_0__inst_mult_25_17_q ;
wire Xd_0__inst_mult_25_18_q ;
wire Xd_0__inst_mult_22_16_q ;
wire Xd_0__inst_mult_22_17_q ;
wire Xd_0__inst_mult_22_18_q ;
wire Xd_0__inst_mult_23_16_q ;
wire Xd_0__inst_mult_23_17_q ;
wire Xd_0__inst_mult_23_18_q ;
wire Xd_0__inst_mult_20_16_q ;
wire Xd_0__inst_mult_20_17_q ;
wire Xd_0__inst_mult_20_18_q ;
wire Xd_0__inst_mult_21_16_q ;
wire Xd_0__inst_mult_21_17_q ;
wire Xd_0__inst_mult_21_18_q ;
wire Xd_0__inst_mult_18_16_q ;
wire Xd_0__inst_mult_18_17_q ;
wire Xd_0__inst_mult_18_18_q ;
wire Xd_0__inst_mult_19_16_q ;
wire Xd_0__inst_mult_19_17_q ;
wire Xd_0__inst_mult_19_18_q ;
wire Xd_0__inst_mult_16_16_q ;
wire Xd_0__inst_mult_16_17_q ;
wire Xd_0__inst_mult_16_18_q ;
wire Xd_0__inst_mult_17_16_q ;
wire Xd_0__inst_mult_17_17_q ;
wire Xd_0__inst_mult_17_18_q ;
wire Xd_0__inst_mult_14_16_q ;
wire Xd_0__inst_mult_14_17_q ;
wire Xd_0__inst_mult_14_18_q ;
wire Xd_0__inst_mult_15_16_q ;
wire Xd_0__inst_mult_15_17_q ;
wire Xd_0__inst_mult_15_18_q ;
wire Xd_0__inst_mult_12_16_q ;
wire Xd_0__inst_mult_12_17_q ;
wire Xd_0__inst_mult_12_18_q ;
wire Xd_0__inst_mult_13_16_q ;
wire Xd_0__inst_mult_13_17_q ;
wire Xd_0__inst_mult_13_18_q ;
wire Xd_0__inst_mult_10_16_q ;
wire Xd_0__inst_mult_10_17_q ;
wire Xd_0__inst_mult_10_18_q ;
wire Xd_0__inst_mult_11_16_q ;
wire Xd_0__inst_mult_11_17_q ;
wire Xd_0__inst_mult_11_18_q ;
wire Xd_0__inst_mult_8_16_q ;
wire Xd_0__inst_mult_8_17_q ;
wire Xd_0__inst_mult_8_18_q ;
wire Xd_0__inst_mult_9_16_q ;
wire Xd_0__inst_mult_9_17_q ;
wire Xd_0__inst_mult_9_18_q ;
wire Xd_0__inst_mult_6_16_q ;
wire Xd_0__inst_mult_6_17_q ;
wire Xd_0__inst_mult_6_18_q ;
wire Xd_0__inst_mult_7_16_q ;
wire Xd_0__inst_mult_7_17_q ;
wire Xd_0__inst_mult_7_18_q ;
wire Xd_0__inst_mult_4_16_q ;
wire Xd_0__inst_mult_4_17_q ;
wire Xd_0__inst_mult_4_18_q ;
wire Xd_0__inst_mult_5_16_q ;
wire Xd_0__inst_mult_5_17_q ;
wire Xd_0__inst_mult_5_18_q ;
wire Xd_0__inst_mult_2_16_q ;
wire Xd_0__inst_mult_2_17_q ;
wire Xd_0__inst_mult_2_18_q ;
wire Xd_0__inst_mult_3_16_q ;
wire Xd_0__inst_mult_3_17_q ;
wire Xd_0__inst_mult_3_18_q ;
wire Xd_0__inst_mult_0_16_q ;
wire Xd_0__inst_mult_0_17_q ;
wire Xd_0__inst_mult_0_18_q ;
wire Xd_0__inst_mult_1_16_q ;
wire Xd_0__inst_mult_1_17_q ;
wire Xd_0__inst_mult_1_18_q ;
wire Xd_0__inst_mult_28_19_q ;
wire Xd_0__inst_mult_28_20_q ;
wire Xd_0__inst_mult_29_19_q ;
wire Xd_0__inst_mult_29_20_q ;
wire Xd_0__inst_mult_26_19_q ;
wire Xd_0__inst_mult_26_20_q ;
wire Xd_0__inst_mult_27_19_q ;
wire Xd_0__inst_mult_27_20_q ;
wire Xd_0__inst_mult_24_19_q ;
wire Xd_0__inst_mult_24_20_q ;
wire Xd_0__inst_mult_25_19_q ;
wire Xd_0__inst_mult_25_20_q ;
wire Xd_0__inst_mult_22_19_q ;
wire Xd_0__inst_mult_22_20_q ;
wire Xd_0__inst_mult_23_19_q ;
wire Xd_0__inst_mult_23_20_q ;
wire Xd_0__inst_mult_20_19_q ;
wire Xd_0__inst_mult_20_20_q ;
wire Xd_0__inst_mult_21_19_q ;
wire Xd_0__inst_mult_21_20_q ;
wire Xd_0__inst_mult_18_19_q ;
wire Xd_0__inst_mult_18_20_q ;
wire Xd_0__inst_mult_19_19_q ;
wire Xd_0__inst_mult_19_20_q ;
wire Xd_0__inst_mult_16_19_q ;
wire Xd_0__inst_mult_16_20_q ;
wire Xd_0__inst_mult_17_19_q ;
wire Xd_0__inst_mult_17_20_q ;
wire Xd_0__inst_mult_14_19_q ;
wire Xd_0__inst_mult_14_20_q ;
wire Xd_0__inst_mult_15_19_q ;
wire Xd_0__inst_mult_15_20_q ;
wire Xd_0__inst_mult_12_19_q ;
wire Xd_0__inst_mult_12_20_q ;
wire Xd_0__inst_mult_13_19_q ;
wire Xd_0__inst_mult_13_20_q ;
wire Xd_0__inst_mult_10_19_q ;
wire Xd_0__inst_mult_10_20_q ;
wire Xd_0__inst_mult_11_19_q ;
wire Xd_0__inst_mult_11_20_q ;
wire Xd_0__inst_mult_8_19_q ;
wire Xd_0__inst_mult_8_20_q ;
wire Xd_0__inst_mult_9_19_q ;
wire Xd_0__inst_mult_9_20_q ;
wire Xd_0__inst_mult_6_19_q ;
wire Xd_0__inst_mult_6_20_q ;
wire Xd_0__inst_mult_7_19_q ;
wire Xd_0__inst_mult_7_20_q ;
wire Xd_0__inst_mult_4_19_q ;
wire Xd_0__inst_mult_4_20_q ;
wire Xd_0__inst_mult_5_19_q ;
wire Xd_0__inst_mult_5_20_q ;
wire Xd_0__inst_mult_2_19_q ;
wire Xd_0__inst_mult_2_20_q ;
wire Xd_0__inst_mult_3_19_q ;
wire Xd_0__inst_mult_3_20_q ;
wire Xd_0__inst_mult_0_19_q ;
wire Xd_0__inst_mult_0_20_q ;
wire Xd_0__inst_mult_1_19_q ;
wire Xd_0__inst_mult_1_20_q ;
wire Xd_0__inst_mult_28_0_q ;
wire Xd_0__inst_mult_29_0_q ;
wire Xd_0__inst_mult_26_0_q ;
wire Xd_0__inst_mult_27_0_q ;
wire Xd_0__inst_mult_24_0_q ;
wire Xd_0__inst_mult_25_0_q ;
wire Xd_0__inst_mult_22_0_q ;
wire Xd_0__inst_mult_23_0_q ;
wire Xd_0__inst_mult_20_0_q ;
wire Xd_0__inst_mult_21_0_q ;
wire Xd_0__inst_mult_18_0_q ;
wire Xd_0__inst_mult_19_0_q ;
wire Xd_0__inst_mult_16_0_q ;
wire Xd_0__inst_mult_17_0_q ;
wire Xd_0__inst_mult_14_0_q ;
wire Xd_0__inst_mult_15_0_q ;
wire Xd_0__inst_mult_12_0_q ;
wire Xd_0__inst_mult_13_0_q ;
wire Xd_0__inst_mult_10_0_q ;
wire Xd_0__inst_mult_11_0_q ;
wire Xd_0__inst_mult_8_0_q ;
wire Xd_0__inst_mult_9_0_q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_1_0_q ;
wire [17:0] Xd_0__inst_inst_inst_inst_dout ;
wire [13:0] Xd_0__inst_a1_0__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_1__adder1_inst_dout ;
wire [0:31] Xd_0__inst_sign1 ;
wire [13:0] Xd_0__inst_a1_2__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_3__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_4__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_5__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_12__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_13__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_14__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_15__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_11__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_10__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_9__adder1_inst_dout ;
wire [0:31] Xd_0__inst_sign ;
wire [13:0] Xd_0__inst_a1_8__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_7__adder1_inst_dout ;
wire [13:0] Xd_0__inst_a1_6__adder1_inst_dout ;


twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_1_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__0__q  ) + ( Xd_0__inst_inst_inst_first_level_0__0__q  ) + ( Xd_0__inst_i19_2  ))
// Xd_0__inst_inst_inst_inst_add_0_2  = CARRY(( Xd_0__inst_inst_inst_first_level_1__0__q  ) + ( Xd_0__inst_inst_inst_first_level_0__0__q  ) + ( Xd_0__inst_i19_2  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__0__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__0__q ),
	.datag(gnd),
	.cin(Xd_0__inst_i19_2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_5_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__1__q  ) + ( Xd_0__inst_inst_inst_first_level_0__1__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_inst_add_0_6  = CARRY(( Xd_0__inst_inst_inst_first_level_1__1__q  ) + ( Xd_0__inst_inst_inst_first_level_0__1__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_2  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__1__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__1__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_6 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_9_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__2__q  ) + ( Xd_0__inst_inst_inst_first_level_0__2__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_inst_add_0_10  = CARRY(( Xd_0__inst_inst_inst_first_level_1__2__q  ) + ( Xd_0__inst_inst_inst_first_level_0__2__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_6  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__2__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__2__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_10 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_13_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__3__q  ) + ( Xd_0__inst_inst_inst_first_level_0__3__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_inst_add_0_14  = CARRY(( Xd_0__inst_inst_inst_first_level_1__3__q  ) + ( Xd_0__inst_inst_inst_first_level_0__3__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_10  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__3__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__3__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_10 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_14 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_17_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__4__q  ) + ( Xd_0__inst_inst_inst_first_level_0__4__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_inst_add_0_18  = CARRY(( Xd_0__inst_inst_inst_first_level_1__4__q  ) + ( Xd_0__inst_inst_inst_first_level_0__4__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_14  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__4__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__4__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_14 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_18 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_21_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__5__q  ) + ( Xd_0__inst_inst_inst_first_level_0__5__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_inst_add_0_22  = CARRY(( Xd_0__inst_inst_inst_first_level_1__5__q  ) + ( Xd_0__inst_inst_inst_first_level_0__5__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_18  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__5__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__5__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_18 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_25_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__6__q  ) + ( Xd_0__inst_inst_inst_first_level_0__6__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_inst_add_0_26  = CARRY(( Xd_0__inst_inst_inst_first_level_1__6__q  ) + ( Xd_0__inst_inst_inst_first_level_0__6__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_22  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__6__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__6__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_26 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_29_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__7__q  ) + ( Xd_0__inst_inst_inst_first_level_0__7__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_inst_add_0_30  = CARRY(( Xd_0__inst_inst_inst_first_level_1__7__q  ) + ( Xd_0__inst_inst_inst_first_level_0__7__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_26  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__7__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__7__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_26 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_30 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_33_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__8__q  ) + ( Xd_0__inst_inst_inst_first_level_0__8__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_inst_add_0_34  = CARRY(( Xd_0__inst_inst_inst_first_level_1__8__q  ) + ( Xd_0__inst_inst_inst_first_level_0__8__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_30  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__8__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__8__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_30 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_34 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_37_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__9__q  ) + ( Xd_0__inst_inst_inst_first_level_0__9__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_inst_add_0_38  = CARRY(( Xd_0__inst_inst_inst_first_level_1__9__q  ) + ( Xd_0__inst_inst_inst_first_level_0__9__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_34  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__9__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__9__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_34 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_38 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_41_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__10__q  ) + ( Xd_0__inst_inst_inst_first_level_0__10__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_inst_add_0_42  = CARRY(( Xd_0__inst_inst_inst_first_level_1__10__q  ) + ( Xd_0__inst_inst_inst_first_level_0__10__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_38  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__10__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__10__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_38 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_45_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__11__q  ) + ( Xd_0__inst_inst_inst_first_level_0__11__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_inst_add_0_46  = CARRY(( Xd_0__inst_inst_inst_first_level_1__11__q  ) + ( Xd_0__inst_inst_inst_first_level_0__11__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_42  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__11__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__11__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_46 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_49_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__12__q  ) + ( Xd_0__inst_inst_inst_first_level_0__12__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_inst_add_0_50  = CARRY(( Xd_0__inst_inst_inst_first_level_1__12__q  ) + ( Xd_0__inst_inst_inst_first_level_0__12__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_46  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__12__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__12__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_46 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_50 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_53_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__13__q  ) + ( Xd_0__inst_inst_inst_first_level_0__13__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_inst_add_0_54  = CARRY(( Xd_0__inst_inst_inst_first_level_1__13__q  ) + ( Xd_0__inst_inst_inst_first_level_0__13__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_50  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__13__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__13__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_50 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_54 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_57_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__14__q  ) + ( Xd_0__inst_inst_inst_first_level_0__14__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_inst_add_0_58  = CARRY(( Xd_0__inst_inst_inst_first_level_1__14__q  ) + ( Xd_0__inst_inst_inst_first_level_0__14__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_54  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__14__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__14__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_54 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_58 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_61_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__15__q  ) + ( Xd_0__inst_inst_inst_first_level_0__15__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_58  ))
// Xd_0__inst_inst_inst_inst_add_0_62  = CARRY(( Xd_0__inst_inst_inst_first_level_1__15__q  ) + ( Xd_0__inst_inst_inst_first_level_0__15__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_58  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__15__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__15__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_58 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_65 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_65_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__16__q  ) + ( Xd_0__inst_inst_inst_first_level_0__16__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_62  ))
// Xd_0__inst_inst_inst_inst_add_0_66  = CARRY(( Xd_0__inst_inst_inst_first_level_1__16__q  ) + ( Xd_0__inst_inst_inst_first_level_0__16__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_62  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__16__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__16__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_62 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_65_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_66 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FF00000000FF),
	.shared_arith("off")
) Xd_0__inst_inst_inst_inst_add_0_69 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_69_sumout  = SUM(( Xd_0__inst_inst_inst_first_level_1__17__q  ) + ( Xd_0__inst_inst_inst_first_level_0__17__q  ) + ( Xd_0__inst_inst_inst_inst_add_0_66  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__17__q ),
	.datae(gnd),
	.dataf(!Xd_0__inst_inst_inst_first_level_0__17__q ),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_66 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_69_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00006666),
	.shared_arith("off")
) Xd_0__inst_i19_1 (
// Equation(s):
// Xd_0__inst_i19_1_sumout  = SUM(( !din_a[202] $ (!din_b[202]) ) + ( GND ) + ( Xd_0__inst_i19_6  ))
// Xd_0__inst_i19_2  = CARRY(( !din_a[202] $ (!din_b[202]) ) + ( GND ) + ( Xd_0__inst_i19_6  ))

	.dataa(!din_a[202]),
	.datab(!din_b[202]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_6 ),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_1_sumout ),
	.cout(Xd_0__inst_i19_2 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_1 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__0__q  $ (!Xd_0__inst_inst_first_level_3__0__q  $ (Xd_0__inst_inst_first_level_5__0__q )) ) + ( Xd_0__inst_i19_11  ) + ( Xd_0__inst_i19_10  ))
// Xd_0__inst_inst_inst_add_3_2  = CARRY(( !Xd_0__inst_inst_first_level_4__0__q  $ (!Xd_0__inst_inst_first_level_3__0__q  $ (Xd_0__inst_inst_first_level_5__0__q )) ) + ( Xd_0__inst_i19_11  ) + ( Xd_0__inst_i19_10  ))
// Xd_0__inst_inst_inst_add_3_3  = SHARE((!Xd_0__inst_inst_first_level_4__0__q  & (Xd_0__inst_inst_first_level_3__0__q  & Xd_0__inst_inst_first_level_5__0__q )) # (Xd_0__inst_inst_first_level_4__0__q  & ((Xd_0__inst_inst_first_level_5__0__q ) # 
// (Xd_0__inst_inst_first_level_3__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__0__q ),
	.datac(!Xd_0__inst_inst_first_level_3__0__q ),
	.datad(!Xd_0__inst_inst_first_level_5__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_10 ),
	.sharein(Xd_0__inst_i19_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_2 ),
	.shareout(Xd_0__inst_inst_inst_add_3_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_i19_15  ) + ( Xd_0__inst_i19_14  ))
// Xd_0__inst_inst_inst_add_0_2  = CARRY(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_i19_15  ) + ( Xd_0__inst_i19_14  ))
// Xd_0__inst_inst_inst_add_0_3  = SHARE((!Xd_0__inst_inst_first_level_2__0__q  & (Xd_0__inst_inst_first_level_1__0__q  & Xd_0__inst_inst_first_level_0__0__q )) # (Xd_0__inst_inst_first_level_2__0__q  & ((Xd_0__inst_inst_first_level_0__0__q ) # 
// (Xd_0__inst_inst_first_level_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__0__q ),
	.datac(!Xd_0__inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_14 ),
	.sharein(Xd_0__inst_i19_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00006666),
	.shared_arith("off")
) Xd_0__inst_i19_5 (
// Equation(s):
// Xd_0__inst_i19_5_sumout  = SUM(( !din_a[209] $ (!din_b[209]) ) + ( GND ) + ( !VCC ))
// Xd_0__inst_i19_6  = CARRY(( !din_a[209] $ (!din_b[209]) ) + ( GND ) + ( !VCC ))

	.dataa(!din_a[209]),
	.datab(!din_b[209]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_5_sumout ),
	.cout(Xd_0__inst_i19_6 ),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_5 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__1__q  $ (!Xd_0__inst_inst_first_level_3__1__q  $ (Xd_0__inst_inst_first_level_5__1__q )) ) + ( Xd_0__inst_inst_inst_add_3_3  ) + ( Xd_0__inst_inst_inst_add_3_2  ))
// Xd_0__inst_inst_inst_add_3_6  = CARRY(( !Xd_0__inst_inst_first_level_4__1__q  $ (!Xd_0__inst_inst_first_level_3__1__q  $ (Xd_0__inst_inst_first_level_5__1__q )) ) + ( Xd_0__inst_inst_inst_add_3_3  ) + ( Xd_0__inst_inst_inst_add_3_2  ))
// Xd_0__inst_inst_inst_add_3_7  = SHARE((!Xd_0__inst_inst_first_level_4__1__q  & (Xd_0__inst_inst_first_level_3__1__q  & Xd_0__inst_inst_first_level_5__1__q )) # (Xd_0__inst_inst_first_level_4__1__q  & ((Xd_0__inst_inst_first_level_5__1__q ) # 
// (Xd_0__inst_inst_first_level_3__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__1__q ),
	.datac(!Xd_0__inst_inst_first_level_3__1__q ),
	.datad(!Xd_0__inst_inst_first_level_5__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_2 ),
	.sharein(Xd_0__inst_inst_inst_add_3_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_5_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_6 ),
	.shareout(Xd_0__inst_inst_inst_add_3_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_6  = CARRY(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_7  = SHARE((!Xd_0__inst_inst_first_level_2__1__q  & (Xd_0__inst_inst_first_level_1__1__q  & Xd_0__inst_inst_first_level_0__1__q )) # (Xd_0__inst_inst_first_level_2__1__q  & ((Xd_0__inst_inst_first_level_0__1__q ) # 
// (Xd_0__inst_inst_first_level_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__1__q ),
	.datac(!Xd_0__inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_9 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__2__q  $ (!Xd_0__inst_inst_first_level_3__2__q  $ (Xd_0__inst_inst_first_level_5__2__q )) ) + ( Xd_0__inst_inst_inst_add_3_7  ) + ( Xd_0__inst_inst_inst_add_3_6  ))
// Xd_0__inst_inst_inst_add_3_10  = CARRY(( !Xd_0__inst_inst_first_level_4__2__q  $ (!Xd_0__inst_inst_first_level_3__2__q  $ (Xd_0__inst_inst_first_level_5__2__q )) ) + ( Xd_0__inst_inst_inst_add_3_7  ) + ( Xd_0__inst_inst_inst_add_3_6  ))
// Xd_0__inst_inst_inst_add_3_11  = SHARE((!Xd_0__inst_inst_first_level_4__2__q  & (Xd_0__inst_inst_first_level_3__2__q  & Xd_0__inst_inst_first_level_5__2__q )) # (Xd_0__inst_inst_first_level_4__2__q  & ((Xd_0__inst_inst_first_level_5__2__q ) # 
// (Xd_0__inst_inst_first_level_3__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__2__q ),
	.datac(!Xd_0__inst_inst_first_level_3__2__q ),
	.datad(!Xd_0__inst_inst_first_level_5__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_6 ),
	.sharein(Xd_0__inst_inst_inst_add_3_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_9_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_10 ),
	.shareout(Xd_0__inst_inst_inst_add_3_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_10  = CARRY(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_11  = SHARE((!Xd_0__inst_inst_first_level_2__2__q  & (Xd_0__inst_inst_first_level_1__2__q  & Xd_0__inst_inst_first_level_0__2__q )) # (Xd_0__inst_inst_first_level_2__2__q  & ((Xd_0__inst_inst_first_level_0__2__q ) # 
// (Xd_0__inst_inst_first_level_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__2__q ),
	.datac(!Xd_0__inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_13 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__3__q  $ (!Xd_0__inst_inst_first_level_3__3__q  $ (Xd_0__inst_inst_first_level_5__3__q )) ) + ( Xd_0__inst_inst_inst_add_3_11  ) + ( Xd_0__inst_inst_inst_add_3_10  ))
// Xd_0__inst_inst_inst_add_3_14  = CARRY(( !Xd_0__inst_inst_first_level_4__3__q  $ (!Xd_0__inst_inst_first_level_3__3__q  $ (Xd_0__inst_inst_first_level_5__3__q )) ) + ( Xd_0__inst_inst_inst_add_3_11  ) + ( Xd_0__inst_inst_inst_add_3_10  ))
// Xd_0__inst_inst_inst_add_3_15  = SHARE((!Xd_0__inst_inst_first_level_4__3__q  & (Xd_0__inst_inst_first_level_3__3__q  & Xd_0__inst_inst_first_level_5__3__q )) # (Xd_0__inst_inst_first_level_4__3__q  & ((Xd_0__inst_inst_first_level_5__3__q ) # 
// (Xd_0__inst_inst_first_level_3__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__3__q ),
	.datac(!Xd_0__inst_inst_first_level_3__3__q ),
	.datad(!Xd_0__inst_inst_first_level_5__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_10 ),
	.sharein(Xd_0__inst_inst_inst_add_3_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_13_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_14 ),
	.shareout(Xd_0__inst_inst_inst_add_3_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_14  = CARRY(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_15  = SHARE((!Xd_0__inst_inst_first_level_2__3__q  & (Xd_0__inst_inst_first_level_1__3__q  & Xd_0__inst_inst_first_level_0__3__q )) # (Xd_0__inst_inst_first_level_2__3__q  & ((Xd_0__inst_inst_first_level_0__3__q ) # 
// (Xd_0__inst_inst_first_level_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__3__q ),
	.datac(!Xd_0__inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_17 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__4__q  $ (!Xd_0__inst_inst_first_level_3__4__q  $ (Xd_0__inst_inst_first_level_5__4__q )) ) + ( Xd_0__inst_inst_inst_add_3_15  ) + ( Xd_0__inst_inst_inst_add_3_14  ))
// Xd_0__inst_inst_inst_add_3_18  = CARRY(( !Xd_0__inst_inst_first_level_4__4__q  $ (!Xd_0__inst_inst_first_level_3__4__q  $ (Xd_0__inst_inst_first_level_5__4__q )) ) + ( Xd_0__inst_inst_inst_add_3_15  ) + ( Xd_0__inst_inst_inst_add_3_14  ))
// Xd_0__inst_inst_inst_add_3_19  = SHARE((!Xd_0__inst_inst_first_level_4__4__q  & (Xd_0__inst_inst_first_level_3__4__q  & Xd_0__inst_inst_first_level_5__4__q )) # (Xd_0__inst_inst_first_level_4__4__q  & ((Xd_0__inst_inst_first_level_5__4__q ) # 
// (Xd_0__inst_inst_first_level_3__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__4__q ),
	.datac(!Xd_0__inst_inst_first_level_3__4__q ),
	.datad(!Xd_0__inst_inst_first_level_5__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_14 ),
	.sharein(Xd_0__inst_inst_inst_add_3_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_17_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_18 ),
	.shareout(Xd_0__inst_inst_inst_add_3_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_18  = CARRY(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_19  = SHARE((!Xd_0__inst_inst_first_level_2__4__q  & (Xd_0__inst_inst_first_level_1__4__q  & Xd_0__inst_inst_first_level_0__4__q )) # (Xd_0__inst_inst_first_level_2__4__q  & ((Xd_0__inst_inst_first_level_0__4__q ) # 
// (Xd_0__inst_inst_first_level_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__4__q ),
	.datac(!Xd_0__inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_21 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__5__q  $ (!Xd_0__inst_inst_first_level_3__5__q  $ (Xd_0__inst_inst_first_level_5__5__q )) ) + ( Xd_0__inst_inst_inst_add_3_19  ) + ( Xd_0__inst_inst_inst_add_3_18  ))
// Xd_0__inst_inst_inst_add_3_22  = CARRY(( !Xd_0__inst_inst_first_level_4__5__q  $ (!Xd_0__inst_inst_first_level_3__5__q  $ (Xd_0__inst_inst_first_level_5__5__q )) ) + ( Xd_0__inst_inst_inst_add_3_19  ) + ( Xd_0__inst_inst_inst_add_3_18  ))
// Xd_0__inst_inst_inst_add_3_23  = SHARE((!Xd_0__inst_inst_first_level_4__5__q  & (Xd_0__inst_inst_first_level_3__5__q  & Xd_0__inst_inst_first_level_5__5__q )) # (Xd_0__inst_inst_first_level_4__5__q  & ((Xd_0__inst_inst_first_level_5__5__q ) # 
// (Xd_0__inst_inst_first_level_3__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__5__q ),
	.datac(!Xd_0__inst_inst_first_level_3__5__q ),
	.datad(!Xd_0__inst_inst_first_level_5__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_18 ),
	.sharein(Xd_0__inst_inst_inst_add_3_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_22 ),
	.shareout(Xd_0__inst_inst_inst_add_3_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_22  = CARRY(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_23  = SHARE((!Xd_0__inst_inst_first_level_2__5__q  & (Xd_0__inst_inst_first_level_1__5__q  & Xd_0__inst_inst_first_level_0__5__q )) # (Xd_0__inst_inst_first_level_2__5__q  & ((Xd_0__inst_inst_first_level_0__5__q ) # 
// (Xd_0__inst_inst_first_level_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__5__q ),
	.datac(!Xd_0__inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_25 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__6__q  $ (!Xd_0__inst_inst_first_level_3__6__q  $ (Xd_0__inst_inst_first_level_5__6__q )) ) + ( Xd_0__inst_inst_inst_add_3_23  ) + ( Xd_0__inst_inst_inst_add_3_22  ))
// Xd_0__inst_inst_inst_add_3_26  = CARRY(( !Xd_0__inst_inst_first_level_4__6__q  $ (!Xd_0__inst_inst_first_level_3__6__q  $ (Xd_0__inst_inst_first_level_5__6__q )) ) + ( Xd_0__inst_inst_inst_add_3_23  ) + ( Xd_0__inst_inst_inst_add_3_22  ))
// Xd_0__inst_inst_inst_add_3_27  = SHARE((!Xd_0__inst_inst_first_level_4__6__q  & (Xd_0__inst_inst_first_level_3__6__q  & Xd_0__inst_inst_first_level_5__6__q )) # (Xd_0__inst_inst_first_level_4__6__q  & ((Xd_0__inst_inst_first_level_5__6__q ) # 
// (Xd_0__inst_inst_first_level_3__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__6__q ),
	.datac(!Xd_0__inst_inst_first_level_3__6__q ),
	.datad(!Xd_0__inst_inst_first_level_5__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_22 ),
	.sharein(Xd_0__inst_inst_inst_add_3_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_25_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_26 ),
	.shareout(Xd_0__inst_inst_inst_add_3_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_26  = CARRY(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_27  = SHARE((!Xd_0__inst_inst_first_level_2__6__q  & (Xd_0__inst_inst_first_level_1__6__q  & Xd_0__inst_inst_first_level_0__6__q )) # (Xd_0__inst_inst_first_level_2__6__q  & ((Xd_0__inst_inst_first_level_0__6__q ) # 
// (Xd_0__inst_inst_first_level_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__6__q ),
	.datac(!Xd_0__inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_29 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__7__q  $ (!Xd_0__inst_inst_first_level_3__7__q  $ (Xd_0__inst_inst_first_level_5__7__q )) ) + ( Xd_0__inst_inst_inst_add_3_27  ) + ( Xd_0__inst_inst_inst_add_3_26  ))
// Xd_0__inst_inst_inst_add_3_30  = CARRY(( !Xd_0__inst_inst_first_level_4__7__q  $ (!Xd_0__inst_inst_first_level_3__7__q  $ (Xd_0__inst_inst_first_level_5__7__q )) ) + ( Xd_0__inst_inst_inst_add_3_27  ) + ( Xd_0__inst_inst_inst_add_3_26  ))
// Xd_0__inst_inst_inst_add_3_31  = SHARE((!Xd_0__inst_inst_first_level_4__7__q  & (Xd_0__inst_inst_first_level_3__7__q  & Xd_0__inst_inst_first_level_5__7__q )) # (Xd_0__inst_inst_first_level_4__7__q  & ((Xd_0__inst_inst_first_level_5__7__q ) # 
// (Xd_0__inst_inst_first_level_3__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__7__q ),
	.datac(!Xd_0__inst_inst_first_level_3__7__q ),
	.datad(!Xd_0__inst_inst_first_level_5__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_26 ),
	.sharein(Xd_0__inst_inst_inst_add_3_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_29_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_30 ),
	.shareout(Xd_0__inst_inst_inst_add_3_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_30  = CARRY(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_31  = SHARE((!Xd_0__inst_inst_first_level_2__7__q  & (Xd_0__inst_inst_first_level_1__7__q  & Xd_0__inst_inst_first_level_0__7__q )) # (Xd_0__inst_inst_first_level_2__7__q  & ((Xd_0__inst_inst_first_level_0__7__q ) # 
// (Xd_0__inst_inst_first_level_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__7__q ),
	.datac(!Xd_0__inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_33 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__8__q  $ (!Xd_0__inst_inst_first_level_3__8__q  $ (Xd_0__inst_inst_first_level_5__8__q )) ) + ( Xd_0__inst_inst_inst_add_3_31  ) + ( Xd_0__inst_inst_inst_add_3_30  ))
// Xd_0__inst_inst_inst_add_3_34  = CARRY(( !Xd_0__inst_inst_first_level_4__8__q  $ (!Xd_0__inst_inst_first_level_3__8__q  $ (Xd_0__inst_inst_first_level_5__8__q )) ) + ( Xd_0__inst_inst_inst_add_3_31  ) + ( Xd_0__inst_inst_inst_add_3_30  ))
// Xd_0__inst_inst_inst_add_3_35  = SHARE((!Xd_0__inst_inst_first_level_4__8__q  & (Xd_0__inst_inst_first_level_3__8__q  & Xd_0__inst_inst_first_level_5__8__q )) # (Xd_0__inst_inst_first_level_4__8__q  & ((Xd_0__inst_inst_first_level_5__8__q ) # 
// (Xd_0__inst_inst_first_level_3__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__8__q ),
	.datac(!Xd_0__inst_inst_first_level_3__8__q ),
	.datad(!Xd_0__inst_inst_first_level_5__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_30 ),
	.sharein(Xd_0__inst_inst_inst_add_3_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_33_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_34 ),
	.shareout(Xd_0__inst_inst_inst_add_3_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_34  = CARRY(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_35  = SHARE((!Xd_0__inst_inst_first_level_2__8__q  & (Xd_0__inst_inst_first_level_1__8__q  & Xd_0__inst_inst_first_level_0__8__q )) # (Xd_0__inst_inst_first_level_2__8__q  & ((Xd_0__inst_inst_first_level_0__8__q ) # 
// (Xd_0__inst_inst_first_level_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__8__q ),
	.datac(!Xd_0__inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_37 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__9__q  $ (!Xd_0__inst_inst_first_level_3__9__q  $ (Xd_0__inst_inst_first_level_5__9__q )) ) + ( Xd_0__inst_inst_inst_add_3_35  ) + ( Xd_0__inst_inst_inst_add_3_34  ))
// Xd_0__inst_inst_inst_add_3_38  = CARRY(( !Xd_0__inst_inst_first_level_4__9__q  $ (!Xd_0__inst_inst_first_level_3__9__q  $ (Xd_0__inst_inst_first_level_5__9__q )) ) + ( Xd_0__inst_inst_inst_add_3_35  ) + ( Xd_0__inst_inst_inst_add_3_34  ))
// Xd_0__inst_inst_inst_add_3_39  = SHARE((!Xd_0__inst_inst_first_level_4__9__q  & (Xd_0__inst_inst_first_level_3__9__q  & Xd_0__inst_inst_first_level_5__9__q )) # (Xd_0__inst_inst_first_level_4__9__q  & ((Xd_0__inst_inst_first_level_5__9__q ) # 
// (Xd_0__inst_inst_first_level_3__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__9__q ),
	.datac(!Xd_0__inst_inst_first_level_3__9__q ),
	.datad(!Xd_0__inst_inst_first_level_5__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_34 ),
	.sharein(Xd_0__inst_inst_inst_add_3_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_37_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_38 ),
	.shareout(Xd_0__inst_inst_inst_add_3_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_38  = CARRY(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_39  = SHARE((!Xd_0__inst_inst_first_level_2__9__q  & (Xd_0__inst_inst_first_level_1__9__q  & Xd_0__inst_inst_first_level_0__9__q )) # (Xd_0__inst_inst_first_level_2__9__q  & ((Xd_0__inst_inst_first_level_0__9__q ) # 
// (Xd_0__inst_inst_first_level_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__9__q ),
	.datac(!Xd_0__inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_41 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__10__q  $ (!Xd_0__inst_inst_first_level_3__10__q  $ (Xd_0__inst_inst_first_level_5__10__q )) ) + ( Xd_0__inst_inst_inst_add_3_39  ) + ( Xd_0__inst_inst_inst_add_3_38  ))
// Xd_0__inst_inst_inst_add_3_42  = CARRY(( !Xd_0__inst_inst_first_level_4__10__q  $ (!Xd_0__inst_inst_first_level_3__10__q  $ (Xd_0__inst_inst_first_level_5__10__q )) ) + ( Xd_0__inst_inst_inst_add_3_39  ) + ( Xd_0__inst_inst_inst_add_3_38  ))
// Xd_0__inst_inst_inst_add_3_43  = SHARE((!Xd_0__inst_inst_first_level_4__10__q  & (Xd_0__inst_inst_first_level_3__10__q  & Xd_0__inst_inst_first_level_5__10__q )) # (Xd_0__inst_inst_first_level_4__10__q  & ((Xd_0__inst_inst_first_level_5__10__q ) # 
// (Xd_0__inst_inst_first_level_3__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__10__q ),
	.datac(!Xd_0__inst_inst_first_level_3__10__q ),
	.datad(!Xd_0__inst_inst_first_level_5__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_38 ),
	.sharein(Xd_0__inst_inst_inst_add_3_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_42 ),
	.shareout(Xd_0__inst_inst_inst_add_3_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_42  = CARRY(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_43  = SHARE((!Xd_0__inst_inst_first_level_2__10__q  & (Xd_0__inst_inst_first_level_1__10__q  & Xd_0__inst_inst_first_level_0__10__q )) # (Xd_0__inst_inst_first_level_2__10__q  & ((Xd_0__inst_inst_first_level_0__10__q ) # 
// (Xd_0__inst_inst_first_level_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__10__q ),
	.datac(!Xd_0__inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_45 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__11__q  $ (!Xd_0__inst_inst_first_level_3__11__q  $ (Xd_0__inst_inst_first_level_5__11__q )) ) + ( Xd_0__inst_inst_inst_add_3_43  ) + ( Xd_0__inst_inst_inst_add_3_42  ))
// Xd_0__inst_inst_inst_add_3_46  = CARRY(( !Xd_0__inst_inst_first_level_4__11__q  $ (!Xd_0__inst_inst_first_level_3__11__q  $ (Xd_0__inst_inst_first_level_5__11__q )) ) + ( Xd_0__inst_inst_inst_add_3_43  ) + ( Xd_0__inst_inst_inst_add_3_42  ))
// Xd_0__inst_inst_inst_add_3_47  = SHARE((!Xd_0__inst_inst_first_level_4__11__q  & (Xd_0__inst_inst_first_level_3__11__q  & Xd_0__inst_inst_first_level_5__11__q )) # (Xd_0__inst_inst_first_level_4__11__q  & ((Xd_0__inst_inst_first_level_5__11__q ) # 
// (Xd_0__inst_inst_first_level_3__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__11__q ),
	.datac(!Xd_0__inst_inst_first_level_3__11__q ),
	.datad(!Xd_0__inst_inst_first_level_5__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_42 ),
	.sharein(Xd_0__inst_inst_inst_add_3_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_45_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_46 ),
	.shareout(Xd_0__inst_inst_inst_add_3_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_46  = CARRY(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_47  = SHARE((!Xd_0__inst_inst_first_level_2__11__q  & (Xd_0__inst_inst_first_level_1__11__q  & Xd_0__inst_inst_first_level_0__11__q )) # (Xd_0__inst_inst_first_level_2__11__q  & ((Xd_0__inst_inst_first_level_0__11__q ) # 
// (Xd_0__inst_inst_first_level_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__11__q ),
	.datac(!Xd_0__inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_49 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__12__q  $ (!Xd_0__inst_inst_first_level_3__12__q  $ (Xd_0__inst_inst_first_level_5__12__q )) ) + ( Xd_0__inst_inst_inst_add_3_47  ) + ( Xd_0__inst_inst_inst_add_3_46  ))
// Xd_0__inst_inst_inst_add_3_50  = CARRY(( !Xd_0__inst_inst_first_level_4__12__q  $ (!Xd_0__inst_inst_first_level_3__12__q  $ (Xd_0__inst_inst_first_level_5__12__q )) ) + ( Xd_0__inst_inst_inst_add_3_47  ) + ( Xd_0__inst_inst_inst_add_3_46  ))
// Xd_0__inst_inst_inst_add_3_51  = SHARE((!Xd_0__inst_inst_first_level_4__12__q  & (Xd_0__inst_inst_first_level_3__12__q  & Xd_0__inst_inst_first_level_5__12__q )) # (Xd_0__inst_inst_first_level_4__12__q  & ((Xd_0__inst_inst_first_level_5__12__q ) # 
// (Xd_0__inst_inst_first_level_3__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__12__q ),
	.datac(!Xd_0__inst_inst_first_level_3__12__q ),
	.datad(!Xd_0__inst_inst_first_level_5__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_46 ),
	.sharein(Xd_0__inst_inst_inst_add_3_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_49_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_50 ),
	.shareout(Xd_0__inst_inst_inst_add_3_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_50  = CARRY(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_51  = SHARE((!Xd_0__inst_inst_first_level_2__12__q  & (Xd_0__inst_inst_first_level_1__12__q  & Xd_0__inst_inst_first_level_0__12__q )) # (Xd_0__inst_inst_first_level_2__12__q  & ((Xd_0__inst_inst_first_level_0__12__q ) # 
// (Xd_0__inst_inst_first_level_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__12__q ),
	.datac(!Xd_0__inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_53 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_51  ) + ( Xd_0__inst_inst_inst_add_3_50  ))
// Xd_0__inst_inst_inst_add_3_54  = CARRY(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_51  ) + ( Xd_0__inst_inst_inst_add_3_50  ))
// Xd_0__inst_inst_inst_add_3_55  = SHARE((!Xd_0__inst_inst_first_level_4__13__q  & (Xd_0__inst_inst_first_level_3__13__q  & Xd_0__inst_inst_first_level_5__15__q )) # (Xd_0__inst_inst_first_level_4__13__q  & ((Xd_0__inst_inst_first_level_5__15__q ) # 
// (Xd_0__inst_inst_first_level_3__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__13__q ),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_5__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_50 ),
	.sharein(Xd_0__inst_inst_inst_add_3_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_53_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_54 ),
	.shareout(Xd_0__inst_inst_inst_add_3_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_54  = CARRY(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_55  = SHARE((!Xd_0__inst_inst_first_level_2__13__q  & (Xd_0__inst_inst_first_level_1__13__q  & Xd_0__inst_inst_first_level_0__13__q )) # (Xd_0__inst_inst_first_level_2__13__q  & ((Xd_0__inst_inst_first_level_0__13__q ) # 
// (Xd_0__inst_inst_first_level_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__13__q ),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_57 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__14__q  $ (!Xd_0__inst_inst_first_level_3__14__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_55  ) + ( Xd_0__inst_inst_inst_add_3_54  ))
// Xd_0__inst_inst_inst_add_3_58  = CARRY(( !Xd_0__inst_inst_first_level_4__14__q  $ (!Xd_0__inst_inst_first_level_3__14__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_55  ) + ( Xd_0__inst_inst_inst_add_3_54  ))
// Xd_0__inst_inst_inst_add_3_59  = SHARE((!Xd_0__inst_inst_first_level_4__14__q  & (Xd_0__inst_inst_first_level_3__14__q  & Xd_0__inst_inst_first_level_5__15__q )) # (Xd_0__inst_inst_first_level_4__14__q  & ((Xd_0__inst_inst_first_level_5__15__q ) # 
// (Xd_0__inst_inst_first_level_3__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__14__q ),
	.datac(!Xd_0__inst_inst_first_level_3__14__q ),
	.datad(!Xd_0__inst_inst_first_level_5__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_54 ),
	.sharein(Xd_0__inst_inst_inst_add_3_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_57_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_58 ),
	.shareout(Xd_0__inst_inst_inst_add_3_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q  $ (Xd_0__inst_inst_first_level_0__14__q )) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_58  = CARRY(( !Xd_0__inst_inst_first_level_2__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q  $ (Xd_0__inst_inst_first_level_0__14__q )) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_59  = SHARE((!Xd_0__inst_inst_first_level_2__14__q  & (Xd_0__inst_inst_first_level_1__14__q  & Xd_0__inst_inst_first_level_0__14__q )) # (Xd_0__inst_inst_first_level_2__14__q  & ((Xd_0__inst_inst_first_level_0__14__q ) # 
// (Xd_0__inst_inst_first_level_1__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__14__q ),
	.datac(!Xd_0__inst_inst_first_level_1__14__q ),
	.datad(!Xd_0__inst_inst_first_level_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_61 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__15__q  $ (!Xd_0__inst_inst_first_level_3__15__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_59  ) + ( Xd_0__inst_inst_inst_add_3_58  ))
// Xd_0__inst_inst_inst_add_3_62  = CARRY(( !Xd_0__inst_inst_first_level_4__15__q  $ (!Xd_0__inst_inst_first_level_3__15__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_59  ) + ( Xd_0__inst_inst_inst_add_3_58  ))
// Xd_0__inst_inst_inst_add_3_63  = SHARE((!Xd_0__inst_inst_first_level_4__15__q  & (Xd_0__inst_inst_first_level_3__15__q  & Xd_0__inst_inst_first_level_5__15__q )) # (Xd_0__inst_inst_first_level_4__15__q  & ((Xd_0__inst_inst_first_level_5__15__q ) # 
// (Xd_0__inst_inst_first_level_3__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__15__q ),
	.datac(!Xd_0__inst_inst_first_level_3__15__q ),
	.datad(!Xd_0__inst_inst_first_level_5__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_58 ),
	.sharein(Xd_0__inst_inst_inst_add_3_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_62 ),
	.shareout(Xd_0__inst_inst_inst_add_3_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_add_0_58  ))
// Xd_0__inst_inst_inst_add_0_62  = CARRY(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_add_0_58  ))
// Xd_0__inst_inst_inst_add_0_63  = SHARE((!Xd_0__inst_inst_first_level_2__15__q  & (Xd_0__inst_inst_first_level_1__15__q  & Xd_0__inst_inst_first_level_0__15__q )) # (Xd_0__inst_inst_first_level_2__15__q  & ((Xd_0__inst_inst_first_level_0__15__q ) # 
// (Xd_0__inst_inst_first_level_1__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__15__q ),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_62 ),
	.shareout(Xd_0__inst_inst_inst_add_0_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_65 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_65_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__15__q  $ (!Xd_0__inst_inst_first_level_3__15__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_63  ) + ( Xd_0__inst_inst_inst_add_3_62  ))
// Xd_0__inst_inst_inst_add_3_66  = CARRY(( !Xd_0__inst_inst_first_level_4__15__q  $ (!Xd_0__inst_inst_first_level_3__15__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_63  ) + ( Xd_0__inst_inst_inst_add_3_62  ))
// Xd_0__inst_inst_inst_add_3_67  = SHARE((!Xd_0__inst_inst_first_level_4__15__q  & (Xd_0__inst_inst_first_level_3__15__q  & Xd_0__inst_inst_first_level_5__15__q )) # (Xd_0__inst_inst_first_level_4__15__q  & ((Xd_0__inst_inst_first_level_5__15__q ) # 
// (Xd_0__inst_inst_first_level_3__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__15__q ),
	.datac(!Xd_0__inst_inst_first_level_3__15__q ),
	.datad(!Xd_0__inst_inst_first_level_5__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_62 ),
	.sharein(Xd_0__inst_inst_inst_add_3_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_65_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_66 ),
	.shareout(Xd_0__inst_inst_inst_add_3_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_65 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_65_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_add_0_63  ) + ( Xd_0__inst_inst_inst_add_0_62  ))
// Xd_0__inst_inst_inst_add_0_66  = CARRY(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_add_0_63  ) + ( Xd_0__inst_inst_inst_add_0_62  ))
// Xd_0__inst_inst_inst_add_0_67  = SHARE((!Xd_0__inst_inst_first_level_2__15__q  & (Xd_0__inst_inst_first_level_1__15__q  & Xd_0__inst_inst_first_level_0__15__q )) # (Xd_0__inst_inst_first_level_2__15__q  & ((Xd_0__inst_inst_first_level_0__15__q ) # 
// (Xd_0__inst_inst_first_level_1__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__15__q ),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_62 ),
	.sharein(Xd_0__inst_inst_inst_add_0_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_65_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_66 ),
	.shareout(Xd_0__inst_inst_inst_add_0_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_69 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_69_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__15__q  $ (!Xd_0__inst_inst_first_level_3__15__q  $ (Xd_0__inst_inst_first_level_5__15__q )) ) + ( Xd_0__inst_inst_inst_add_3_67  ) + ( Xd_0__inst_inst_inst_add_3_66  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__15__q ),
	.datac(!Xd_0__inst_inst_first_level_3__15__q ),
	.datad(!Xd_0__inst_inst_first_level_5__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_66 ),
	.sharein(Xd_0__inst_inst_inst_add_3_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_69_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_69 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_69_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q  $ (Xd_0__inst_inst_first_level_0__15__q )) ) + ( Xd_0__inst_inst_inst_add_0_67  ) + ( Xd_0__inst_inst_inst_add_0_66  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__15__q ),
	.datac(!Xd_0__inst_inst_first_level_1__15__q ),
	.datad(!Xd_0__inst_inst_first_level_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_66 ),
	.sharein(Xd_0__inst_inst_inst_add_0_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_69_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_9 (
// Equation(s):
// Xd_0__inst_i19_9_sumout  = SUM(( !din_a[125] $ (!din_b[125]) ) + ( Xd_0__inst_i19_19  ) + ( Xd_0__inst_i19_18  ))
// Xd_0__inst_i19_10  = CARRY(( !din_a[125] $ (!din_b[125]) ) + ( Xd_0__inst_i19_19  ) + ( Xd_0__inst_i19_18  ))
// Xd_0__inst_i19_11  = SHARE(GND)

	.dataa(!din_a[125]),
	.datab(!din_b[125]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_18 ),
	.sharein(Xd_0__inst_i19_19 ),
	.combout(),
	.sumout(Xd_0__inst_i19_9_sumout ),
	.cout(Xd_0__inst_i19_10 ),
	.shareout(Xd_0__inst_i19_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_13 (
// Equation(s):
// Xd_0__inst_i19_13_sumout  = SUM(( !din_a[223] $ (!din_b[223]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_14  = CARRY(( !din_a[223] $ (!din_b[223]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_15  = SHARE(GND)

	.dataa(!din_a[223]),
	.datab(!din_b[223]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_13_sumout ),
	.cout(Xd_0__inst_i19_14 ),
	.shareout(Xd_0__inst_i19_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_1 (
// Equation(s):
// Xd_0__inst_inst_add_8_1_sumout  = SUM(( !Xd_0__inst_r_sum1_14__0__q  $ (!Xd_0__inst_r_sum1_13__0__q  $ (Xd_0__inst_r_sum1_12__0__q )) ) + ( Xd_0__inst_i19_23  ) + ( Xd_0__inst_i19_22  ))
// Xd_0__inst_inst_add_8_2  = CARRY(( !Xd_0__inst_r_sum1_14__0__q  $ (!Xd_0__inst_r_sum1_13__0__q  $ (Xd_0__inst_r_sum1_12__0__q )) ) + ( Xd_0__inst_i19_23  ) + ( Xd_0__inst_i19_22  ))
// Xd_0__inst_inst_add_8_3  = SHARE((!Xd_0__inst_r_sum1_14__0__q  & (Xd_0__inst_r_sum1_13__0__q  & Xd_0__inst_r_sum1_12__0__q )) # (Xd_0__inst_r_sum1_14__0__q  & ((Xd_0__inst_r_sum1_12__0__q ) # (Xd_0__inst_r_sum1_13__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__0__q ),
	.datac(!Xd_0__inst_r_sum1_13__0__q ),
	.datad(!Xd_0__inst_r_sum1_12__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_22 ),
	.sharein(Xd_0__inst_i19_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_1_sumout ),
	.cout(Xd_0__inst_inst_add_8_2 ),
	.shareout(Xd_0__inst_inst_add_8_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_1 (
// Equation(s):
// Xd_0__inst_inst_add_6_1_sumout  = SUM(( !Xd_0__inst_r_sum1_11__0__q  $ (!Xd_0__inst_r_sum1_10__0__q  $ (Xd_0__inst_r_sum1_9__0__q )) ) + ( Xd_0__inst_i19_27  ) + ( Xd_0__inst_i19_26  ))
// Xd_0__inst_inst_add_6_2  = CARRY(( !Xd_0__inst_r_sum1_11__0__q  $ (!Xd_0__inst_r_sum1_10__0__q  $ (Xd_0__inst_r_sum1_9__0__q )) ) + ( Xd_0__inst_i19_27  ) + ( Xd_0__inst_i19_26  ))
// Xd_0__inst_inst_add_6_3  = SHARE((!Xd_0__inst_r_sum1_11__0__q  & (Xd_0__inst_r_sum1_10__0__q  & Xd_0__inst_r_sum1_9__0__q )) # (Xd_0__inst_r_sum1_11__0__q  & ((Xd_0__inst_r_sum1_9__0__q ) # (Xd_0__inst_r_sum1_10__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__0__q ),
	.datac(!Xd_0__inst_r_sum1_10__0__q ),
	.datad(!Xd_0__inst_r_sum1_9__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_26 ),
	.sharein(Xd_0__inst_i19_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_1_sumout ),
	.cout(Xd_0__inst_inst_add_6_2 ),
	.shareout(Xd_0__inst_inst_add_6_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_17 (
// Equation(s):
// Xd_0__inst_i19_17_sumout  = SUM(( !din_a[216] $ (!din_b[216]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_18  = CARRY(( !din_a[216] $ (!din_b[216]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_19  = SHARE(GND)

	.dataa(!din_a[216]),
	.datab(!din_b[216]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_17_sumout ),
	.cout(Xd_0__inst_i19_18 ),
	.shareout(Xd_0__inst_i19_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_1 (
// Equation(s):
// Xd_0__inst_inst_add_4_1_sumout  = SUM(( !Xd_0__inst_r_sum1_8__0__q  $ (!Xd_0__inst_r_sum1_7__0__q  $ (Xd_0__inst_r_sum1_6__0__q )) ) + ( Xd_0__inst_i19_31  ) + ( Xd_0__inst_i19_30  ))
// Xd_0__inst_inst_add_4_2  = CARRY(( !Xd_0__inst_r_sum1_8__0__q  $ (!Xd_0__inst_r_sum1_7__0__q  $ (Xd_0__inst_r_sum1_6__0__q )) ) + ( Xd_0__inst_i19_31  ) + ( Xd_0__inst_i19_30  ))
// Xd_0__inst_inst_add_4_3  = SHARE((!Xd_0__inst_r_sum1_8__0__q  & (Xd_0__inst_r_sum1_7__0__q  & Xd_0__inst_r_sum1_6__0__q )) # (Xd_0__inst_r_sum1_8__0__q  & ((Xd_0__inst_r_sum1_6__0__q ) # (Xd_0__inst_r_sum1_7__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__0__q ),
	.datac(!Xd_0__inst_r_sum1_7__0__q ),
	.datad(!Xd_0__inst_r_sum1_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_30 ),
	.sharein(Xd_0__inst_i19_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_1_sumout ),
	.cout(Xd_0__inst_inst_add_4_2 ),
	.shareout(Xd_0__inst_inst_add_4_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_1 (
// Equation(s):
// Xd_0__inst_inst_add_2_1_sumout  = SUM(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_i19_35  ) + ( Xd_0__inst_i19_34  ))
// Xd_0__inst_inst_add_2_2  = CARRY(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_i19_35  ) + ( Xd_0__inst_i19_34  ))
// Xd_0__inst_inst_add_2_3  = SHARE((!Xd_0__inst_r_sum1_5__0__q  & (Xd_0__inst_r_sum1_4__0__q  & Xd_0__inst_r_sum1_3__0__q )) # (Xd_0__inst_r_sum1_5__0__q  & ((Xd_0__inst_r_sum1_3__0__q ) # (Xd_0__inst_r_sum1_4__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__0__q ),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sum1_3__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_34 ),
	.sharein(Xd_0__inst_i19_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_1_sumout ),
	.cout(Xd_0__inst_inst_add_2_2 ),
	.shareout(Xd_0__inst_inst_add_2_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_i19_39  ) + ( Xd_0__inst_i19_38  ))
// Xd_0__inst_inst_add_0_2  = CARRY(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_i19_39  ) + ( Xd_0__inst_i19_38  ))
// Xd_0__inst_inst_add_0_3  = SHARE((!Xd_0__inst_r_sum1_2__0__q  & (Xd_0__inst_r_sum1_1__0__q  & Xd_0__inst_r_sum1_0__0__q )) # (Xd_0__inst_r_sum1_2__0__q  & ((Xd_0__inst_r_sum1_0__0__q ) # (Xd_0__inst_r_sum1_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__0__q ),
	.datac(!Xd_0__inst_r_sum1_1__0__q ),
	.datad(!Xd_0__inst_r_sum1_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_38 ),
	.sharein(Xd_0__inst_i19_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_5 (
// Equation(s):
// Xd_0__inst_inst_add_8_5_sumout  = SUM(( !Xd_0__inst_r_sum1_14__1__q  $ (!Xd_0__inst_r_sum1_13__1__q  $ (Xd_0__inst_r_sum1_12__1__q )) ) + ( Xd_0__inst_inst_add_8_3  ) + ( Xd_0__inst_inst_add_8_2  ))
// Xd_0__inst_inst_add_8_6  = CARRY(( !Xd_0__inst_r_sum1_14__1__q  $ (!Xd_0__inst_r_sum1_13__1__q  $ (Xd_0__inst_r_sum1_12__1__q )) ) + ( Xd_0__inst_inst_add_8_3  ) + ( Xd_0__inst_inst_add_8_2  ))
// Xd_0__inst_inst_add_8_7  = SHARE((!Xd_0__inst_r_sum1_14__1__q  & (Xd_0__inst_r_sum1_13__1__q  & Xd_0__inst_r_sum1_12__1__q )) # (Xd_0__inst_r_sum1_14__1__q  & ((Xd_0__inst_r_sum1_12__1__q ) # (Xd_0__inst_r_sum1_13__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__1__q ),
	.datac(!Xd_0__inst_r_sum1_13__1__q ),
	.datad(!Xd_0__inst_r_sum1_12__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_2 ),
	.sharein(Xd_0__inst_inst_add_8_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_5_sumout ),
	.cout(Xd_0__inst_inst_add_8_6 ),
	.shareout(Xd_0__inst_inst_add_8_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_5 (
// Equation(s):
// Xd_0__inst_inst_add_6_5_sumout  = SUM(( !Xd_0__inst_r_sum1_11__1__q  $ (!Xd_0__inst_r_sum1_10__1__q  $ (Xd_0__inst_r_sum1_9__1__q )) ) + ( Xd_0__inst_inst_add_6_3  ) + ( Xd_0__inst_inst_add_6_2  ))
// Xd_0__inst_inst_add_6_6  = CARRY(( !Xd_0__inst_r_sum1_11__1__q  $ (!Xd_0__inst_r_sum1_10__1__q  $ (Xd_0__inst_r_sum1_9__1__q )) ) + ( Xd_0__inst_inst_add_6_3  ) + ( Xd_0__inst_inst_add_6_2  ))
// Xd_0__inst_inst_add_6_7  = SHARE((!Xd_0__inst_r_sum1_11__1__q  & (Xd_0__inst_r_sum1_10__1__q  & Xd_0__inst_r_sum1_9__1__q )) # (Xd_0__inst_r_sum1_11__1__q  & ((Xd_0__inst_r_sum1_9__1__q ) # (Xd_0__inst_r_sum1_10__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__1__q ),
	.datac(!Xd_0__inst_r_sum1_10__1__q ),
	.datad(!Xd_0__inst_r_sum1_9__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_2 ),
	.sharein(Xd_0__inst_inst_add_6_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_5_sumout ),
	.cout(Xd_0__inst_inst_add_6_6 ),
	.shareout(Xd_0__inst_inst_add_6_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_5 (
// Equation(s):
// Xd_0__inst_inst_add_4_5_sumout  = SUM(( !Xd_0__inst_r_sum1_8__1__q  $ (!Xd_0__inst_r_sum1_7__1__q  $ (Xd_0__inst_r_sum1_6__1__q )) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_6  = CARRY(( !Xd_0__inst_r_sum1_8__1__q  $ (!Xd_0__inst_r_sum1_7__1__q  $ (Xd_0__inst_r_sum1_6__1__q )) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_7  = SHARE((!Xd_0__inst_r_sum1_8__1__q  & (Xd_0__inst_r_sum1_7__1__q  & Xd_0__inst_r_sum1_6__1__q )) # (Xd_0__inst_r_sum1_8__1__q  & ((Xd_0__inst_r_sum1_6__1__q ) # (Xd_0__inst_r_sum1_7__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__1__q ),
	.datac(!Xd_0__inst_r_sum1_7__1__q ),
	.datad(!Xd_0__inst_r_sum1_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_2 ),
	.sharein(Xd_0__inst_inst_add_4_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_5_sumout ),
	.cout(Xd_0__inst_inst_add_4_6 ),
	.shareout(Xd_0__inst_inst_add_4_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_5 (
// Equation(s):
// Xd_0__inst_inst_add_2_5_sumout  = SUM(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_6  = CARRY(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_7  = SHARE((!Xd_0__inst_r_sum1_5__1__q  & (Xd_0__inst_r_sum1_4__1__q  & Xd_0__inst_r_sum1_3__1__q )) # (Xd_0__inst_r_sum1_5__1__q  & ((Xd_0__inst_r_sum1_3__1__q ) # (Xd_0__inst_r_sum1_4__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__1__q ),
	.datac(!Xd_0__inst_r_sum1_4__1__q ),
	.datad(!Xd_0__inst_r_sum1_3__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_2 ),
	.sharein(Xd_0__inst_inst_add_2_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_5_sumout ),
	.cout(Xd_0__inst_inst_add_2_6 ),
	.shareout(Xd_0__inst_inst_add_2_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_6  = CARRY(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_7  = SHARE((!Xd_0__inst_r_sum1_2__1__q  & (Xd_0__inst_r_sum1_1__1__q  & Xd_0__inst_r_sum1_0__1__q )) # (Xd_0__inst_r_sum1_2__1__q  & ((Xd_0__inst_r_sum1_0__1__q ) # (Xd_0__inst_r_sum1_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__1__q ),
	.datad(!Xd_0__inst_r_sum1_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_9 (
// Equation(s):
// Xd_0__inst_inst_add_8_9_sumout  = SUM(( !Xd_0__inst_r_sum1_14__2__q  $ (!Xd_0__inst_r_sum1_13__2__q  $ (Xd_0__inst_r_sum1_12__2__q )) ) + ( Xd_0__inst_inst_add_8_7  ) + ( Xd_0__inst_inst_add_8_6  ))
// Xd_0__inst_inst_add_8_10  = CARRY(( !Xd_0__inst_r_sum1_14__2__q  $ (!Xd_0__inst_r_sum1_13__2__q  $ (Xd_0__inst_r_sum1_12__2__q )) ) + ( Xd_0__inst_inst_add_8_7  ) + ( Xd_0__inst_inst_add_8_6  ))
// Xd_0__inst_inst_add_8_11  = SHARE((!Xd_0__inst_r_sum1_14__2__q  & (Xd_0__inst_r_sum1_13__2__q  & Xd_0__inst_r_sum1_12__2__q )) # (Xd_0__inst_r_sum1_14__2__q  & ((Xd_0__inst_r_sum1_12__2__q ) # (Xd_0__inst_r_sum1_13__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__2__q ),
	.datac(!Xd_0__inst_r_sum1_13__2__q ),
	.datad(!Xd_0__inst_r_sum1_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_6 ),
	.sharein(Xd_0__inst_inst_add_8_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_9_sumout ),
	.cout(Xd_0__inst_inst_add_8_10 ),
	.shareout(Xd_0__inst_inst_add_8_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_9 (
// Equation(s):
// Xd_0__inst_inst_add_6_9_sumout  = SUM(( !Xd_0__inst_r_sum1_11__2__q  $ (!Xd_0__inst_r_sum1_10__2__q  $ (Xd_0__inst_r_sum1_9__2__q )) ) + ( Xd_0__inst_inst_add_6_7  ) + ( Xd_0__inst_inst_add_6_6  ))
// Xd_0__inst_inst_add_6_10  = CARRY(( !Xd_0__inst_r_sum1_11__2__q  $ (!Xd_0__inst_r_sum1_10__2__q  $ (Xd_0__inst_r_sum1_9__2__q )) ) + ( Xd_0__inst_inst_add_6_7  ) + ( Xd_0__inst_inst_add_6_6  ))
// Xd_0__inst_inst_add_6_11  = SHARE((!Xd_0__inst_r_sum1_11__2__q  & (Xd_0__inst_r_sum1_10__2__q  & Xd_0__inst_r_sum1_9__2__q )) # (Xd_0__inst_r_sum1_11__2__q  & ((Xd_0__inst_r_sum1_9__2__q ) # (Xd_0__inst_r_sum1_10__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__2__q ),
	.datac(!Xd_0__inst_r_sum1_10__2__q ),
	.datad(!Xd_0__inst_r_sum1_9__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_6 ),
	.sharein(Xd_0__inst_inst_add_6_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_9_sumout ),
	.cout(Xd_0__inst_inst_add_6_10 ),
	.shareout(Xd_0__inst_inst_add_6_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_9 (
// Equation(s):
// Xd_0__inst_inst_add_4_9_sumout  = SUM(( !Xd_0__inst_r_sum1_8__2__q  $ (!Xd_0__inst_r_sum1_7__2__q  $ (Xd_0__inst_r_sum1_6__2__q )) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_10  = CARRY(( !Xd_0__inst_r_sum1_8__2__q  $ (!Xd_0__inst_r_sum1_7__2__q  $ (Xd_0__inst_r_sum1_6__2__q )) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_11  = SHARE((!Xd_0__inst_r_sum1_8__2__q  & (Xd_0__inst_r_sum1_7__2__q  & Xd_0__inst_r_sum1_6__2__q )) # (Xd_0__inst_r_sum1_8__2__q  & ((Xd_0__inst_r_sum1_6__2__q ) # (Xd_0__inst_r_sum1_7__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__2__q ),
	.datac(!Xd_0__inst_r_sum1_7__2__q ),
	.datad(!Xd_0__inst_r_sum1_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_6 ),
	.sharein(Xd_0__inst_inst_add_4_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_9_sumout ),
	.cout(Xd_0__inst_inst_add_4_10 ),
	.shareout(Xd_0__inst_inst_add_4_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_9 (
// Equation(s):
// Xd_0__inst_inst_add_2_9_sumout  = SUM(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_10  = CARRY(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_11  = SHARE((!Xd_0__inst_r_sum1_5__2__q  & (Xd_0__inst_r_sum1_4__2__q  & Xd_0__inst_r_sum1_3__2__q )) # (Xd_0__inst_r_sum1_5__2__q  & ((Xd_0__inst_r_sum1_3__2__q ) # (Xd_0__inst_r_sum1_4__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__2__q ),
	.datac(!Xd_0__inst_r_sum1_4__2__q ),
	.datad(!Xd_0__inst_r_sum1_3__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_6 ),
	.sharein(Xd_0__inst_inst_add_2_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_9_sumout ),
	.cout(Xd_0__inst_inst_add_2_10 ),
	.shareout(Xd_0__inst_inst_add_2_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_10  = CARRY(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_11  = SHARE((!Xd_0__inst_r_sum1_2__2__q  & (Xd_0__inst_r_sum1_1__2__q  & Xd_0__inst_r_sum1_0__2__q )) # (Xd_0__inst_r_sum1_2__2__q  & ((Xd_0__inst_r_sum1_0__2__q ) # (Xd_0__inst_r_sum1_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__2__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_13 (
// Equation(s):
// Xd_0__inst_inst_add_8_13_sumout  = SUM(( !Xd_0__inst_r_sum1_14__3__q  $ (!Xd_0__inst_r_sum1_13__3__q  $ (Xd_0__inst_r_sum1_12__3__q )) ) + ( Xd_0__inst_inst_add_8_11  ) + ( Xd_0__inst_inst_add_8_10  ))
// Xd_0__inst_inst_add_8_14  = CARRY(( !Xd_0__inst_r_sum1_14__3__q  $ (!Xd_0__inst_r_sum1_13__3__q  $ (Xd_0__inst_r_sum1_12__3__q )) ) + ( Xd_0__inst_inst_add_8_11  ) + ( Xd_0__inst_inst_add_8_10  ))
// Xd_0__inst_inst_add_8_15  = SHARE((!Xd_0__inst_r_sum1_14__3__q  & (Xd_0__inst_r_sum1_13__3__q  & Xd_0__inst_r_sum1_12__3__q )) # (Xd_0__inst_r_sum1_14__3__q  & ((Xd_0__inst_r_sum1_12__3__q ) # (Xd_0__inst_r_sum1_13__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__3__q ),
	.datac(!Xd_0__inst_r_sum1_13__3__q ),
	.datad(!Xd_0__inst_r_sum1_12__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_10 ),
	.sharein(Xd_0__inst_inst_add_8_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_13_sumout ),
	.cout(Xd_0__inst_inst_add_8_14 ),
	.shareout(Xd_0__inst_inst_add_8_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_13 (
// Equation(s):
// Xd_0__inst_inst_add_6_13_sumout  = SUM(( !Xd_0__inst_r_sum1_11__3__q  $ (!Xd_0__inst_r_sum1_10__3__q  $ (Xd_0__inst_r_sum1_9__3__q )) ) + ( Xd_0__inst_inst_add_6_11  ) + ( Xd_0__inst_inst_add_6_10  ))
// Xd_0__inst_inst_add_6_14  = CARRY(( !Xd_0__inst_r_sum1_11__3__q  $ (!Xd_0__inst_r_sum1_10__3__q  $ (Xd_0__inst_r_sum1_9__3__q )) ) + ( Xd_0__inst_inst_add_6_11  ) + ( Xd_0__inst_inst_add_6_10  ))
// Xd_0__inst_inst_add_6_15  = SHARE((!Xd_0__inst_r_sum1_11__3__q  & (Xd_0__inst_r_sum1_10__3__q  & Xd_0__inst_r_sum1_9__3__q )) # (Xd_0__inst_r_sum1_11__3__q  & ((Xd_0__inst_r_sum1_9__3__q ) # (Xd_0__inst_r_sum1_10__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__3__q ),
	.datac(!Xd_0__inst_r_sum1_10__3__q ),
	.datad(!Xd_0__inst_r_sum1_9__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_10 ),
	.sharein(Xd_0__inst_inst_add_6_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_13_sumout ),
	.cout(Xd_0__inst_inst_add_6_14 ),
	.shareout(Xd_0__inst_inst_add_6_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_13 (
// Equation(s):
// Xd_0__inst_inst_add_4_13_sumout  = SUM(( !Xd_0__inst_r_sum1_8__3__q  $ (!Xd_0__inst_r_sum1_7__3__q  $ (Xd_0__inst_r_sum1_6__3__q )) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_14  = CARRY(( !Xd_0__inst_r_sum1_8__3__q  $ (!Xd_0__inst_r_sum1_7__3__q  $ (Xd_0__inst_r_sum1_6__3__q )) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_15  = SHARE((!Xd_0__inst_r_sum1_8__3__q  & (Xd_0__inst_r_sum1_7__3__q  & Xd_0__inst_r_sum1_6__3__q )) # (Xd_0__inst_r_sum1_8__3__q  & ((Xd_0__inst_r_sum1_6__3__q ) # (Xd_0__inst_r_sum1_7__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__3__q ),
	.datac(!Xd_0__inst_r_sum1_7__3__q ),
	.datad(!Xd_0__inst_r_sum1_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_10 ),
	.sharein(Xd_0__inst_inst_add_4_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_13_sumout ),
	.cout(Xd_0__inst_inst_add_4_14 ),
	.shareout(Xd_0__inst_inst_add_4_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_13 (
// Equation(s):
// Xd_0__inst_inst_add_2_13_sumout  = SUM(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_14  = CARRY(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_15  = SHARE((!Xd_0__inst_r_sum1_5__3__q  & (Xd_0__inst_r_sum1_4__3__q  & Xd_0__inst_r_sum1_3__3__q )) # (Xd_0__inst_r_sum1_5__3__q  & ((Xd_0__inst_r_sum1_3__3__q ) # (Xd_0__inst_r_sum1_4__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__3__q ),
	.datac(!Xd_0__inst_r_sum1_4__3__q ),
	.datad(!Xd_0__inst_r_sum1_3__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_10 ),
	.sharein(Xd_0__inst_inst_add_2_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_13_sumout ),
	.cout(Xd_0__inst_inst_add_2_14 ),
	.shareout(Xd_0__inst_inst_add_2_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_14  = CARRY(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_15  = SHARE((!Xd_0__inst_r_sum1_2__3__q  & (Xd_0__inst_r_sum1_1__3__q  & Xd_0__inst_r_sum1_0__3__q )) # (Xd_0__inst_r_sum1_2__3__q  & ((Xd_0__inst_r_sum1_0__3__q ) # (Xd_0__inst_r_sum1_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__3__q ),
	.datad(!Xd_0__inst_r_sum1_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_17 (
// Equation(s):
// Xd_0__inst_inst_add_8_17_sumout  = SUM(( !Xd_0__inst_r_sum1_14__4__q  $ (!Xd_0__inst_r_sum1_13__4__q  $ (Xd_0__inst_r_sum1_12__4__q )) ) + ( Xd_0__inst_inst_add_8_15  ) + ( Xd_0__inst_inst_add_8_14  ))
// Xd_0__inst_inst_add_8_18  = CARRY(( !Xd_0__inst_r_sum1_14__4__q  $ (!Xd_0__inst_r_sum1_13__4__q  $ (Xd_0__inst_r_sum1_12__4__q )) ) + ( Xd_0__inst_inst_add_8_15  ) + ( Xd_0__inst_inst_add_8_14  ))
// Xd_0__inst_inst_add_8_19  = SHARE((!Xd_0__inst_r_sum1_14__4__q  & (Xd_0__inst_r_sum1_13__4__q  & Xd_0__inst_r_sum1_12__4__q )) # (Xd_0__inst_r_sum1_14__4__q  & ((Xd_0__inst_r_sum1_12__4__q ) # (Xd_0__inst_r_sum1_13__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__4__q ),
	.datac(!Xd_0__inst_r_sum1_13__4__q ),
	.datad(!Xd_0__inst_r_sum1_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_14 ),
	.sharein(Xd_0__inst_inst_add_8_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_17_sumout ),
	.cout(Xd_0__inst_inst_add_8_18 ),
	.shareout(Xd_0__inst_inst_add_8_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_17 (
// Equation(s):
// Xd_0__inst_inst_add_6_17_sumout  = SUM(( !Xd_0__inst_r_sum1_11__4__q  $ (!Xd_0__inst_r_sum1_10__4__q  $ (Xd_0__inst_r_sum1_9__4__q )) ) + ( Xd_0__inst_inst_add_6_15  ) + ( Xd_0__inst_inst_add_6_14  ))
// Xd_0__inst_inst_add_6_18  = CARRY(( !Xd_0__inst_r_sum1_11__4__q  $ (!Xd_0__inst_r_sum1_10__4__q  $ (Xd_0__inst_r_sum1_9__4__q )) ) + ( Xd_0__inst_inst_add_6_15  ) + ( Xd_0__inst_inst_add_6_14  ))
// Xd_0__inst_inst_add_6_19  = SHARE((!Xd_0__inst_r_sum1_11__4__q  & (Xd_0__inst_r_sum1_10__4__q  & Xd_0__inst_r_sum1_9__4__q )) # (Xd_0__inst_r_sum1_11__4__q  & ((Xd_0__inst_r_sum1_9__4__q ) # (Xd_0__inst_r_sum1_10__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__4__q ),
	.datac(!Xd_0__inst_r_sum1_10__4__q ),
	.datad(!Xd_0__inst_r_sum1_9__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_14 ),
	.sharein(Xd_0__inst_inst_add_6_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_17_sumout ),
	.cout(Xd_0__inst_inst_add_6_18 ),
	.shareout(Xd_0__inst_inst_add_6_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_17 (
// Equation(s):
// Xd_0__inst_inst_add_4_17_sumout  = SUM(( !Xd_0__inst_r_sum1_8__4__q  $ (!Xd_0__inst_r_sum1_7__4__q  $ (Xd_0__inst_r_sum1_6__4__q )) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_18  = CARRY(( !Xd_0__inst_r_sum1_8__4__q  $ (!Xd_0__inst_r_sum1_7__4__q  $ (Xd_0__inst_r_sum1_6__4__q )) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_19  = SHARE((!Xd_0__inst_r_sum1_8__4__q  & (Xd_0__inst_r_sum1_7__4__q  & Xd_0__inst_r_sum1_6__4__q )) # (Xd_0__inst_r_sum1_8__4__q  & ((Xd_0__inst_r_sum1_6__4__q ) # (Xd_0__inst_r_sum1_7__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__4__q ),
	.datac(!Xd_0__inst_r_sum1_7__4__q ),
	.datad(!Xd_0__inst_r_sum1_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_14 ),
	.sharein(Xd_0__inst_inst_add_4_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_17_sumout ),
	.cout(Xd_0__inst_inst_add_4_18 ),
	.shareout(Xd_0__inst_inst_add_4_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_17 (
// Equation(s):
// Xd_0__inst_inst_add_2_17_sumout  = SUM(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_18  = CARRY(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_19  = SHARE((!Xd_0__inst_r_sum1_5__4__q  & (Xd_0__inst_r_sum1_4__4__q  & Xd_0__inst_r_sum1_3__4__q )) # (Xd_0__inst_r_sum1_5__4__q  & ((Xd_0__inst_r_sum1_3__4__q ) # (Xd_0__inst_r_sum1_4__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__4__q ),
	.datac(!Xd_0__inst_r_sum1_4__4__q ),
	.datad(!Xd_0__inst_r_sum1_3__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_14 ),
	.sharein(Xd_0__inst_inst_add_2_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_17_sumout ),
	.cout(Xd_0__inst_inst_add_2_18 ),
	.shareout(Xd_0__inst_inst_add_2_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_18  = CARRY(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_19  = SHARE((!Xd_0__inst_r_sum1_2__4__q  & (Xd_0__inst_r_sum1_1__4__q  & Xd_0__inst_r_sum1_0__4__q )) # (Xd_0__inst_r_sum1_2__4__q  & ((Xd_0__inst_r_sum1_0__4__q ) # (Xd_0__inst_r_sum1_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__4__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_21 (
// Equation(s):
// Xd_0__inst_inst_add_8_21_sumout  = SUM(( !Xd_0__inst_r_sum1_14__5__q  $ (!Xd_0__inst_r_sum1_13__5__q  $ (Xd_0__inst_r_sum1_12__5__q )) ) + ( Xd_0__inst_inst_add_8_19  ) + ( Xd_0__inst_inst_add_8_18  ))
// Xd_0__inst_inst_add_8_22  = CARRY(( !Xd_0__inst_r_sum1_14__5__q  $ (!Xd_0__inst_r_sum1_13__5__q  $ (Xd_0__inst_r_sum1_12__5__q )) ) + ( Xd_0__inst_inst_add_8_19  ) + ( Xd_0__inst_inst_add_8_18  ))
// Xd_0__inst_inst_add_8_23  = SHARE((!Xd_0__inst_r_sum1_14__5__q  & (Xd_0__inst_r_sum1_13__5__q  & Xd_0__inst_r_sum1_12__5__q )) # (Xd_0__inst_r_sum1_14__5__q  & ((Xd_0__inst_r_sum1_12__5__q ) # (Xd_0__inst_r_sum1_13__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__5__q ),
	.datac(!Xd_0__inst_r_sum1_13__5__q ),
	.datad(!Xd_0__inst_r_sum1_12__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_18 ),
	.sharein(Xd_0__inst_inst_add_8_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_21_sumout ),
	.cout(Xd_0__inst_inst_add_8_22 ),
	.shareout(Xd_0__inst_inst_add_8_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_21 (
// Equation(s):
// Xd_0__inst_inst_add_6_21_sumout  = SUM(( !Xd_0__inst_r_sum1_11__5__q  $ (!Xd_0__inst_r_sum1_10__5__q  $ (Xd_0__inst_r_sum1_9__5__q )) ) + ( Xd_0__inst_inst_add_6_19  ) + ( Xd_0__inst_inst_add_6_18  ))
// Xd_0__inst_inst_add_6_22  = CARRY(( !Xd_0__inst_r_sum1_11__5__q  $ (!Xd_0__inst_r_sum1_10__5__q  $ (Xd_0__inst_r_sum1_9__5__q )) ) + ( Xd_0__inst_inst_add_6_19  ) + ( Xd_0__inst_inst_add_6_18  ))
// Xd_0__inst_inst_add_6_23  = SHARE((!Xd_0__inst_r_sum1_11__5__q  & (Xd_0__inst_r_sum1_10__5__q  & Xd_0__inst_r_sum1_9__5__q )) # (Xd_0__inst_r_sum1_11__5__q  & ((Xd_0__inst_r_sum1_9__5__q ) # (Xd_0__inst_r_sum1_10__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__5__q ),
	.datac(!Xd_0__inst_r_sum1_10__5__q ),
	.datad(!Xd_0__inst_r_sum1_9__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_18 ),
	.sharein(Xd_0__inst_inst_add_6_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_21_sumout ),
	.cout(Xd_0__inst_inst_add_6_22 ),
	.shareout(Xd_0__inst_inst_add_6_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_21 (
// Equation(s):
// Xd_0__inst_inst_add_4_21_sumout  = SUM(( !Xd_0__inst_r_sum1_8__5__q  $ (!Xd_0__inst_r_sum1_7__5__q  $ (Xd_0__inst_r_sum1_6__5__q )) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_22  = CARRY(( !Xd_0__inst_r_sum1_8__5__q  $ (!Xd_0__inst_r_sum1_7__5__q  $ (Xd_0__inst_r_sum1_6__5__q )) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_23  = SHARE((!Xd_0__inst_r_sum1_8__5__q  & (Xd_0__inst_r_sum1_7__5__q  & Xd_0__inst_r_sum1_6__5__q )) # (Xd_0__inst_r_sum1_8__5__q  & ((Xd_0__inst_r_sum1_6__5__q ) # (Xd_0__inst_r_sum1_7__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__5__q ),
	.datac(!Xd_0__inst_r_sum1_7__5__q ),
	.datad(!Xd_0__inst_r_sum1_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_18 ),
	.sharein(Xd_0__inst_inst_add_4_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_21_sumout ),
	.cout(Xd_0__inst_inst_add_4_22 ),
	.shareout(Xd_0__inst_inst_add_4_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_21 (
// Equation(s):
// Xd_0__inst_inst_add_2_21_sumout  = SUM(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_22  = CARRY(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_23  = SHARE((!Xd_0__inst_r_sum1_5__5__q  & (Xd_0__inst_r_sum1_4__5__q  & Xd_0__inst_r_sum1_3__5__q )) # (Xd_0__inst_r_sum1_5__5__q  & ((Xd_0__inst_r_sum1_3__5__q ) # (Xd_0__inst_r_sum1_4__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__5__q ),
	.datac(!Xd_0__inst_r_sum1_4__5__q ),
	.datad(!Xd_0__inst_r_sum1_3__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_18 ),
	.sharein(Xd_0__inst_inst_add_2_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_21_sumout ),
	.cout(Xd_0__inst_inst_add_2_22 ),
	.shareout(Xd_0__inst_inst_add_2_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_22  = CARRY(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_23  = SHARE((!Xd_0__inst_r_sum1_2__5__q  & (Xd_0__inst_r_sum1_1__5__q  & Xd_0__inst_r_sum1_0__5__q )) # (Xd_0__inst_r_sum1_2__5__q  & ((Xd_0__inst_r_sum1_0__5__q ) # (Xd_0__inst_r_sum1_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__5__q ),
	.datad(!Xd_0__inst_r_sum1_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_25 (
// Equation(s):
// Xd_0__inst_inst_add_8_25_sumout  = SUM(( !Xd_0__inst_r_sum1_14__6__q  $ (!Xd_0__inst_r_sum1_13__6__q  $ (Xd_0__inst_r_sum1_12__6__q )) ) + ( Xd_0__inst_inst_add_8_23  ) + ( Xd_0__inst_inst_add_8_22  ))
// Xd_0__inst_inst_add_8_26  = CARRY(( !Xd_0__inst_r_sum1_14__6__q  $ (!Xd_0__inst_r_sum1_13__6__q  $ (Xd_0__inst_r_sum1_12__6__q )) ) + ( Xd_0__inst_inst_add_8_23  ) + ( Xd_0__inst_inst_add_8_22  ))
// Xd_0__inst_inst_add_8_27  = SHARE((!Xd_0__inst_r_sum1_14__6__q  & (Xd_0__inst_r_sum1_13__6__q  & Xd_0__inst_r_sum1_12__6__q )) # (Xd_0__inst_r_sum1_14__6__q  & ((Xd_0__inst_r_sum1_12__6__q ) # (Xd_0__inst_r_sum1_13__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__6__q ),
	.datac(!Xd_0__inst_r_sum1_13__6__q ),
	.datad(!Xd_0__inst_r_sum1_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_22 ),
	.sharein(Xd_0__inst_inst_add_8_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_25_sumout ),
	.cout(Xd_0__inst_inst_add_8_26 ),
	.shareout(Xd_0__inst_inst_add_8_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_25 (
// Equation(s):
// Xd_0__inst_inst_add_6_25_sumout  = SUM(( !Xd_0__inst_r_sum1_11__6__q  $ (!Xd_0__inst_r_sum1_10__6__q  $ (Xd_0__inst_r_sum1_9__6__q )) ) + ( Xd_0__inst_inst_add_6_23  ) + ( Xd_0__inst_inst_add_6_22  ))
// Xd_0__inst_inst_add_6_26  = CARRY(( !Xd_0__inst_r_sum1_11__6__q  $ (!Xd_0__inst_r_sum1_10__6__q  $ (Xd_0__inst_r_sum1_9__6__q )) ) + ( Xd_0__inst_inst_add_6_23  ) + ( Xd_0__inst_inst_add_6_22  ))
// Xd_0__inst_inst_add_6_27  = SHARE((!Xd_0__inst_r_sum1_11__6__q  & (Xd_0__inst_r_sum1_10__6__q  & Xd_0__inst_r_sum1_9__6__q )) # (Xd_0__inst_r_sum1_11__6__q  & ((Xd_0__inst_r_sum1_9__6__q ) # (Xd_0__inst_r_sum1_10__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__6__q ),
	.datac(!Xd_0__inst_r_sum1_10__6__q ),
	.datad(!Xd_0__inst_r_sum1_9__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_22 ),
	.sharein(Xd_0__inst_inst_add_6_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_25_sumout ),
	.cout(Xd_0__inst_inst_add_6_26 ),
	.shareout(Xd_0__inst_inst_add_6_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_25 (
// Equation(s):
// Xd_0__inst_inst_add_4_25_sumout  = SUM(( !Xd_0__inst_r_sum1_8__6__q  $ (!Xd_0__inst_r_sum1_7__6__q  $ (Xd_0__inst_r_sum1_6__6__q )) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_26  = CARRY(( !Xd_0__inst_r_sum1_8__6__q  $ (!Xd_0__inst_r_sum1_7__6__q  $ (Xd_0__inst_r_sum1_6__6__q )) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_27  = SHARE((!Xd_0__inst_r_sum1_8__6__q  & (Xd_0__inst_r_sum1_7__6__q  & Xd_0__inst_r_sum1_6__6__q )) # (Xd_0__inst_r_sum1_8__6__q  & ((Xd_0__inst_r_sum1_6__6__q ) # (Xd_0__inst_r_sum1_7__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__6__q ),
	.datac(!Xd_0__inst_r_sum1_7__6__q ),
	.datad(!Xd_0__inst_r_sum1_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_22 ),
	.sharein(Xd_0__inst_inst_add_4_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_25_sumout ),
	.cout(Xd_0__inst_inst_add_4_26 ),
	.shareout(Xd_0__inst_inst_add_4_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_25 (
// Equation(s):
// Xd_0__inst_inst_add_2_25_sumout  = SUM(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_26  = CARRY(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_27  = SHARE((!Xd_0__inst_r_sum1_5__6__q  & (Xd_0__inst_r_sum1_4__6__q  & Xd_0__inst_r_sum1_3__6__q )) # (Xd_0__inst_r_sum1_5__6__q  & ((Xd_0__inst_r_sum1_3__6__q ) # (Xd_0__inst_r_sum1_4__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__6__q ),
	.datac(!Xd_0__inst_r_sum1_4__6__q ),
	.datad(!Xd_0__inst_r_sum1_3__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_22 ),
	.sharein(Xd_0__inst_inst_add_2_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_25_sumout ),
	.cout(Xd_0__inst_inst_add_2_26 ),
	.shareout(Xd_0__inst_inst_add_2_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_26  = CARRY(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_27  = SHARE((!Xd_0__inst_r_sum1_2__6__q  & (Xd_0__inst_r_sum1_1__6__q  & Xd_0__inst_r_sum1_0__6__q )) # (Xd_0__inst_r_sum1_2__6__q  & ((Xd_0__inst_r_sum1_0__6__q ) # (Xd_0__inst_r_sum1_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__6__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_29 (
// Equation(s):
// Xd_0__inst_inst_add_8_29_sumout  = SUM(( !Xd_0__inst_r_sum1_14__7__q  $ (!Xd_0__inst_r_sum1_13__7__q  $ (Xd_0__inst_r_sum1_12__7__q )) ) + ( Xd_0__inst_inst_add_8_27  ) + ( Xd_0__inst_inst_add_8_26  ))
// Xd_0__inst_inst_add_8_30  = CARRY(( !Xd_0__inst_r_sum1_14__7__q  $ (!Xd_0__inst_r_sum1_13__7__q  $ (Xd_0__inst_r_sum1_12__7__q )) ) + ( Xd_0__inst_inst_add_8_27  ) + ( Xd_0__inst_inst_add_8_26  ))
// Xd_0__inst_inst_add_8_31  = SHARE((!Xd_0__inst_r_sum1_14__7__q  & (Xd_0__inst_r_sum1_13__7__q  & Xd_0__inst_r_sum1_12__7__q )) # (Xd_0__inst_r_sum1_14__7__q  & ((Xd_0__inst_r_sum1_12__7__q ) # (Xd_0__inst_r_sum1_13__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__7__q ),
	.datac(!Xd_0__inst_r_sum1_13__7__q ),
	.datad(!Xd_0__inst_r_sum1_12__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_26 ),
	.sharein(Xd_0__inst_inst_add_8_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_29_sumout ),
	.cout(Xd_0__inst_inst_add_8_30 ),
	.shareout(Xd_0__inst_inst_add_8_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_29 (
// Equation(s):
// Xd_0__inst_inst_add_6_29_sumout  = SUM(( !Xd_0__inst_r_sum1_11__7__q  $ (!Xd_0__inst_r_sum1_10__7__q  $ (Xd_0__inst_r_sum1_9__7__q )) ) + ( Xd_0__inst_inst_add_6_27  ) + ( Xd_0__inst_inst_add_6_26  ))
// Xd_0__inst_inst_add_6_30  = CARRY(( !Xd_0__inst_r_sum1_11__7__q  $ (!Xd_0__inst_r_sum1_10__7__q  $ (Xd_0__inst_r_sum1_9__7__q )) ) + ( Xd_0__inst_inst_add_6_27  ) + ( Xd_0__inst_inst_add_6_26  ))
// Xd_0__inst_inst_add_6_31  = SHARE((!Xd_0__inst_r_sum1_11__7__q  & (Xd_0__inst_r_sum1_10__7__q  & Xd_0__inst_r_sum1_9__7__q )) # (Xd_0__inst_r_sum1_11__7__q  & ((Xd_0__inst_r_sum1_9__7__q ) # (Xd_0__inst_r_sum1_10__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__7__q ),
	.datac(!Xd_0__inst_r_sum1_10__7__q ),
	.datad(!Xd_0__inst_r_sum1_9__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_26 ),
	.sharein(Xd_0__inst_inst_add_6_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_29_sumout ),
	.cout(Xd_0__inst_inst_add_6_30 ),
	.shareout(Xd_0__inst_inst_add_6_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_29 (
// Equation(s):
// Xd_0__inst_inst_add_4_29_sumout  = SUM(( !Xd_0__inst_r_sum1_8__7__q  $ (!Xd_0__inst_r_sum1_7__7__q  $ (Xd_0__inst_r_sum1_6__7__q )) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_30  = CARRY(( !Xd_0__inst_r_sum1_8__7__q  $ (!Xd_0__inst_r_sum1_7__7__q  $ (Xd_0__inst_r_sum1_6__7__q )) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_31  = SHARE((!Xd_0__inst_r_sum1_8__7__q  & (Xd_0__inst_r_sum1_7__7__q  & Xd_0__inst_r_sum1_6__7__q )) # (Xd_0__inst_r_sum1_8__7__q  & ((Xd_0__inst_r_sum1_6__7__q ) # (Xd_0__inst_r_sum1_7__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__7__q ),
	.datac(!Xd_0__inst_r_sum1_7__7__q ),
	.datad(!Xd_0__inst_r_sum1_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_26 ),
	.sharein(Xd_0__inst_inst_add_4_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_29_sumout ),
	.cout(Xd_0__inst_inst_add_4_30 ),
	.shareout(Xd_0__inst_inst_add_4_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_29 (
// Equation(s):
// Xd_0__inst_inst_add_2_29_sumout  = SUM(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_30  = CARRY(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_31  = SHARE((!Xd_0__inst_r_sum1_5__7__q  & (Xd_0__inst_r_sum1_4__7__q  & Xd_0__inst_r_sum1_3__7__q )) # (Xd_0__inst_r_sum1_5__7__q  & ((Xd_0__inst_r_sum1_3__7__q ) # (Xd_0__inst_r_sum1_4__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__7__q ),
	.datac(!Xd_0__inst_r_sum1_4__7__q ),
	.datad(!Xd_0__inst_r_sum1_3__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_26 ),
	.sharein(Xd_0__inst_inst_add_2_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_29_sumout ),
	.cout(Xd_0__inst_inst_add_2_30 ),
	.shareout(Xd_0__inst_inst_add_2_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_30  = CARRY(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_31  = SHARE((!Xd_0__inst_r_sum1_2__7__q  & (Xd_0__inst_r_sum1_1__7__q  & Xd_0__inst_r_sum1_0__7__q )) # (Xd_0__inst_r_sum1_2__7__q  & ((Xd_0__inst_r_sum1_0__7__q ) # (Xd_0__inst_r_sum1_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__7__q ),
	.datad(!Xd_0__inst_r_sum1_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_33 (
// Equation(s):
// Xd_0__inst_inst_add_8_33_sumout  = SUM(( !Xd_0__inst_r_sum1_14__8__q  $ (!Xd_0__inst_r_sum1_13__8__q  $ (Xd_0__inst_r_sum1_12__8__q )) ) + ( Xd_0__inst_inst_add_8_31  ) + ( Xd_0__inst_inst_add_8_30  ))
// Xd_0__inst_inst_add_8_34  = CARRY(( !Xd_0__inst_r_sum1_14__8__q  $ (!Xd_0__inst_r_sum1_13__8__q  $ (Xd_0__inst_r_sum1_12__8__q )) ) + ( Xd_0__inst_inst_add_8_31  ) + ( Xd_0__inst_inst_add_8_30  ))
// Xd_0__inst_inst_add_8_35  = SHARE((!Xd_0__inst_r_sum1_14__8__q  & (Xd_0__inst_r_sum1_13__8__q  & Xd_0__inst_r_sum1_12__8__q )) # (Xd_0__inst_r_sum1_14__8__q  & ((Xd_0__inst_r_sum1_12__8__q ) # (Xd_0__inst_r_sum1_13__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__8__q ),
	.datac(!Xd_0__inst_r_sum1_13__8__q ),
	.datad(!Xd_0__inst_r_sum1_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_30 ),
	.sharein(Xd_0__inst_inst_add_8_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_33_sumout ),
	.cout(Xd_0__inst_inst_add_8_34 ),
	.shareout(Xd_0__inst_inst_add_8_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_33 (
// Equation(s):
// Xd_0__inst_inst_add_6_33_sumout  = SUM(( !Xd_0__inst_r_sum1_11__8__q  $ (!Xd_0__inst_r_sum1_10__8__q  $ (Xd_0__inst_r_sum1_9__8__q )) ) + ( Xd_0__inst_inst_add_6_31  ) + ( Xd_0__inst_inst_add_6_30  ))
// Xd_0__inst_inst_add_6_34  = CARRY(( !Xd_0__inst_r_sum1_11__8__q  $ (!Xd_0__inst_r_sum1_10__8__q  $ (Xd_0__inst_r_sum1_9__8__q )) ) + ( Xd_0__inst_inst_add_6_31  ) + ( Xd_0__inst_inst_add_6_30  ))
// Xd_0__inst_inst_add_6_35  = SHARE((!Xd_0__inst_r_sum1_11__8__q  & (Xd_0__inst_r_sum1_10__8__q  & Xd_0__inst_r_sum1_9__8__q )) # (Xd_0__inst_r_sum1_11__8__q  & ((Xd_0__inst_r_sum1_9__8__q ) # (Xd_0__inst_r_sum1_10__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__8__q ),
	.datac(!Xd_0__inst_r_sum1_10__8__q ),
	.datad(!Xd_0__inst_r_sum1_9__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_30 ),
	.sharein(Xd_0__inst_inst_add_6_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_33_sumout ),
	.cout(Xd_0__inst_inst_add_6_34 ),
	.shareout(Xd_0__inst_inst_add_6_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_33 (
// Equation(s):
// Xd_0__inst_inst_add_4_33_sumout  = SUM(( !Xd_0__inst_r_sum1_8__8__q  $ (!Xd_0__inst_r_sum1_7__8__q  $ (Xd_0__inst_r_sum1_6__8__q )) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_34  = CARRY(( !Xd_0__inst_r_sum1_8__8__q  $ (!Xd_0__inst_r_sum1_7__8__q  $ (Xd_0__inst_r_sum1_6__8__q )) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_35  = SHARE((!Xd_0__inst_r_sum1_8__8__q  & (Xd_0__inst_r_sum1_7__8__q  & Xd_0__inst_r_sum1_6__8__q )) # (Xd_0__inst_r_sum1_8__8__q  & ((Xd_0__inst_r_sum1_6__8__q ) # (Xd_0__inst_r_sum1_7__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__8__q ),
	.datac(!Xd_0__inst_r_sum1_7__8__q ),
	.datad(!Xd_0__inst_r_sum1_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_30 ),
	.sharein(Xd_0__inst_inst_add_4_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_33_sumout ),
	.cout(Xd_0__inst_inst_add_4_34 ),
	.shareout(Xd_0__inst_inst_add_4_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_33 (
// Equation(s):
// Xd_0__inst_inst_add_2_33_sumout  = SUM(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_34  = CARRY(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_35  = SHARE((!Xd_0__inst_r_sum1_5__8__q  & (Xd_0__inst_r_sum1_4__8__q  & Xd_0__inst_r_sum1_3__8__q )) # (Xd_0__inst_r_sum1_5__8__q  & ((Xd_0__inst_r_sum1_3__8__q ) # (Xd_0__inst_r_sum1_4__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__8__q ),
	.datac(!Xd_0__inst_r_sum1_4__8__q ),
	.datad(!Xd_0__inst_r_sum1_3__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_30 ),
	.sharein(Xd_0__inst_inst_add_2_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_33_sumout ),
	.cout(Xd_0__inst_inst_add_2_34 ),
	.shareout(Xd_0__inst_inst_add_2_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_34  = CARRY(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_35  = SHARE((!Xd_0__inst_r_sum1_2__8__q  & (Xd_0__inst_r_sum1_1__8__q  & Xd_0__inst_r_sum1_0__8__q )) # (Xd_0__inst_r_sum1_2__8__q  & ((Xd_0__inst_r_sum1_0__8__q ) # (Xd_0__inst_r_sum1_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__8__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_37 (
// Equation(s):
// Xd_0__inst_inst_add_8_37_sumout  = SUM(( !Xd_0__inst_r_sum1_14__9__q  $ (!Xd_0__inst_r_sum1_13__9__q  $ (Xd_0__inst_r_sum1_12__9__q )) ) + ( Xd_0__inst_inst_add_8_35  ) + ( Xd_0__inst_inst_add_8_34  ))
// Xd_0__inst_inst_add_8_38  = CARRY(( !Xd_0__inst_r_sum1_14__9__q  $ (!Xd_0__inst_r_sum1_13__9__q  $ (Xd_0__inst_r_sum1_12__9__q )) ) + ( Xd_0__inst_inst_add_8_35  ) + ( Xd_0__inst_inst_add_8_34  ))
// Xd_0__inst_inst_add_8_39  = SHARE((!Xd_0__inst_r_sum1_14__9__q  & (Xd_0__inst_r_sum1_13__9__q  & Xd_0__inst_r_sum1_12__9__q )) # (Xd_0__inst_r_sum1_14__9__q  & ((Xd_0__inst_r_sum1_12__9__q ) # (Xd_0__inst_r_sum1_13__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__9__q ),
	.datac(!Xd_0__inst_r_sum1_13__9__q ),
	.datad(!Xd_0__inst_r_sum1_12__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_34 ),
	.sharein(Xd_0__inst_inst_add_8_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_37_sumout ),
	.cout(Xd_0__inst_inst_add_8_38 ),
	.shareout(Xd_0__inst_inst_add_8_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_37 (
// Equation(s):
// Xd_0__inst_inst_add_6_37_sumout  = SUM(( !Xd_0__inst_r_sum1_11__9__q  $ (!Xd_0__inst_r_sum1_10__9__q  $ (Xd_0__inst_r_sum1_9__9__q )) ) + ( Xd_0__inst_inst_add_6_35  ) + ( Xd_0__inst_inst_add_6_34  ))
// Xd_0__inst_inst_add_6_38  = CARRY(( !Xd_0__inst_r_sum1_11__9__q  $ (!Xd_0__inst_r_sum1_10__9__q  $ (Xd_0__inst_r_sum1_9__9__q )) ) + ( Xd_0__inst_inst_add_6_35  ) + ( Xd_0__inst_inst_add_6_34  ))
// Xd_0__inst_inst_add_6_39  = SHARE((!Xd_0__inst_r_sum1_11__9__q  & (Xd_0__inst_r_sum1_10__9__q  & Xd_0__inst_r_sum1_9__9__q )) # (Xd_0__inst_r_sum1_11__9__q  & ((Xd_0__inst_r_sum1_9__9__q ) # (Xd_0__inst_r_sum1_10__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__9__q ),
	.datac(!Xd_0__inst_r_sum1_10__9__q ),
	.datad(!Xd_0__inst_r_sum1_9__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_34 ),
	.sharein(Xd_0__inst_inst_add_6_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_37_sumout ),
	.cout(Xd_0__inst_inst_add_6_38 ),
	.shareout(Xd_0__inst_inst_add_6_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_37 (
// Equation(s):
// Xd_0__inst_inst_add_4_37_sumout  = SUM(( !Xd_0__inst_r_sum1_8__9__q  $ (!Xd_0__inst_r_sum1_7__9__q  $ (Xd_0__inst_r_sum1_6__9__q )) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_38  = CARRY(( !Xd_0__inst_r_sum1_8__9__q  $ (!Xd_0__inst_r_sum1_7__9__q  $ (Xd_0__inst_r_sum1_6__9__q )) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_39  = SHARE((!Xd_0__inst_r_sum1_8__9__q  & (Xd_0__inst_r_sum1_7__9__q  & Xd_0__inst_r_sum1_6__9__q )) # (Xd_0__inst_r_sum1_8__9__q  & ((Xd_0__inst_r_sum1_6__9__q ) # (Xd_0__inst_r_sum1_7__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__9__q ),
	.datac(!Xd_0__inst_r_sum1_7__9__q ),
	.datad(!Xd_0__inst_r_sum1_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_34 ),
	.sharein(Xd_0__inst_inst_add_4_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_37_sumout ),
	.cout(Xd_0__inst_inst_add_4_38 ),
	.shareout(Xd_0__inst_inst_add_4_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_37 (
// Equation(s):
// Xd_0__inst_inst_add_2_37_sumout  = SUM(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_38  = CARRY(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_39  = SHARE((!Xd_0__inst_r_sum1_5__9__q  & (Xd_0__inst_r_sum1_4__9__q  & Xd_0__inst_r_sum1_3__9__q )) # (Xd_0__inst_r_sum1_5__9__q  & ((Xd_0__inst_r_sum1_3__9__q ) # (Xd_0__inst_r_sum1_4__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__9__q ),
	.datac(!Xd_0__inst_r_sum1_4__9__q ),
	.datad(!Xd_0__inst_r_sum1_3__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_34 ),
	.sharein(Xd_0__inst_inst_add_2_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_37_sumout ),
	.cout(Xd_0__inst_inst_add_2_38 ),
	.shareout(Xd_0__inst_inst_add_2_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_38  = CARRY(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_39  = SHARE((!Xd_0__inst_r_sum1_2__9__q  & (Xd_0__inst_r_sum1_1__9__q  & Xd_0__inst_r_sum1_0__9__q )) # (Xd_0__inst_r_sum1_2__9__q  & ((Xd_0__inst_r_sum1_0__9__q ) # (Xd_0__inst_r_sum1_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__9__q ),
	.datad(!Xd_0__inst_r_sum1_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_41 (
// Equation(s):
// Xd_0__inst_inst_add_8_41_sumout  = SUM(( !Xd_0__inst_r_sum1_14__10__q  $ (!Xd_0__inst_r_sum1_13__10__q  $ (Xd_0__inst_r_sum1_12__10__q )) ) + ( Xd_0__inst_inst_add_8_39  ) + ( Xd_0__inst_inst_add_8_38  ))
// Xd_0__inst_inst_add_8_42  = CARRY(( !Xd_0__inst_r_sum1_14__10__q  $ (!Xd_0__inst_r_sum1_13__10__q  $ (Xd_0__inst_r_sum1_12__10__q )) ) + ( Xd_0__inst_inst_add_8_39  ) + ( Xd_0__inst_inst_add_8_38  ))
// Xd_0__inst_inst_add_8_43  = SHARE((!Xd_0__inst_r_sum1_14__10__q  & (Xd_0__inst_r_sum1_13__10__q  & Xd_0__inst_r_sum1_12__10__q )) # (Xd_0__inst_r_sum1_14__10__q  & ((Xd_0__inst_r_sum1_12__10__q ) # (Xd_0__inst_r_sum1_13__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__10__q ),
	.datac(!Xd_0__inst_r_sum1_13__10__q ),
	.datad(!Xd_0__inst_r_sum1_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_38 ),
	.sharein(Xd_0__inst_inst_add_8_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_41_sumout ),
	.cout(Xd_0__inst_inst_add_8_42 ),
	.shareout(Xd_0__inst_inst_add_8_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_41 (
// Equation(s):
// Xd_0__inst_inst_add_6_41_sumout  = SUM(( !Xd_0__inst_r_sum1_11__10__q  $ (!Xd_0__inst_r_sum1_10__10__q  $ (Xd_0__inst_r_sum1_9__10__q )) ) + ( Xd_0__inst_inst_add_6_39  ) + ( Xd_0__inst_inst_add_6_38  ))
// Xd_0__inst_inst_add_6_42  = CARRY(( !Xd_0__inst_r_sum1_11__10__q  $ (!Xd_0__inst_r_sum1_10__10__q  $ (Xd_0__inst_r_sum1_9__10__q )) ) + ( Xd_0__inst_inst_add_6_39  ) + ( Xd_0__inst_inst_add_6_38  ))
// Xd_0__inst_inst_add_6_43  = SHARE((!Xd_0__inst_r_sum1_11__10__q  & (Xd_0__inst_r_sum1_10__10__q  & Xd_0__inst_r_sum1_9__10__q )) # (Xd_0__inst_r_sum1_11__10__q  & ((Xd_0__inst_r_sum1_9__10__q ) # (Xd_0__inst_r_sum1_10__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__10__q ),
	.datac(!Xd_0__inst_r_sum1_10__10__q ),
	.datad(!Xd_0__inst_r_sum1_9__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_38 ),
	.sharein(Xd_0__inst_inst_add_6_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_41_sumout ),
	.cout(Xd_0__inst_inst_add_6_42 ),
	.shareout(Xd_0__inst_inst_add_6_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_41 (
// Equation(s):
// Xd_0__inst_inst_add_4_41_sumout  = SUM(( !Xd_0__inst_r_sum1_8__10__q  $ (!Xd_0__inst_r_sum1_7__10__q  $ (Xd_0__inst_r_sum1_6__10__q )) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_42  = CARRY(( !Xd_0__inst_r_sum1_8__10__q  $ (!Xd_0__inst_r_sum1_7__10__q  $ (Xd_0__inst_r_sum1_6__10__q )) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_43  = SHARE((!Xd_0__inst_r_sum1_8__10__q  & (Xd_0__inst_r_sum1_7__10__q  & Xd_0__inst_r_sum1_6__10__q )) # (Xd_0__inst_r_sum1_8__10__q  & ((Xd_0__inst_r_sum1_6__10__q ) # (Xd_0__inst_r_sum1_7__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__10__q ),
	.datac(!Xd_0__inst_r_sum1_7__10__q ),
	.datad(!Xd_0__inst_r_sum1_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_38 ),
	.sharein(Xd_0__inst_inst_add_4_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_41_sumout ),
	.cout(Xd_0__inst_inst_add_4_42 ),
	.shareout(Xd_0__inst_inst_add_4_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_41 (
// Equation(s):
// Xd_0__inst_inst_add_2_41_sumout  = SUM(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_42  = CARRY(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_43  = SHARE((!Xd_0__inst_r_sum1_5__10__q  & (Xd_0__inst_r_sum1_4__10__q  & Xd_0__inst_r_sum1_3__10__q )) # (Xd_0__inst_r_sum1_5__10__q  & ((Xd_0__inst_r_sum1_3__10__q ) # (Xd_0__inst_r_sum1_4__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__10__q ),
	.datac(!Xd_0__inst_r_sum1_4__10__q ),
	.datad(!Xd_0__inst_r_sum1_3__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_38 ),
	.sharein(Xd_0__inst_inst_add_2_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_41_sumout ),
	.cout(Xd_0__inst_inst_add_2_42 ),
	.shareout(Xd_0__inst_inst_add_2_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_42  = CARRY(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_43  = SHARE((!Xd_0__inst_r_sum1_2__10__q  & (Xd_0__inst_r_sum1_1__10__q  & Xd_0__inst_r_sum1_0__10__q )) # (Xd_0__inst_r_sum1_2__10__q  & ((Xd_0__inst_r_sum1_0__10__q ) # (Xd_0__inst_r_sum1_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__10__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_45 (
// Equation(s):
// Xd_0__inst_inst_add_8_45_sumout  = SUM(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_43  ) + ( Xd_0__inst_inst_add_8_42  ))
// Xd_0__inst_inst_add_8_46  = CARRY(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_43  ) + ( Xd_0__inst_inst_add_8_42  ))
// Xd_0__inst_inst_add_8_47  = SHARE((!Xd_0__inst_r_sum1_14__11__q  & (Xd_0__inst_r_sum1_13__11__q  & Xd_0__inst_r_sum1_12__11__q )) # (Xd_0__inst_r_sum1_14__11__q  & ((Xd_0__inst_r_sum1_12__11__q ) # (Xd_0__inst_r_sum1_13__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__11__q ),
	.datad(!Xd_0__inst_r_sum1_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_42 ),
	.sharein(Xd_0__inst_inst_add_8_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_45_sumout ),
	.cout(Xd_0__inst_inst_add_8_46 ),
	.shareout(Xd_0__inst_inst_add_8_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_45 (
// Equation(s):
// Xd_0__inst_inst_add_6_45_sumout  = SUM(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_43  ) + ( Xd_0__inst_inst_add_6_42  ))
// Xd_0__inst_inst_add_6_46  = CARRY(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_43  ) + ( Xd_0__inst_inst_add_6_42  ))
// Xd_0__inst_inst_add_6_47  = SHARE((!Xd_0__inst_r_sum1_11__11__q  & (Xd_0__inst_r_sum1_10__11__q  & Xd_0__inst_r_sum1_9__11__q )) # (Xd_0__inst_r_sum1_11__11__q  & ((Xd_0__inst_r_sum1_9__11__q ) # (Xd_0__inst_r_sum1_10__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__11__q ),
	.datad(!Xd_0__inst_r_sum1_9__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_42 ),
	.sharein(Xd_0__inst_inst_add_6_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_45_sumout ),
	.cout(Xd_0__inst_inst_add_6_46 ),
	.shareout(Xd_0__inst_inst_add_6_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_45 (
// Equation(s):
// Xd_0__inst_inst_add_4_45_sumout  = SUM(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_46  = CARRY(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_47  = SHARE((!Xd_0__inst_r_sum1_8__11__q  & (Xd_0__inst_r_sum1_7__11__q  & Xd_0__inst_r_sum1_6__11__q )) # (Xd_0__inst_r_sum1_8__11__q  & ((Xd_0__inst_r_sum1_6__11__q ) # (Xd_0__inst_r_sum1_7__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__11__q ),
	.datad(!Xd_0__inst_r_sum1_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_42 ),
	.sharein(Xd_0__inst_inst_add_4_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_45_sumout ),
	.cout(Xd_0__inst_inst_add_4_46 ),
	.shareout(Xd_0__inst_inst_add_4_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_45 (
// Equation(s):
// Xd_0__inst_inst_add_2_45_sumout  = SUM(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_46  = CARRY(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_47  = SHARE((!Xd_0__inst_r_sum1_5__11__q  & (Xd_0__inst_r_sum1_4__11__q  & Xd_0__inst_r_sum1_3__11__q )) # (Xd_0__inst_r_sum1_5__11__q  & ((Xd_0__inst_r_sum1_3__11__q ) # (Xd_0__inst_r_sum1_4__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__11__q ),
	.datad(!Xd_0__inst_r_sum1_3__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_42 ),
	.sharein(Xd_0__inst_inst_add_2_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_45_sumout ),
	.cout(Xd_0__inst_inst_add_2_46 ),
	.shareout(Xd_0__inst_inst_add_2_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_46  = CARRY(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_47  = SHARE((!Xd_0__inst_r_sum1_2__11__q  & (Xd_0__inst_r_sum1_1__11__q  & Xd_0__inst_r_sum1_0__11__q )) # (Xd_0__inst_r_sum1_2__11__q  & ((Xd_0__inst_r_sum1_0__11__q ) # (Xd_0__inst_r_sum1_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_49 (
// Equation(s):
// Xd_0__inst_inst_add_8_49_sumout  = SUM(( !Xd_0__inst_r_sum1_14__12__q  $ (!Xd_0__inst_r_sum1_13__12__q  $ (Xd_0__inst_r_sum1_12__12__q )) ) + ( Xd_0__inst_inst_add_8_47  ) + ( Xd_0__inst_inst_add_8_46  ))
// Xd_0__inst_inst_add_8_50  = CARRY(( !Xd_0__inst_r_sum1_14__12__q  $ (!Xd_0__inst_r_sum1_13__12__q  $ (Xd_0__inst_r_sum1_12__12__q )) ) + ( Xd_0__inst_inst_add_8_47  ) + ( Xd_0__inst_inst_add_8_46  ))
// Xd_0__inst_inst_add_8_51  = SHARE((!Xd_0__inst_r_sum1_14__12__q  & (Xd_0__inst_r_sum1_13__12__q  & Xd_0__inst_r_sum1_12__12__q )) # (Xd_0__inst_r_sum1_14__12__q  & ((Xd_0__inst_r_sum1_12__12__q ) # (Xd_0__inst_r_sum1_13__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__12__q ),
	.datac(!Xd_0__inst_r_sum1_13__12__q ),
	.datad(!Xd_0__inst_r_sum1_12__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_46 ),
	.sharein(Xd_0__inst_inst_add_8_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_49_sumout ),
	.cout(Xd_0__inst_inst_add_8_50 ),
	.shareout(Xd_0__inst_inst_add_8_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_49 (
// Equation(s):
// Xd_0__inst_inst_add_6_49_sumout  = SUM(( !Xd_0__inst_r_sum1_11__12__q  $ (!Xd_0__inst_r_sum1_10__12__q  $ (Xd_0__inst_r_sum1_9__12__q )) ) + ( Xd_0__inst_inst_add_6_47  ) + ( Xd_0__inst_inst_add_6_46  ))
// Xd_0__inst_inst_add_6_50  = CARRY(( !Xd_0__inst_r_sum1_11__12__q  $ (!Xd_0__inst_r_sum1_10__12__q  $ (Xd_0__inst_r_sum1_9__12__q )) ) + ( Xd_0__inst_inst_add_6_47  ) + ( Xd_0__inst_inst_add_6_46  ))
// Xd_0__inst_inst_add_6_51  = SHARE((!Xd_0__inst_r_sum1_11__12__q  & (Xd_0__inst_r_sum1_10__12__q  & Xd_0__inst_r_sum1_9__12__q )) # (Xd_0__inst_r_sum1_11__12__q  & ((Xd_0__inst_r_sum1_9__12__q ) # (Xd_0__inst_r_sum1_10__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__12__q ),
	.datac(!Xd_0__inst_r_sum1_10__12__q ),
	.datad(!Xd_0__inst_r_sum1_9__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_46 ),
	.sharein(Xd_0__inst_inst_add_6_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_49_sumout ),
	.cout(Xd_0__inst_inst_add_6_50 ),
	.shareout(Xd_0__inst_inst_add_6_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_49 (
// Equation(s):
// Xd_0__inst_inst_add_4_49_sumout  = SUM(( !Xd_0__inst_r_sum1_8__12__q  $ (!Xd_0__inst_r_sum1_7__12__q  $ (Xd_0__inst_r_sum1_6__12__q )) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_50  = CARRY(( !Xd_0__inst_r_sum1_8__12__q  $ (!Xd_0__inst_r_sum1_7__12__q  $ (Xd_0__inst_r_sum1_6__12__q )) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_51  = SHARE((!Xd_0__inst_r_sum1_8__12__q  & (Xd_0__inst_r_sum1_7__12__q  & Xd_0__inst_r_sum1_6__12__q )) # (Xd_0__inst_r_sum1_8__12__q  & ((Xd_0__inst_r_sum1_6__12__q ) # (Xd_0__inst_r_sum1_7__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__12__q ),
	.datac(!Xd_0__inst_r_sum1_7__12__q ),
	.datad(!Xd_0__inst_r_sum1_6__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_46 ),
	.sharein(Xd_0__inst_inst_add_4_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_49_sumout ),
	.cout(Xd_0__inst_inst_add_4_50 ),
	.shareout(Xd_0__inst_inst_add_4_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_49 (
// Equation(s):
// Xd_0__inst_inst_add_2_49_sumout  = SUM(( !Xd_0__inst_r_sum1_5__12__q  $ (!Xd_0__inst_r_sum1_4__12__q  $ (Xd_0__inst_r_sum1_3__12__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_50  = CARRY(( !Xd_0__inst_r_sum1_5__12__q  $ (!Xd_0__inst_r_sum1_4__12__q  $ (Xd_0__inst_r_sum1_3__12__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_51  = SHARE((!Xd_0__inst_r_sum1_5__12__q  & (Xd_0__inst_r_sum1_4__12__q  & Xd_0__inst_r_sum1_3__12__q )) # (Xd_0__inst_r_sum1_5__12__q  & ((Xd_0__inst_r_sum1_3__12__q ) # (Xd_0__inst_r_sum1_4__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__12__q ),
	.datac(!Xd_0__inst_r_sum1_4__12__q ),
	.datad(!Xd_0__inst_r_sum1_3__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_46 ),
	.sharein(Xd_0__inst_inst_add_2_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_49_sumout ),
	.cout(Xd_0__inst_inst_add_2_50 ),
	.shareout(Xd_0__inst_inst_add_2_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_50  = CARRY(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_51  = SHARE((!Xd_0__inst_r_sum1_2__12__q  & (Xd_0__inst_r_sum1_1__12__q  & Xd_0__inst_r_sum1_0__12__q )) # (Xd_0__inst_r_sum1_2__12__q  & ((Xd_0__inst_r_sum1_0__12__q ) # (Xd_0__inst_r_sum1_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__12__q ),
	.datac(!Xd_0__inst_r_sum1_1__12__q ),
	.datad(!Xd_0__inst_r_sum1_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_53 (
// Equation(s):
// Xd_0__inst_inst_add_8_53_sumout  = SUM(( !Xd_0__inst_r_sum1_14__13__q  $ (!Xd_0__inst_r_sum1_13__13__q  $ (Xd_0__inst_r_sum1_12__13__q )) ) + ( Xd_0__inst_inst_add_8_51  ) + ( Xd_0__inst_inst_add_8_50  ))
// Xd_0__inst_inst_add_8_54  = CARRY(( !Xd_0__inst_r_sum1_14__13__q  $ (!Xd_0__inst_r_sum1_13__13__q  $ (Xd_0__inst_r_sum1_12__13__q )) ) + ( Xd_0__inst_inst_add_8_51  ) + ( Xd_0__inst_inst_add_8_50  ))
// Xd_0__inst_inst_add_8_55  = SHARE((!Xd_0__inst_r_sum1_14__13__q  & (Xd_0__inst_r_sum1_13__13__q  & Xd_0__inst_r_sum1_12__13__q )) # (Xd_0__inst_r_sum1_14__13__q  & ((Xd_0__inst_r_sum1_12__13__q ) # (Xd_0__inst_r_sum1_13__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__13__q ),
	.datac(!Xd_0__inst_r_sum1_13__13__q ),
	.datad(!Xd_0__inst_r_sum1_12__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_50 ),
	.sharein(Xd_0__inst_inst_add_8_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_53_sumout ),
	.cout(Xd_0__inst_inst_add_8_54 ),
	.shareout(Xd_0__inst_inst_add_8_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_53 (
// Equation(s):
// Xd_0__inst_inst_add_6_53_sumout  = SUM(( !Xd_0__inst_r_sum1_11__13__q  $ (!Xd_0__inst_r_sum1_10__13__q  $ (Xd_0__inst_r_sum1_9__13__q )) ) + ( Xd_0__inst_inst_add_6_51  ) + ( Xd_0__inst_inst_add_6_50  ))
// Xd_0__inst_inst_add_6_54  = CARRY(( !Xd_0__inst_r_sum1_11__13__q  $ (!Xd_0__inst_r_sum1_10__13__q  $ (Xd_0__inst_r_sum1_9__13__q )) ) + ( Xd_0__inst_inst_add_6_51  ) + ( Xd_0__inst_inst_add_6_50  ))
// Xd_0__inst_inst_add_6_55  = SHARE((!Xd_0__inst_r_sum1_11__13__q  & (Xd_0__inst_r_sum1_10__13__q  & Xd_0__inst_r_sum1_9__13__q )) # (Xd_0__inst_r_sum1_11__13__q  & ((Xd_0__inst_r_sum1_9__13__q ) # (Xd_0__inst_r_sum1_10__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__13__q ),
	.datac(!Xd_0__inst_r_sum1_10__13__q ),
	.datad(!Xd_0__inst_r_sum1_9__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_50 ),
	.sharein(Xd_0__inst_inst_add_6_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_53_sumout ),
	.cout(Xd_0__inst_inst_add_6_54 ),
	.shareout(Xd_0__inst_inst_add_6_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_53 (
// Equation(s):
// Xd_0__inst_inst_add_4_53_sumout  = SUM(( !Xd_0__inst_r_sum1_8__13__q  $ (!Xd_0__inst_r_sum1_7__13__q  $ (Xd_0__inst_r_sum1_6__13__q )) ) + ( Xd_0__inst_inst_add_4_51  ) + ( Xd_0__inst_inst_add_4_50  ))
// Xd_0__inst_inst_add_4_54  = CARRY(( !Xd_0__inst_r_sum1_8__13__q  $ (!Xd_0__inst_r_sum1_7__13__q  $ (Xd_0__inst_r_sum1_6__13__q )) ) + ( Xd_0__inst_inst_add_4_51  ) + ( Xd_0__inst_inst_add_4_50  ))
// Xd_0__inst_inst_add_4_55  = SHARE((!Xd_0__inst_r_sum1_8__13__q  & (Xd_0__inst_r_sum1_7__13__q  & Xd_0__inst_r_sum1_6__13__q )) # (Xd_0__inst_r_sum1_8__13__q  & ((Xd_0__inst_r_sum1_6__13__q ) # (Xd_0__inst_r_sum1_7__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__13__q ),
	.datac(!Xd_0__inst_r_sum1_7__13__q ),
	.datad(!Xd_0__inst_r_sum1_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_50 ),
	.sharein(Xd_0__inst_inst_add_4_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_53_sumout ),
	.cout(Xd_0__inst_inst_add_4_54 ),
	.shareout(Xd_0__inst_inst_add_4_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_53 (
// Equation(s):
// Xd_0__inst_inst_add_2_53_sumout  = SUM(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_51  ) + ( Xd_0__inst_inst_add_2_50  ))
// Xd_0__inst_inst_add_2_54  = CARRY(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_51  ) + ( Xd_0__inst_inst_add_2_50  ))
// Xd_0__inst_inst_add_2_55  = SHARE((!Xd_0__inst_r_sum1_5__13__q  & (Xd_0__inst_r_sum1_4__13__q  & Xd_0__inst_r_sum1_3__13__q )) # (Xd_0__inst_r_sum1_5__13__q  & ((Xd_0__inst_r_sum1_3__13__q ) # (Xd_0__inst_r_sum1_4__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__13__q ),
	.datad(!Xd_0__inst_r_sum1_3__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_50 ),
	.sharein(Xd_0__inst_inst_add_2_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_53_sumout ),
	.cout(Xd_0__inst_inst_add_2_54 ),
	.shareout(Xd_0__inst_inst_add_2_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_54  = CARRY(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_55  = SHARE((!Xd_0__inst_r_sum1_2__13__q  & (Xd_0__inst_r_sum1_1__13__q  & Xd_0__inst_r_sum1_0__13__q )) # (Xd_0__inst_r_sum1_2__13__q  & ((Xd_0__inst_r_sum1_0__13__q ) # (Xd_0__inst_r_sum1_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__13__q ),
	.datad(!Xd_0__inst_r_sum1_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_57 (
// Equation(s):
// Xd_0__inst_inst_add_8_57_sumout  = SUM(( !Xd_0__inst_r_sum1_14__13__q  $ (!Xd_0__inst_r_sum1_13__13__q  $ (Xd_0__inst_r_sum1_12__13__q )) ) + ( Xd_0__inst_inst_add_8_55  ) + ( Xd_0__inst_inst_add_8_54  ))
// Xd_0__inst_inst_add_8_58  = CARRY(( !Xd_0__inst_r_sum1_14__13__q  $ (!Xd_0__inst_r_sum1_13__13__q  $ (Xd_0__inst_r_sum1_12__13__q )) ) + ( Xd_0__inst_inst_add_8_55  ) + ( Xd_0__inst_inst_add_8_54  ))
// Xd_0__inst_inst_add_8_59  = SHARE((!Xd_0__inst_r_sum1_14__13__q  & (Xd_0__inst_r_sum1_13__13__q  & Xd_0__inst_r_sum1_12__13__q )) # (Xd_0__inst_r_sum1_14__13__q  & ((Xd_0__inst_r_sum1_12__13__q ) # (Xd_0__inst_r_sum1_13__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__13__q ),
	.datac(!Xd_0__inst_r_sum1_13__13__q ),
	.datad(!Xd_0__inst_r_sum1_12__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_54 ),
	.sharein(Xd_0__inst_inst_add_8_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_57_sumout ),
	.cout(Xd_0__inst_inst_add_8_58 ),
	.shareout(Xd_0__inst_inst_add_8_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_57 (
// Equation(s):
// Xd_0__inst_inst_add_6_57_sumout  = SUM(( !Xd_0__inst_r_sum1_11__13__q  $ (!Xd_0__inst_r_sum1_10__13__q  $ (Xd_0__inst_r_sum1_9__13__q )) ) + ( Xd_0__inst_inst_add_6_55  ) + ( Xd_0__inst_inst_add_6_54  ))
// Xd_0__inst_inst_add_6_58  = CARRY(( !Xd_0__inst_r_sum1_11__13__q  $ (!Xd_0__inst_r_sum1_10__13__q  $ (Xd_0__inst_r_sum1_9__13__q )) ) + ( Xd_0__inst_inst_add_6_55  ) + ( Xd_0__inst_inst_add_6_54  ))
// Xd_0__inst_inst_add_6_59  = SHARE((!Xd_0__inst_r_sum1_11__13__q  & (Xd_0__inst_r_sum1_10__13__q  & Xd_0__inst_r_sum1_9__13__q )) # (Xd_0__inst_r_sum1_11__13__q  & ((Xd_0__inst_r_sum1_9__13__q ) # (Xd_0__inst_r_sum1_10__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__13__q ),
	.datac(!Xd_0__inst_r_sum1_10__13__q ),
	.datad(!Xd_0__inst_r_sum1_9__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_54 ),
	.sharein(Xd_0__inst_inst_add_6_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_57_sumout ),
	.cout(Xd_0__inst_inst_add_6_58 ),
	.shareout(Xd_0__inst_inst_add_6_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_57 (
// Equation(s):
// Xd_0__inst_inst_add_4_57_sumout  = SUM(( !Xd_0__inst_r_sum1_8__13__q  $ (!Xd_0__inst_r_sum1_7__13__q  $ (Xd_0__inst_r_sum1_6__13__q )) ) + ( Xd_0__inst_inst_add_4_55  ) + ( Xd_0__inst_inst_add_4_54  ))
// Xd_0__inst_inst_add_4_58  = CARRY(( !Xd_0__inst_r_sum1_8__13__q  $ (!Xd_0__inst_r_sum1_7__13__q  $ (Xd_0__inst_r_sum1_6__13__q )) ) + ( Xd_0__inst_inst_add_4_55  ) + ( Xd_0__inst_inst_add_4_54  ))
// Xd_0__inst_inst_add_4_59  = SHARE((!Xd_0__inst_r_sum1_8__13__q  & (Xd_0__inst_r_sum1_7__13__q  & Xd_0__inst_r_sum1_6__13__q )) # (Xd_0__inst_r_sum1_8__13__q  & ((Xd_0__inst_r_sum1_6__13__q ) # (Xd_0__inst_r_sum1_7__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__13__q ),
	.datac(!Xd_0__inst_r_sum1_7__13__q ),
	.datad(!Xd_0__inst_r_sum1_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_54 ),
	.sharein(Xd_0__inst_inst_add_4_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_57_sumout ),
	.cout(Xd_0__inst_inst_add_4_58 ),
	.shareout(Xd_0__inst_inst_add_4_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_57 (
// Equation(s):
// Xd_0__inst_inst_add_2_57_sumout  = SUM(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_55  ) + ( Xd_0__inst_inst_add_2_54  ))
// Xd_0__inst_inst_add_2_58  = CARRY(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_55  ) + ( Xd_0__inst_inst_add_2_54  ))
// Xd_0__inst_inst_add_2_59  = SHARE((!Xd_0__inst_r_sum1_5__13__q  & (Xd_0__inst_r_sum1_4__13__q  & Xd_0__inst_r_sum1_3__13__q )) # (Xd_0__inst_r_sum1_5__13__q  & ((Xd_0__inst_r_sum1_3__13__q ) # (Xd_0__inst_r_sum1_4__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__13__q ),
	.datad(!Xd_0__inst_r_sum1_3__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_54 ),
	.sharein(Xd_0__inst_inst_add_2_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_57_sumout ),
	.cout(Xd_0__inst_inst_add_2_58 ),
	.shareout(Xd_0__inst_inst_add_2_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_58  = CARRY(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_59  = SHARE((!Xd_0__inst_r_sum1_2__13__q  & (Xd_0__inst_r_sum1_1__13__q  & Xd_0__inst_r_sum1_0__13__q )) # (Xd_0__inst_r_sum1_2__13__q  & ((Xd_0__inst_r_sum1_0__13__q ) # (Xd_0__inst_r_sum1_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__13__q ),
	.datad(!Xd_0__inst_r_sum1_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_61 (
// Equation(s):
// Xd_0__inst_inst_add_8_61_sumout  = SUM(( !Xd_0__inst_r_sum1_14__13__q  $ (!Xd_0__inst_r_sum1_13__13__q  $ (Xd_0__inst_r_sum1_12__13__q )) ) + ( Xd_0__inst_inst_add_8_59  ) + ( Xd_0__inst_inst_add_8_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__13__q ),
	.datac(!Xd_0__inst_r_sum1_13__13__q ),
	.datad(!Xd_0__inst_r_sum1_12__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_58 ),
	.sharein(Xd_0__inst_inst_add_8_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_61 (
// Equation(s):
// Xd_0__inst_inst_add_6_61_sumout  = SUM(( !Xd_0__inst_r_sum1_11__13__q  $ (!Xd_0__inst_r_sum1_10__13__q  $ (Xd_0__inst_r_sum1_9__13__q )) ) + ( Xd_0__inst_inst_add_6_59  ) + ( Xd_0__inst_inst_add_6_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__13__q ),
	.datac(!Xd_0__inst_r_sum1_10__13__q ),
	.datad(!Xd_0__inst_r_sum1_9__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_58 ),
	.sharein(Xd_0__inst_inst_add_6_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_61 (
// Equation(s):
// Xd_0__inst_inst_add_4_61_sumout  = SUM(( !Xd_0__inst_r_sum1_8__13__q  $ (!Xd_0__inst_r_sum1_7__13__q  $ (Xd_0__inst_r_sum1_6__13__q )) ) + ( Xd_0__inst_inst_add_4_59  ) + ( Xd_0__inst_inst_add_4_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__13__q ),
	.datac(!Xd_0__inst_r_sum1_7__13__q ),
	.datad(!Xd_0__inst_r_sum1_6__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_58 ),
	.sharein(Xd_0__inst_inst_add_4_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_61 (
// Equation(s):
// Xd_0__inst_inst_add_2_61_sumout  = SUM(( !Xd_0__inst_r_sum1_5__13__q  $ (!Xd_0__inst_r_sum1_4__13__q  $ (Xd_0__inst_r_sum1_3__13__q )) ) + ( Xd_0__inst_inst_add_2_59  ) + ( Xd_0__inst_inst_add_2_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__13__q ),
	.datac(!Xd_0__inst_r_sum1_4__13__q ),
	.datad(!Xd_0__inst_r_sum1_3__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_58 ),
	.sharein(Xd_0__inst_inst_add_2_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_59  ) + ( Xd_0__inst_inst_add_0_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__13__q ),
	.datad(!Xd_0__inst_r_sum1_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_21 (
// Equation(s):
// Xd_0__inst_i19_21_sumout  = SUM(( !din_a[188] $ (!din_b[188]) ) + ( Xd_0__inst_i19_43  ) + ( Xd_0__inst_i19_42  ))
// Xd_0__inst_i19_22  = CARRY(( !din_a[188] $ (!din_b[188]) ) + ( Xd_0__inst_i19_43  ) + ( Xd_0__inst_i19_42  ))
// Xd_0__inst_i19_23  = SHARE(GND)

	.dataa(!din_a[188]),
	.datab(!din_b[188]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_42 ),
	.sharein(Xd_0__inst_i19_43 ),
	.combout(),
	.sumout(Xd_0__inst_i19_21_sumout ),
	.cout(Xd_0__inst_i19_22 ),
	.shareout(Xd_0__inst_i19_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_25 (
// Equation(s):
// Xd_0__inst_i19_25_sumout  = SUM(( !din_a[160] $ (!din_b[160]) ) + ( Xd_0__inst_i19_47  ) + ( Xd_0__inst_i19_46  ))
// Xd_0__inst_i19_26  = CARRY(( !din_a[160] $ (!din_b[160]) ) + ( Xd_0__inst_i19_47  ) + ( Xd_0__inst_i19_46  ))
// Xd_0__inst_i19_27  = SHARE(GND)

	.dataa(!din_a[160]),
	.datab(!din_b[160]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_46 ),
	.sharein(Xd_0__inst_i19_47 ),
	.combout(),
	.sumout(Xd_0__inst_i19_25_sumout ),
	.cout(Xd_0__inst_i19_26 ),
	.shareout(Xd_0__inst_i19_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_30__0__q  $ (!Xd_0__inst_product_31__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_30__0__q  $ (!Xd_0__inst_product_31__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_30__0__q  & ((!Xd_0__inst_sign [31] & ((Xd_0__inst_sign [30]))) # (Xd_0__inst_sign [31] & (!Xd_0__inst_product_31__0__q )))) # (Xd_0__inst_product_30__0__q  & ((!Xd_0__inst_sign [31] 
// & (Xd_0__inst_product_31__0__q )) # (Xd_0__inst_sign [31] & ((!Xd_0__inst_sign [30]))))))

	.dataa(!Xd_0__inst_product_30__0__q ),
	.datab(!Xd_0__inst_product_31__0__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_29 (
// Equation(s):
// Xd_0__inst_i19_29_sumout  = SUM(( !din_a[132] $ (!din_b[132]) ) + ( Xd_0__inst_i19_51  ) + ( Xd_0__inst_i19_50  ))
// Xd_0__inst_i19_30  = CARRY(( !din_a[132] $ (!din_b[132]) ) + ( Xd_0__inst_i19_51  ) + ( Xd_0__inst_i19_50  ))
// Xd_0__inst_i19_31  = SHARE(GND)

	.dataa(!din_a[132]),
	.datab(!din_b[132]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_50 ),
	.sharein(Xd_0__inst_i19_51 ),
	.combout(),
	.sumout(Xd_0__inst_i19_29_sumout ),
	.cout(Xd_0__inst_i19_30 ),
	.shareout(Xd_0__inst_i19_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_33 (
// Equation(s):
// Xd_0__inst_i19_33_sumout  = SUM(( !din_a[104] $ (!din_b[104]) ) + ( Xd_0__inst_i19_55  ) + ( Xd_0__inst_i19_54  ))
// Xd_0__inst_i19_34  = CARRY(( !din_a[104] $ (!din_b[104]) ) + ( Xd_0__inst_i19_55  ) + ( Xd_0__inst_i19_54  ))
// Xd_0__inst_i19_35  = SHARE(GND)

	.dataa(!din_a[104]),
	.datab(!din_b[104]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_54 ),
	.sharein(Xd_0__inst_i19_55 ),
	.combout(),
	.sumout(Xd_0__inst_i19_33_sumout ),
	.cout(Xd_0__inst_i19_34 ),
	.shareout(Xd_0__inst_i19_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_37 (
// Equation(s):
// Xd_0__inst_i19_37_sumout  = SUM(( !din_a[76] $ (!din_b[76]) ) + ( Xd_0__inst_i19_59  ) + ( Xd_0__inst_i19_58  ))
// Xd_0__inst_i19_38  = CARRY(( !din_a[76] $ (!din_b[76]) ) + ( Xd_0__inst_i19_59  ) + ( Xd_0__inst_i19_58  ))
// Xd_0__inst_i19_39  = SHARE(GND)

	.dataa(!din_a[76]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_58 ),
	.sharein(Xd_0__inst_i19_59 ),
	.combout(),
	.sumout(Xd_0__inst_i19_37_sumout ),
	.cout(Xd_0__inst_i19_38 ),
	.shareout(Xd_0__inst_i19_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_30__1__q  $ (!Xd_0__inst_product_31__1__q  $ (((Xd_0__inst_sign [31]) # (Xd_0__inst_sign [30])))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_30__1__q  $ (!Xd_0__inst_product_31__1__q  $ (((Xd_0__inst_sign [31]) # (Xd_0__inst_sign [30])))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [30] & (Xd_0__inst_product_30__1__q  & (!Xd_0__inst_product_31__1__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_sign [30] & ((!Xd_0__inst_product_31__1__q  & ((Xd_0__inst_sign [31]))) 
// # (Xd_0__inst_product_31__1__q  & (!Xd_0__inst_product_30__1__q )))))

	.dataa(!Xd_0__inst_product_30__1__q ),
	.datab(!Xd_0__inst_product_31__1__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_30__2__q  $ (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_30__2__q  $ (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__2__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__2__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__2__q ),
	.datab(!Xd_0__inst_product_31__2__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_30__3__q  $ (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_30__3__q  $ (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__3__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__3__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__3__q ),
	.datab(!Xd_0__inst_product_31__3__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_30__4__q  $ (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_30__4__q  $ (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__4__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__4__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__4__q ),
	.datab(!Xd_0__inst_product_31__4__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_30__5__q  $ (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_30__5__q  $ (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__5__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__5__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__5__q ),
	.datab(!Xd_0__inst_product_31__5__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_30__6__q  $ (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_30__6__q  $ (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__6__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__6__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__6__q ),
	.datab(!Xd_0__inst_product_31__6__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_30__7__q  $ (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_30__7__q  $ (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__7__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__7__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__7__q ),
	.datab(!Xd_0__inst_product_31__7__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_30__8__q  $ (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_30__8__q  $ (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__8__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__8__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__8__q ),
	.datab(!Xd_0__inst_product_31__8__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_30__9__q  $ (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_30__9__q  $ (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__9__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__9__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__9__q ),
	.datab(!Xd_0__inst_product_31__9__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_30__10__q  $ (!Xd_0__inst_product_31__10__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_30__10__q  $ (!Xd_0__inst_product_31__10__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__10__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__10__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__10__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__10__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__10__q ),
	.datab(!Xd_0__inst_product_31__10__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_30__11__q  $ (!Xd_0__inst_product_31__11__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_30__11__q  $ (!Xd_0__inst_product_31__11__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__11__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__11__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__11__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__11__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__11__q ),
	.datab(!Xd_0__inst_product_31__11__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [30] & Xd_0__inst_sign [31]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_28__0__q  $ (!Xd_0__inst_product_29__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_28__0__q  $ (!Xd_0__inst_product_29__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_28__0__q  & ((!Xd_0__inst_sign [29] & ((Xd_0__inst_sign [28]))) # (Xd_0__inst_sign [29] & (!Xd_0__inst_product_29__0__q )))) # (Xd_0__inst_product_28__0__q  & ((!Xd_0__inst_sign [29] 
// & (Xd_0__inst_product_29__0__q )) # (Xd_0__inst_sign [29] & ((!Xd_0__inst_sign [28]))))))

	.dataa(!Xd_0__inst_product_28__0__q ),
	.datab(!Xd_0__inst_product_29__0__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_26__0__q  $ (!Xd_0__inst_product_27__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_26__0__q  $ (!Xd_0__inst_product_27__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_26__0__q  & ((!Xd_0__inst_sign [27] & ((Xd_0__inst_sign [26]))) # (Xd_0__inst_sign [27] & (!Xd_0__inst_product_27__0__q )))) # (Xd_0__inst_product_26__0__q  & ((!Xd_0__inst_sign [27] 
// & (Xd_0__inst_product_27__0__q )) # (Xd_0__inst_sign [27] & ((!Xd_0__inst_sign [26]))))))

	.dataa(!Xd_0__inst_product_26__0__q ),
	.datab(!Xd_0__inst_product_27__0__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_24__0__q  $ (!Xd_0__inst_product_25__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_24__0__q  $ (!Xd_0__inst_product_25__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_24__0__q  & ((!Xd_0__inst_sign [25] & ((Xd_0__inst_sign [24]))) # (Xd_0__inst_sign [25] & (!Xd_0__inst_product_25__0__q )))) # (Xd_0__inst_product_24__0__q  & ((!Xd_0__inst_sign [25] 
// & (Xd_0__inst_product_25__0__q )) # (Xd_0__inst_sign [25] & ((!Xd_0__inst_sign [24]))))))

	.dataa(!Xd_0__inst_product_24__0__q ),
	.datab(!Xd_0__inst_product_25__0__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_41 (
// Equation(s):
// Xd_0__inst_i19_41_sumout  = SUM(( !din_a[195] $ (!din_b[195]) ) + ( Xd_0__inst_i19_63  ) + ( Xd_0__inst_i19_62  ))
// Xd_0__inst_i19_42  = CARRY(( !din_a[195] $ (!din_b[195]) ) + ( Xd_0__inst_i19_63  ) + ( Xd_0__inst_i19_62  ))
// Xd_0__inst_i19_43  = SHARE(GND)

	.dataa(!din_a[195]),
	.datab(!din_b[195]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_62 ),
	.sharein(Xd_0__inst_i19_63 ),
	.combout(),
	.sumout(Xd_0__inst_i19_41_sumout ),
	.cout(Xd_0__inst_i19_42 ),
	.shareout(Xd_0__inst_i19_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_22__0__q  $ (!Xd_0__inst_product_23__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_22__0__q  $ (!Xd_0__inst_product_23__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_22__0__q  & ((!Xd_0__inst_sign [23] & ((Xd_0__inst_sign [22]))) # (Xd_0__inst_sign [23] & (!Xd_0__inst_product_23__0__q )))) # (Xd_0__inst_product_22__0__q  & ((!Xd_0__inst_sign [23] 
// & (Xd_0__inst_product_23__0__q )) # (Xd_0__inst_sign [23] & ((!Xd_0__inst_sign [22]))))))

	.dataa(!Xd_0__inst_product_22__0__q ),
	.datab(!Xd_0__inst_product_23__0__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_20__0__q  $ (!Xd_0__inst_product_21__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_20__0__q  $ (!Xd_0__inst_product_21__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_20__0__q  & ((!Xd_0__inst_sign [21] & ((Xd_0__inst_sign [20]))) # (Xd_0__inst_sign [21] & (!Xd_0__inst_product_21__0__q )))) # (Xd_0__inst_product_20__0__q  & ((!Xd_0__inst_sign [21] 
// & (Xd_0__inst_product_21__0__q )) # (Xd_0__inst_sign [21] & ((!Xd_0__inst_sign [20]))))))

	.dataa(!Xd_0__inst_product_20__0__q ),
	.datab(!Xd_0__inst_product_21__0__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_18__0__q  $ (!Xd_0__inst_product_19__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_18__0__q  $ (!Xd_0__inst_product_19__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_18__0__q  & ((!Xd_0__inst_sign [19] & ((Xd_0__inst_sign [18]))) # (Xd_0__inst_sign [19] & (!Xd_0__inst_product_19__0__q )))) # (Xd_0__inst_product_18__0__q  & ((!Xd_0__inst_sign [19] 
// & (Xd_0__inst_product_19__0__q )) # (Xd_0__inst_sign [19] & ((!Xd_0__inst_sign [18]))))))

	.dataa(!Xd_0__inst_product_18__0__q ),
	.datab(!Xd_0__inst_product_19__0__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_45 (
// Equation(s):
// Xd_0__inst_i19_45_sumout  = SUM(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i19_67  ) + ( Xd_0__inst_i19_66  ))
// Xd_0__inst_i19_46  = CARRY(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i19_67  ) + ( Xd_0__inst_i19_66  ))
// Xd_0__inst_i19_47  = SHARE(GND)

	.dataa(!din_a[167]),
	.datab(!din_b[167]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_66 ),
	.sharein(Xd_0__inst_i19_67 ),
	.combout(),
	.sumout(Xd_0__inst_i19_45_sumout ),
	.cout(Xd_0__inst_i19_46 ),
	.shareout(Xd_0__inst_i19_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_16__0__q  $ (!Xd_0__inst_product_17__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_16__0__q  $ (!Xd_0__inst_product_17__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_16__0__q  & ((!Xd_0__inst_sign [17] & ((Xd_0__inst_sign [16]))) # (Xd_0__inst_sign [17] & (!Xd_0__inst_product_17__0__q )))) # (Xd_0__inst_product_16__0__q  & ((!Xd_0__inst_sign [17] 
// & (Xd_0__inst_product_17__0__q )) # (Xd_0__inst_sign [17] & ((!Xd_0__inst_sign [16]))))))

	.dataa(!Xd_0__inst_product_16__0__q ),
	.datab(!Xd_0__inst_product_17__0__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] & ((Xd_0__inst_sign [14]))) # (Xd_0__inst_sign [15] & (!Xd_0__inst_product_15__0__q )))) # (Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] 
// & (Xd_0__inst_product_15__0__q )) # (Xd_0__inst_sign [15] & ((!Xd_0__inst_sign [14]))))))

	.dataa(!Xd_0__inst_product_14__0__q ),
	.datab(!Xd_0__inst_product_15__0__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] & ((Xd_0__inst_sign [12]))) # (Xd_0__inst_sign [13] & (!Xd_0__inst_product_13__0__q )))) # (Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] 
// & (Xd_0__inst_product_13__0__q )) # (Xd_0__inst_sign [13] & ((!Xd_0__inst_sign [12]))))))

	.dataa(!Xd_0__inst_product_12__0__q ),
	.datab(!Xd_0__inst_product_13__0__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_49 (
// Equation(s):
// Xd_0__inst_i19_49_sumout  = SUM(( !din_a[139] $ (!din_b[139]) ) + ( Xd_0__inst_i19_71  ) + ( Xd_0__inst_i19_70  ))
// Xd_0__inst_i19_50  = CARRY(( !din_a[139] $ (!din_b[139]) ) + ( Xd_0__inst_i19_71  ) + ( Xd_0__inst_i19_70  ))
// Xd_0__inst_i19_51  = SHARE(GND)

	.dataa(!din_a[139]),
	.datab(!din_b[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_70 ),
	.sharein(Xd_0__inst_i19_71 ),
	.combout(),
	.sumout(Xd_0__inst_i19_49_sumout ),
	.cout(Xd_0__inst_i19_50 ),
	.shareout(Xd_0__inst_i19_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] & ((Xd_0__inst_sign [10]))) # (Xd_0__inst_sign [11] & (!Xd_0__inst_product_11__0__q )))) # (Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] 
// & (Xd_0__inst_product_11__0__q )) # (Xd_0__inst_sign [11] & ((!Xd_0__inst_sign [10]))))))

	.dataa(!Xd_0__inst_product_10__0__q ),
	.datab(!Xd_0__inst_product_11__0__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_4__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & ((Xd_0__inst_sign [8]))) # (Xd_0__inst_sign [9] & (!Xd_0__inst_product_9__0__q )))) # (Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & 
// (Xd_0__inst_product_9__0__q )) # (Xd_0__inst_sign [9] & ((!Xd_0__inst_sign [8]))))))

	.dataa(!Xd_0__inst_product_8__0__q ),
	.datab(!Xd_0__inst_product_9__0__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_3__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & ((Xd_0__inst_sign [6]))) # (Xd_0__inst_sign [7] & (!Xd_0__inst_product_7__0__q )))) # (Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & 
// (Xd_0__inst_product_7__0__q )) # (Xd_0__inst_sign [7] & ((!Xd_0__inst_sign [6]))))))

	.dataa(!Xd_0__inst_product_6__0__q ),
	.datab(!Xd_0__inst_product_7__0__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_53 (
// Equation(s):
// Xd_0__inst_i19_53_sumout  = SUM(( !din_a[111] $ (!din_b[111]) ) + ( Xd_0__inst_i19_75  ) + ( Xd_0__inst_i19_74  ))
// Xd_0__inst_i19_54  = CARRY(( !din_a[111] $ (!din_b[111]) ) + ( Xd_0__inst_i19_75  ) + ( Xd_0__inst_i19_74  ))
// Xd_0__inst_i19_55  = SHARE(GND)

	.dataa(!din_a[111]),
	.datab(!din_b[111]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_74 ),
	.sharein(Xd_0__inst_i19_75 ),
	.combout(),
	.sumout(Xd_0__inst_i19_53_sumout ),
	.cout(Xd_0__inst_i19_54 ),
	.shareout(Xd_0__inst_i19_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_2__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & ((Xd_0__inst_sign [4]))) # (Xd_0__inst_sign [5] & (!Xd_0__inst_product_5__0__q )))) # (Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & 
// (Xd_0__inst_product_5__0__q )) # (Xd_0__inst_sign [5] & ((!Xd_0__inst_sign [4]))))))

	.dataa(!Xd_0__inst_product_4__0__q ),
	.datab(!Xd_0__inst_product_5__0__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_i19_79  ) + ( Xd_0__inst_i19_78  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_i19_79  ) + ( Xd_0__inst_i19_78  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & ((Xd_0__inst_sign [2]))) # (Xd_0__inst_sign [3] & (!Xd_0__inst_product_3__0__q )))) # (Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & 
// (Xd_0__inst_product_3__0__q )) # (Xd_0__inst_sign [3] & ((!Xd_0__inst_sign [2]))))))

	.dataa(!Xd_0__inst_product_2__0__q ),
	.datab(!Xd_0__inst_product_3__0__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_78 ),
	.sharein(Xd_0__inst_i19_79 ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_i19_83  ) + ( Xd_0__inst_i19_82  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_i19_83  ) + ( Xd_0__inst_i19_82  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & ((Xd_0__inst_sign [0]))) # (Xd_0__inst_sign [1] & (!Xd_0__inst_product_1__0__q )))) # (Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & 
// (Xd_0__inst_product_1__0__q )) # (Xd_0__inst_sign [1] & ((!Xd_0__inst_sign [0]))))))

	.dataa(!Xd_0__inst_product_0__0__q ),
	.datab(!Xd_0__inst_product_1__0__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_82 ),
	.sharein(Xd_0__inst_i19_83 ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_57 (
// Equation(s):
// Xd_0__inst_i19_57_sumout  = SUM(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i19_87  ) + ( Xd_0__inst_i19_86  ))
// Xd_0__inst_i19_58  = CARRY(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i19_87  ) + ( Xd_0__inst_i19_86  ))
// Xd_0__inst_i19_59  = SHARE(GND)

	.dataa(!din_a[83]),
	.datab(!din_b[83]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_86 ),
	.sharein(Xd_0__inst_i19_87 ),
	.combout(),
	.sumout(Xd_0__inst_i19_57_sumout ),
	.cout(Xd_0__inst_i19_58 ),
	.shareout(Xd_0__inst_i19_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_28__1__q  $ (!Xd_0__inst_product_29__1__q  $ (((Xd_0__inst_sign [29]) # (Xd_0__inst_sign [28])))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_28__1__q  $ (!Xd_0__inst_product_29__1__q  $ (((Xd_0__inst_sign [29]) # (Xd_0__inst_sign [28])))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [28] & (Xd_0__inst_product_28__1__q  & (!Xd_0__inst_product_29__1__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_sign [28] & ((!Xd_0__inst_product_29__1__q  & ((Xd_0__inst_sign [29]))) 
// # (Xd_0__inst_product_29__1__q  & (!Xd_0__inst_product_28__1__q )))))

	.dataa(!Xd_0__inst_product_28__1__q ),
	.datab(!Xd_0__inst_product_29__1__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_26__1__q  $ (!Xd_0__inst_product_27__1__q  $ (((Xd_0__inst_sign [27]) # (Xd_0__inst_sign [26])))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_26__1__q  $ (!Xd_0__inst_product_27__1__q  $ (((Xd_0__inst_sign [27]) # (Xd_0__inst_sign [26])))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [26] & (Xd_0__inst_product_26__1__q  & (!Xd_0__inst_product_27__1__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_sign [26] & ((!Xd_0__inst_product_27__1__q  & ((Xd_0__inst_sign [27]))) 
// # (Xd_0__inst_product_27__1__q  & (!Xd_0__inst_product_26__1__q )))))

	.dataa(!Xd_0__inst_product_26__1__q ),
	.datab(!Xd_0__inst_product_27__1__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_24__1__q  $ (!Xd_0__inst_product_25__1__q  $ (((Xd_0__inst_sign [25]) # (Xd_0__inst_sign [24])))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_24__1__q  $ (!Xd_0__inst_product_25__1__q  $ (((Xd_0__inst_sign [25]) # (Xd_0__inst_sign [24])))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [24] & (Xd_0__inst_product_24__1__q  & (!Xd_0__inst_product_25__1__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_sign [24] & ((!Xd_0__inst_product_25__1__q  & ((Xd_0__inst_sign [25]))) 
// # (Xd_0__inst_product_25__1__q  & (!Xd_0__inst_product_24__1__q )))))

	.dataa(!Xd_0__inst_product_24__1__q ),
	.datab(!Xd_0__inst_product_25__1__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_22__1__q  $ (!Xd_0__inst_product_23__1__q  $ (((Xd_0__inst_sign [23]) # (Xd_0__inst_sign [22])))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_22__1__q  $ (!Xd_0__inst_product_23__1__q  $ (((Xd_0__inst_sign [23]) # (Xd_0__inst_sign [22])))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [22] & (Xd_0__inst_product_22__1__q  & (!Xd_0__inst_product_23__1__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_sign [22] & ((!Xd_0__inst_product_23__1__q  & ((Xd_0__inst_sign [23]))) 
// # (Xd_0__inst_product_23__1__q  & (!Xd_0__inst_product_22__1__q )))))

	.dataa(!Xd_0__inst_product_22__1__q ),
	.datab(!Xd_0__inst_product_23__1__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_20__1__q  $ (!Xd_0__inst_product_21__1__q  $ (((Xd_0__inst_sign [21]) # (Xd_0__inst_sign [20])))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_20__1__q  $ (!Xd_0__inst_product_21__1__q  $ (((Xd_0__inst_sign [21]) # (Xd_0__inst_sign [20])))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [20] & (Xd_0__inst_product_20__1__q  & (!Xd_0__inst_product_21__1__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_sign [20] & ((!Xd_0__inst_product_21__1__q  & ((Xd_0__inst_sign [21]))) 
// # (Xd_0__inst_product_21__1__q  & (!Xd_0__inst_product_20__1__q )))))

	.dataa(!Xd_0__inst_product_20__1__q ),
	.datab(!Xd_0__inst_product_21__1__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_18__1__q  $ (!Xd_0__inst_product_19__1__q  $ (((Xd_0__inst_sign [19]) # (Xd_0__inst_sign [18])))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_18__1__q  $ (!Xd_0__inst_product_19__1__q  $ (((Xd_0__inst_sign [19]) # (Xd_0__inst_sign [18])))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [18] & (Xd_0__inst_product_18__1__q  & (!Xd_0__inst_product_19__1__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_sign [18] & ((!Xd_0__inst_product_19__1__q  & ((Xd_0__inst_sign [19]))) # 
// (Xd_0__inst_product_19__1__q  & (!Xd_0__inst_product_18__1__q )))))

	.dataa(!Xd_0__inst_product_18__1__q ),
	.datab(!Xd_0__inst_product_19__1__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_16__1__q  $ (!Xd_0__inst_product_17__1__q  $ (((Xd_0__inst_sign [17]) # (Xd_0__inst_sign [16])))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_16__1__q  $ (!Xd_0__inst_product_17__1__q  $ (((Xd_0__inst_sign [17]) # (Xd_0__inst_sign [16])))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [16] & (Xd_0__inst_product_16__1__q  & (!Xd_0__inst_product_17__1__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_sign [16] & ((!Xd_0__inst_product_17__1__q  & ((Xd_0__inst_sign [17]))) # 
// (Xd_0__inst_product_17__1__q  & (!Xd_0__inst_product_16__1__q )))))

	.dataa(!Xd_0__inst_product_16__1__q ),
	.datab(!Xd_0__inst_product_17__1__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [14] & (Xd_0__inst_product_14__1__q  & (!Xd_0__inst_product_15__1__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_sign [14] & ((!Xd_0__inst_product_15__1__q  & ((Xd_0__inst_sign [15]))) # 
// (Xd_0__inst_product_15__1__q  & (!Xd_0__inst_product_14__1__q )))))

	.dataa(!Xd_0__inst_product_14__1__q ),
	.datab(!Xd_0__inst_product_15__1__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [12] & (Xd_0__inst_product_12__1__q  & (!Xd_0__inst_product_13__1__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_sign [12] & ((!Xd_0__inst_product_13__1__q  & ((Xd_0__inst_sign [13]))) # 
// (Xd_0__inst_product_13__1__q  & (!Xd_0__inst_product_12__1__q )))))

	.dataa(!Xd_0__inst_product_12__1__q ),
	.datab(!Xd_0__inst_product_13__1__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [10] & (Xd_0__inst_product_10__1__q  & (!Xd_0__inst_product_11__1__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_sign [10] & ((!Xd_0__inst_product_11__1__q  & ((Xd_0__inst_sign [11]))) # 
// (Xd_0__inst_product_11__1__q  & (!Xd_0__inst_product_10__1__q )))))

	.dataa(!Xd_0__inst_product_10__1__q ),
	.datab(!Xd_0__inst_product_11__1__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [8] & (Xd_0__inst_product_8__1__q  & (!Xd_0__inst_product_9__1__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_sign [8] & ((!Xd_0__inst_product_9__1__q  & ((Xd_0__inst_sign [9]))) # 
// (Xd_0__inst_product_9__1__q  & (!Xd_0__inst_product_8__1__q )))))

	.dataa(!Xd_0__inst_product_8__1__q ),
	.datab(!Xd_0__inst_product_9__1__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [6] & (Xd_0__inst_product_6__1__q  & (!Xd_0__inst_product_7__1__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_sign [6] & ((!Xd_0__inst_product_7__1__q  & ((Xd_0__inst_sign [7]))) # 
// (Xd_0__inst_product_7__1__q  & (!Xd_0__inst_product_6__1__q )))))

	.dataa(!Xd_0__inst_product_6__1__q ),
	.datab(!Xd_0__inst_product_7__1__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [4] & (Xd_0__inst_product_4__1__q  & (!Xd_0__inst_product_5__1__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_sign [4] & ((!Xd_0__inst_product_5__1__q  & ((Xd_0__inst_sign [5]))) # 
// (Xd_0__inst_product_5__1__q  & (!Xd_0__inst_product_4__1__q )))))

	.dataa(!Xd_0__inst_product_4__1__q ),
	.datab(!Xd_0__inst_product_5__1__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [2] & (Xd_0__inst_product_2__1__q  & (!Xd_0__inst_product_3__1__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_sign [2] & ((!Xd_0__inst_product_3__1__q  & ((Xd_0__inst_sign [3]))) # 
// (Xd_0__inst_product_3__1__q  & (!Xd_0__inst_product_2__1__q )))))

	.dataa(!Xd_0__inst_product_2__1__q ),
	.datab(!Xd_0__inst_product_3__1__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [0] & (Xd_0__inst_product_0__1__q  & (!Xd_0__inst_product_1__1__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_sign [0] & ((!Xd_0__inst_product_1__1__q  & ((Xd_0__inst_sign [1]))) # 
// (Xd_0__inst_product_1__1__q  & (!Xd_0__inst_product_0__1__q )))))

	.dataa(!Xd_0__inst_product_0__1__q ),
	.datab(!Xd_0__inst_product_1__1__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_28__2__q  $ (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_28__2__q  $ (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__2__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__2__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__2__q ),
	.datab(!Xd_0__inst_product_29__2__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_26__2__q  $ (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_26__2__q  $ (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__2__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__2__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__2__q ),
	.datab(!Xd_0__inst_product_27__2__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_24__2__q  $ (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_24__2__q  $ (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__2__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__2__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__2__q ),
	.datab(!Xd_0__inst_product_25__2__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_22__2__q  $ (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_22__2__q  $ (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__2__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__2__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__2__q ),
	.datab(!Xd_0__inst_product_23__2__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_20__2__q  $ (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_20__2__q  $ (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__2__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__2__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__2__q ),
	.datab(!Xd_0__inst_product_21__2__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_18__2__q  $ (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_18__2__q  $ (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__2__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__2__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__2__q ),
	.datab(!Xd_0__inst_product_19__2__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_16__2__q  $ (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_16__2__q  $ (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__2__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__2__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__2__q ),
	.datab(!Xd_0__inst_product_17__2__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__2__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__2__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__2__q ),
	.datab(!Xd_0__inst_product_15__2__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__2__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__2__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__2__q ),
	.datab(!Xd_0__inst_product_13__2__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__2__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__2__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__2__q ),
	.datab(!Xd_0__inst_product_11__2__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__2__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__2__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__2__q ),
	.datab(!Xd_0__inst_product_9__2__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__2__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__2__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__2__q ),
	.datab(!Xd_0__inst_product_7__2__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__2__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__2__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__2__q ),
	.datab(!Xd_0__inst_product_5__2__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__2__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__2__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__2__q ),
	.datab(!Xd_0__inst_product_3__2__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__2__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__2__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__2__q ),
	.datab(!Xd_0__inst_product_1__2__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_28__3__q  $ (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_28__3__q  $ (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__3__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__3__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__3__q ),
	.datab(!Xd_0__inst_product_29__3__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_26__3__q  $ (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_26__3__q  $ (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__3__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__3__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__3__q ),
	.datab(!Xd_0__inst_product_27__3__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_24__3__q  $ (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_24__3__q  $ (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__3__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__3__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__3__q ),
	.datab(!Xd_0__inst_product_25__3__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_22__3__q  $ (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_22__3__q  $ (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__3__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__3__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__3__q ),
	.datab(!Xd_0__inst_product_23__3__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_20__3__q  $ (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_20__3__q  $ (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__3__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__3__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__3__q ),
	.datab(!Xd_0__inst_product_21__3__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_18__3__q  $ (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_18__3__q  $ (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__3__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__3__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__3__q ),
	.datab(!Xd_0__inst_product_19__3__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_16__3__q  $ (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_16__3__q  $ (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__3__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__3__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__3__q ),
	.datab(!Xd_0__inst_product_17__3__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__3__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__3__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__3__q ),
	.datab(!Xd_0__inst_product_15__3__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__3__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__3__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__3__q ),
	.datab(!Xd_0__inst_product_13__3__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__3__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__3__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__3__q ),
	.datab(!Xd_0__inst_product_11__3__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__3__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__3__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__3__q ),
	.datab(!Xd_0__inst_product_9__3__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__3__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__3__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__3__q ),
	.datab(!Xd_0__inst_product_7__3__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__3__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__3__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__3__q ),
	.datab(!Xd_0__inst_product_5__3__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__3__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__3__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__3__q ),
	.datab(!Xd_0__inst_product_3__3__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__3__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__3__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__3__q ),
	.datab(!Xd_0__inst_product_1__3__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_28__4__q  $ (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_28__4__q  $ (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__4__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__4__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__4__q ),
	.datab(!Xd_0__inst_product_29__4__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_26__4__q  $ (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_26__4__q  $ (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__4__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__4__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__4__q ),
	.datab(!Xd_0__inst_product_27__4__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_24__4__q  $ (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_24__4__q  $ (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__4__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__4__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__4__q ),
	.datab(!Xd_0__inst_product_25__4__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_22__4__q  $ (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_22__4__q  $ (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__4__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__4__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__4__q ),
	.datab(!Xd_0__inst_product_23__4__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_20__4__q  $ (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_20__4__q  $ (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__4__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__4__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__4__q ),
	.datab(!Xd_0__inst_product_21__4__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_18__4__q  $ (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_18__4__q  $ (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__4__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__4__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__4__q ),
	.datab(!Xd_0__inst_product_19__4__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_16__4__q  $ (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_16__4__q  $ (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__4__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__4__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__4__q ),
	.datab(!Xd_0__inst_product_17__4__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__4__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__4__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__4__q ),
	.datab(!Xd_0__inst_product_15__4__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__4__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__4__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__4__q ),
	.datab(!Xd_0__inst_product_13__4__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__4__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__4__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__4__q ),
	.datab(!Xd_0__inst_product_11__4__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__4__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__4__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__4__q ),
	.datab(!Xd_0__inst_product_9__4__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__4__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__4__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__4__q ),
	.datab(!Xd_0__inst_product_7__4__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__4__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__4__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__4__q ),
	.datab(!Xd_0__inst_product_5__4__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__4__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__4__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__4__q ),
	.datab(!Xd_0__inst_product_3__4__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__4__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__4__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__4__q ),
	.datab(!Xd_0__inst_product_1__4__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_28__5__q  $ (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_28__5__q  $ (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__5__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__5__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__5__q ),
	.datab(!Xd_0__inst_product_29__5__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_26__5__q  $ (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_26__5__q  $ (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__5__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__5__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__5__q ),
	.datab(!Xd_0__inst_product_27__5__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_24__5__q  $ (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_24__5__q  $ (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__5__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__5__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__5__q ),
	.datab(!Xd_0__inst_product_25__5__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_22__5__q  $ (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_22__5__q  $ (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__5__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__5__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__5__q ),
	.datab(!Xd_0__inst_product_23__5__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_20__5__q  $ (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_20__5__q  $ (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__5__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__5__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__5__q ),
	.datab(!Xd_0__inst_product_21__5__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_18__5__q  $ (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_18__5__q  $ (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__5__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__5__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__5__q ),
	.datab(!Xd_0__inst_product_19__5__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_16__5__q  $ (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_16__5__q  $ (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__5__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__5__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__5__q ),
	.datab(!Xd_0__inst_product_17__5__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__5__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__5__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__5__q ),
	.datab(!Xd_0__inst_product_15__5__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__5__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__5__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__5__q ),
	.datab(!Xd_0__inst_product_13__5__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__5__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__5__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__5__q ),
	.datab(!Xd_0__inst_product_11__5__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__5__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__5__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__5__q ),
	.datab(!Xd_0__inst_product_9__5__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__5__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__5__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__5__q ),
	.datab(!Xd_0__inst_product_7__5__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__5__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__5__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__5__q ),
	.datab(!Xd_0__inst_product_5__5__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__5__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__5__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__5__q ),
	.datab(!Xd_0__inst_product_3__5__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__5__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__5__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__5__q ),
	.datab(!Xd_0__inst_product_1__5__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_28__6__q  $ (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_28__6__q  $ (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__6__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__6__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__6__q ),
	.datab(!Xd_0__inst_product_29__6__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_26__6__q  $ (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_26__6__q  $ (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__6__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__6__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__6__q ),
	.datab(!Xd_0__inst_product_27__6__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_24__6__q  $ (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_24__6__q  $ (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__6__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__6__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__6__q ),
	.datab(!Xd_0__inst_product_25__6__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_22__6__q  $ (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_22__6__q  $ (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__6__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__6__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__6__q ),
	.datab(!Xd_0__inst_product_23__6__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_20__6__q  $ (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_20__6__q  $ (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__6__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__6__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__6__q ),
	.datab(!Xd_0__inst_product_21__6__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_18__6__q  $ (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_18__6__q  $ (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__6__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__6__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__6__q ),
	.datab(!Xd_0__inst_product_19__6__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_16__6__q  $ (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_16__6__q  $ (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__6__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__6__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__6__q ),
	.datab(!Xd_0__inst_product_17__6__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__6__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__6__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__6__q ),
	.datab(!Xd_0__inst_product_15__6__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__6__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__6__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__6__q ),
	.datab(!Xd_0__inst_product_13__6__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__6__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__6__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__6__q ),
	.datab(!Xd_0__inst_product_11__6__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__6__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__6__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__6__q ),
	.datab(!Xd_0__inst_product_9__6__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__6__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__6__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__6__q ),
	.datab(!Xd_0__inst_product_7__6__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__6__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__6__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__6__q ),
	.datab(!Xd_0__inst_product_5__6__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__6__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__6__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__6__q ),
	.datab(!Xd_0__inst_product_3__6__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__6__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__6__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__6__q ),
	.datab(!Xd_0__inst_product_1__6__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_28__7__q  $ (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_28__7__q  $ (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__7__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__7__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__7__q ),
	.datab(!Xd_0__inst_product_29__7__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_26__7__q  $ (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_26__7__q  $ (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__7__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__7__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__7__q ),
	.datab(!Xd_0__inst_product_27__7__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_24__7__q  $ (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_24__7__q  $ (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__7__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__7__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__7__q ),
	.datab(!Xd_0__inst_product_25__7__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_22__7__q  $ (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_22__7__q  $ (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__7__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__7__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__7__q ),
	.datab(!Xd_0__inst_product_23__7__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_20__7__q  $ (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_20__7__q  $ (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__7__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__7__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__7__q ),
	.datab(!Xd_0__inst_product_21__7__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_18__7__q  $ (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_18__7__q  $ (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__7__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__7__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__7__q ),
	.datab(!Xd_0__inst_product_19__7__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_16__7__q  $ (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_16__7__q  $ (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__7__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__7__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__7__q ),
	.datab(!Xd_0__inst_product_17__7__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__7__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__7__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__7__q ),
	.datab(!Xd_0__inst_product_15__7__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__7__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__7__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__7__q ),
	.datab(!Xd_0__inst_product_13__7__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__7__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__7__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__7__q ),
	.datab(!Xd_0__inst_product_11__7__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__7__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__7__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__7__q ),
	.datab(!Xd_0__inst_product_9__7__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__7__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__7__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__7__q ),
	.datab(!Xd_0__inst_product_7__7__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__7__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__7__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__7__q ),
	.datab(!Xd_0__inst_product_5__7__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__7__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__7__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__7__q ),
	.datab(!Xd_0__inst_product_3__7__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__7__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__7__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__7__q ),
	.datab(!Xd_0__inst_product_1__7__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_28__8__q  $ (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_28__8__q  $ (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__8__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__8__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__8__q ),
	.datab(!Xd_0__inst_product_29__8__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_26__8__q  $ (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_26__8__q  $ (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__8__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__8__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__8__q ),
	.datab(!Xd_0__inst_product_27__8__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_24__8__q  $ (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_24__8__q  $ (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__8__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__8__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__8__q ),
	.datab(!Xd_0__inst_product_25__8__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_22__8__q  $ (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_22__8__q  $ (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__8__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__8__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__8__q ),
	.datab(!Xd_0__inst_product_23__8__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_20__8__q  $ (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_20__8__q  $ (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__8__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__8__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__8__q ),
	.datab(!Xd_0__inst_product_21__8__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_18__8__q  $ (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_18__8__q  $ (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__8__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__8__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__8__q ),
	.datab(!Xd_0__inst_product_19__8__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_16__8__q  $ (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_16__8__q  $ (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__8__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__8__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__8__q ),
	.datab(!Xd_0__inst_product_17__8__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__8__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__8__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__8__q ),
	.datab(!Xd_0__inst_product_15__8__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__8__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__8__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__8__q ),
	.datab(!Xd_0__inst_product_13__8__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__8__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__8__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__8__q ),
	.datab(!Xd_0__inst_product_11__8__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__8__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__8__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__8__q ),
	.datab(!Xd_0__inst_product_9__8__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__8__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__8__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__8__q ),
	.datab(!Xd_0__inst_product_7__8__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__8__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__8__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__8__q ),
	.datab(!Xd_0__inst_product_5__8__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__8__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__8__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__8__q ),
	.datab(!Xd_0__inst_product_3__8__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__8__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__8__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__8__q ),
	.datab(!Xd_0__inst_product_1__8__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_28__9__q  $ (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_28__9__q  $ (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__9__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__9__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__9__q ),
	.datab(!Xd_0__inst_product_29__9__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_26__9__q  $ (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_26__9__q  $ (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__9__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__9__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__9__q ),
	.datab(!Xd_0__inst_product_27__9__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_24__9__q  $ (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_24__9__q  $ (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__9__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__9__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__9__q ),
	.datab(!Xd_0__inst_product_25__9__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_22__9__q  $ (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_22__9__q  $ (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__9__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__9__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__9__q ),
	.datab(!Xd_0__inst_product_23__9__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_20__9__q  $ (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_20__9__q  $ (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__9__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__9__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__9__q ),
	.datab(!Xd_0__inst_product_21__9__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_18__9__q  $ (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_18__9__q  $ (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__9__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__9__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__9__q ),
	.datab(!Xd_0__inst_product_19__9__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_16__9__q  $ (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_16__9__q  $ (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__9__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__9__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__9__q ),
	.datab(!Xd_0__inst_product_17__9__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__9__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__9__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__9__q ),
	.datab(!Xd_0__inst_product_15__9__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__9__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__9__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__9__q ),
	.datab(!Xd_0__inst_product_13__9__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__9__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__9__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__9__q ),
	.datab(!Xd_0__inst_product_11__9__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__9__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__9__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__9__q ),
	.datab(!Xd_0__inst_product_9__9__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__9__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__9__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__9__q ),
	.datab(!Xd_0__inst_product_7__9__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__9__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__9__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__9__q ),
	.datab(!Xd_0__inst_product_5__9__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__9__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__9__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__9__q ),
	.datab(!Xd_0__inst_product_3__9__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__9__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__9__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__9__q ),
	.datab(!Xd_0__inst_product_1__9__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_28__10__q  $ (!Xd_0__inst_product_29__10__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_28__10__q  $ (!Xd_0__inst_product_29__10__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__10__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__10__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__10__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__10__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__10__q ),
	.datab(!Xd_0__inst_product_29__10__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_26__10__q  $ (!Xd_0__inst_product_27__10__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_26__10__q  $ (!Xd_0__inst_product_27__10__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__10__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__10__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__10__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__10__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__10__q ),
	.datab(!Xd_0__inst_product_27__10__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_24__10__q  $ (!Xd_0__inst_product_25__10__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_24__10__q  $ (!Xd_0__inst_product_25__10__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__10__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__10__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__10__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__10__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__10__q ),
	.datab(!Xd_0__inst_product_25__10__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_22__10__q  $ (!Xd_0__inst_product_23__10__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_22__10__q  $ (!Xd_0__inst_product_23__10__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__10__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__10__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__10__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__10__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__10__q ),
	.datab(!Xd_0__inst_product_23__10__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_20__10__q  $ (!Xd_0__inst_product_21__10__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_20__10__q  $ (!Xd_0__inst_product_21__10__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__10__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__10__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__10__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__10__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__10__q ),
	.datab(!Xd_0__inst_product_21__10__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_18__10__q  $ (!Xd_0__inst_product_19__10__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_18__10__q  $ (!Xd_0__inst_product_19__10__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__10__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__10__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__10__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__10__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__10__q ),
	.datab(!Xd_0__inst_product_19__10__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_16__10__q  $ (!Xd_0__inst_product_17__10__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_16__10__q  $ (!Xd_0__inst_product_17__10__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__10__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__10__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__10__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__10__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__10__q ),
	.datab(!Xd_0__inst_product_17__10__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_14__10__q  $ (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_14__10__q  $ (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__10__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__10__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__10__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__10__q ),
	.datab(!Xd_0__inst_product_15__10__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_12__10__q  $ (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_12__10__q  $ (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__10__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__10__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__10__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__10__q ),
	.datab(!Xd_0__inst_product_13__10__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_10__10__q  $ (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_10__10__q  $ (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__10__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__10__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__10__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__10__q ),
	.datab(!Xd_0__inst_product_11__10__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_8__10__q  $ (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_8__10__q  $ (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__10__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__10__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__10__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__10__q ),
	.datab(!Xd_0__inst_product_9__10__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__10__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__10__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__10__q ),
	.datab(!Xd_0__inst_product_7__10__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__10__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__10__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__10__q ),
	.datab(!Xd_0__inst_product_5__10__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__10__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__10__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__10__q ),
	.datab(!Xd_0__inst_product_3__10__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__10__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__10__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__10__q ),
	.datab(!Xd_0__inst_product_1__10__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_28__11__q  $ (!Xd_0__inst_product_29__11__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_28__11__q  $ (!Xd_0__inst_product_29__11__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__11__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__11__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__11__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__11__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__11__q ),
	.datab(!Xd_0__inst_product_29__11__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_26__11__q  $ (!Xd_0__inst_product_27__11__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_26__11__q  $ (!Xd_0__inst_product_27__11__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__11__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__11__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__11__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__11__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__11__q ),
	.datab(!Xd_0__inst_product_27__11__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_24__11__q  $ (!Xd_0__inst_product_25__11__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_24__11__q  $ (!Xd_0__inst_product_25__11__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__11__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__11__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__11__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__11__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__11__q ),
	.datab(!Xd_0__inst_product_25__11__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_22__11__q  $ (!Xd_0__inst_product_23__11__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_22__11__q  $ (!Xd_0__inst_product_23__11__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__11__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__11__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__11__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__11__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__11__q ),
	.datab(!Xd_0__inst_product_23__11__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_20__11__q  $ (!Xd_0__inst_product_21__11__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_20__11__q  $ (!Xd_0__inst_product_21__11__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__11__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__11__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__11__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__11__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__11__q ),
	.datab(!Xd_0__inst_product_21__11__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_18__11__q  $ (!Xd_0__inst_product_19__11__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_18__11__q  $ (!Xd_0__inst_product_19__11__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__11__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__11__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__11__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__11__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__11__q ),
	.datab(!Xd_0__inst_product_19__11__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_16__11__q  $ (!Xd_0__inst_product_17__11__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_16__11__q  $ (!Xd_0__inst_product_17__11__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__11__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__11__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__11__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__11__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__11__q ),
	.datab(!Xd_0__inst_product_17__11__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_14__11__q  $ (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_14__11__q  $ (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__11__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__11__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__11__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__11__q ),
	.datab(!Xd_0__inst_product_15__11__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_12__11__q  $ (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_12__11__q  $ (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__11__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__11__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__11__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__11__q ),
	.datab(!Xd_0__inst_product_13__11__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_10__11__q  $ (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_10__11__q  $ (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__11__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__11__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__11__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__11__q ),
	.datab(!Xd_0__inst_product_11__11__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_8__11__q  $ (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_8__11__q  $ (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__11__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__11__q  & (!Xd_0__inst_sign [8] & 
// (!Xd_0__inst_product_9__11__q  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__11__q ),
	.datab(!Xd_0__inst_product_9__11__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__11__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__11__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__11__q ),
	.datab(!Xd_0__inst_product_7__11__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__11__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__11__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__11__q ),
	.datab(!Xd_0__inst_product_5__11__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__11__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__11__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__11__q ),
	.datab(!Xd_0__inst_product_3__11__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__11__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__11__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__11__q ),
	.datab(!Xd_0__inst_product_1__11__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [28] & Xd_0__inst_sign [29]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [26] & Xd_0__inst_sign [27]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [24] & Xd_0__inst_sign [25]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [22] & Xd_0__inst_sign [23]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [20] & Xd_0__inst_sign [21]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [18] & Xd_0__inst_sign [19]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [16] & Xd_0__inst_sign [17]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [14] & Xd_0__inst_sign [15]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [12] & Xd_0__inst_sign [13]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [10] & Xd_0__inst_sign [11]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [8] & Xd_0__inst_sign [9]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [6] & Xd_0__inst_sign [7]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [4] & Xd_0__inst_sign [5]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [2] & Xd_0__inst_sign [3]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [12] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [0] & Xd_0__inst_sign [1]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [13] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_61 (
// Equation(s):
// Xd_0__inst_i19_61_sumout  = SUM(( !din_a[174] $ (!din_b[174]) ) + ( Xd_0__inst_i19_91  ) + ( Xd_0__inst_i19_90  ))
// Xd_0__inst_i19_62  = CARRY(( !din_a[174] $ (!din_b[174]) ) + ( Xd_0__inst_i19_91  ) + ( Xd_0__inst_i19_90  ))
// Xd_0__inst_i19_63  = SHARE(GND)

	.dataa(!din_a[174]),
	.datab(!din_b[174]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_90 ),
	.sharein(Xd_0__inst_i19_91 ),
	.combout(),
	.sumout(Xd_0__inst_i19_61_sumout ),
	.cout(Xd_0__inst_i19_62 ),
	.shareout(Xd_0__inst_i19_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_65 (
// Equation(s):
// Xd_0__inst_i19_65_sumout  = SUM(( !din_a[146] $ (!din_b[146]) ) + ( Xd_0__inst_i19_95  ) + ( Xd_0__inst_i19_94  ))
// Xd_0__inst_i19_66  = CARRY(( !din_a[146] $ (!din_b[146]) ) + ( Xd_0__inst_i19_95  ) + ( Xd_0__inst_i19_94  ))
// Xd_0__inst_i19_67  = SHARE(GND)

	.dataa(!din_a[146]),
	.datab(!din_b[146]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_94 ),
	.sharein(Xd_0__inst_i19_95 ),
	.combout(),
	.sumout(Xd_0__inst_i19_65_sumout ),
	.cout(Xd_0__inst_i19_66 ),
	.shareout(Xd_0__inst_i19_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_69 (
// Equation(s):
// Xd_0__inst_i19_69_sumout  = SUM(( !din_a[118] $ (!din_b[118]) ) + ( Xd_0__inst_i19_99  ) + ( Xd_0__inst_i19_98  ))
// Xd_0__inst_i19_70  = CARRY(( !din_a[118] $ (!din_b[118]) ) + ( Xd_0__inst_i19_99  ) + ( Xd_0__inst_i19_98  ))
// Xd_0__inst_i19_71  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[118]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_98 ),
	.sharein(Xd_0__inst_i19_99 ),
	.combout(),
	.sumout(Xd_0__inst_i19_69_sumout ),
	.cout(Xd_0__inst_i19_70 ),
	.shareout(Xd_0__inst_i19_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_73 (
// Equation(s):
// Xd_0__inst_i19_73_sumout  = SUM(( !din_a[90] $ (!din_b[90]) ) + ( Xd_0__inst_i19_103  ) + ( Xd_0__inst_i19_102  ))
// Xd_0__inst_i19_74  = CARRY(( !din_a[90] $ (!din_b[90]) ) + ( Xd_0__inst_i19_103  ) + ( Xd_0__inst_i19_102  ))
// Xd_0__inst_i19_75  = SHARE(GND)

	.dataa(!din_a[90]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_102 ),
	.sharein(Xd_0__inst_i19_103 ),
	.combout(),
	.sumout(Xd_0__inst_i19_73_sumout ),
	.cout(Xd_0__inst_i19_74 ),
	.shareout(Xd_0__inst_i19_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_77 (
// Equation(s):
// Xd_0__inst_i19_77_sumout  = SUM(( !din_a[6] $ (!din_b[6]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_78  = CARRY(( !din_a[6] $ (!din_b[6]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_79  = SHARE(GND)

	.dataa(!din_a[6]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_77_sumout ),
	.cout(Xd_0__inst_i19_78 ),
	.shareout(Xd_0__inst_i19_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_81 (
// Equation(s):
// Xd_0__inst_i19_81_sumout  = SUM(( !din_a[48] $ (!din_b[48]) ) + ( Xd_0__inst_i19_107  ) + ( Xd_0__inst_i19_106  ))
// Xd_0__inst_i19_82  = CARRY(( !din_a[48] $ (!din_b[48]) ) + ( Xd_0__inst_i19_107  ) + ( Xd_0__inst_i19_106  ))
// Xd_0__inst_i19_83  = SHARE(GND)

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_106 ),
	.sharein(Xd_0__inst_i19_107 ),
	.combout(),
	.sumout(Xd_0__inst_i19_81_sumout ),
	.cout(Xd_0__inst_i19_82 ),
	.shareout(Xd_0__inst_i19_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_85 (
// Equation(s):
// Xd_0__inst_i19_85_sumout  = SUM(( !din_a[62] $ (!din_b[62]) ) + ( Xd_0__inst_i19_111  ) + ( Xd_0__inst_i19_110  ))
// Xd_0__inst_i19_86  = CARRY(( !din_a[62] $ (!din_b[62]) ) + ( Xd_0__inst_i19_111  ) + ( Xd_0__inst_i19_110  ))
// Xd_0__inst_i19_87  = SHARE(GND)

	.dataa(!din_a[62]),
	.datab(!din_b[62]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_110 ),
	.sharein(Xd_0__inst_i19_111 ),
	.combout(),
	.sumout(Xd_0__inst_i19_85_sumout ),
	.cout(Xd_0__inst_i19_86 ),
	.shareout(Xd_0__inst_i19_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_30_48 (
// Equation(s):
// Xd_0__inst_mult_30_49  = SUM(( !Xd_0__inst_mult_30_4_q  $ (((!Xd_0__inst_mult_30_2_q ) # (!Xd_0__inst_mult_30_3_q ))) ) + ( Xd_0__inst_mult_30_98  ) + ( Xd_0__inst_mult_30_97  ))
// Xd_0__inst_mult_30_50  = CARRY(( !Xd_0__inst_mult_30_4_q  $ (((!Xd_0__inst_mult_30_2_q ) # (!Xd_0__inst_mult_30_3_q ))) ) + ( Xd_0__inst_mult_30_98  ) + ( Xd_0__inst_mult_30_97  ))
// Xd_0__inst_mult_30_51  = SHARE((Xd_0__inst_mult_30_2_q  & (Xd_0__inst_mult_30_3_q  & Xd_0__inst_mult_30_4_q )))

	.dataa(!Xd_0__inst_mult_30_2_q ),
	.datab(!Xd_0__inst_mult_30_3_q ),
	.datac(!Xd_0__inst_mult_30_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_97 ),
	.sharein(Xd_0__inst_mult_30_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_49 ),
	.cout(Xd_0__inst_mult_30_50 ),
	.shareout(Xd_0__inst_mult_30_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_31_48 (
// Equation(s):
// Xd_0__inst_mult_31_49  = SUM(( !Xd_0__inst_mult_31_4_q  $ (((!Xd_0__inst_mult_31_2_q ) # (!Xd_0__inst_mult_31_3_q ))) ) + ( Xd_0__inst_mult_31_98  ) + ( Xd_0__inst_mult_31_97  ))
// Xd_0__inst_mult_31_50  = CARRY(( !Xd_0__inst_mult_31_4_q  $ (((!Xd_0__inst_mult_31_2_q ) # (!Xd_0__inst_mult_31_3_q ))) ) + ( Xd_0__inst_mult_31_98  ) + ( Xd_0__inst_mult_31_97  ))
// Xd_0__inst_mult_31_51  = SHARE((Xd_0__inst_mult_31_2_q  & (Xd_0__inst_mult_31_3_q  & Xd_0__inst_mult_31_4_q )))

	.dataa(!Xd_0__inst_mult_31_2_q ),
	.datab(!Xd_0__inst_mult_31_3_q ),
	.datac(!Xd_0__inst_mult_31_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_97 ),
	.sharein(Xd_0__inst_mult_31_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_49 ),
	.cout(Xd_0__inst_mult_31_50 ),
	.shareout(Xd_0__inst_mult_31_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_30 (
// Equation(s):
// Xd_0__inst_mult_30_53  = SUM(( !Xd_0__inst_mult_30_5_q  $ (!Xd_0__inst_mult_30_6_q  $ (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_3_q )))) ) + ( Xd_0__inst_mult_30_51  ) + ( Xd_0__inst_mult_30_50  ))
// Xd_0__inst_mult_30_54  = CARRY(( !Xd_0__inst_mult_30_5_q  $ (!Xd_0__inst_mult_30_6_q  $ (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_3_q )))) ) + ( Xd_0__inst_mult_30_51  ) + ( Xd_0__inst_mult_30_50  ))
// Xd_0__inst_mult_30_55  = SHARE((!Xd_0__inst_mult_30_5_q  & (Xd_0__inst_mult_30_6_q  & (Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_3_q ))) # (Xd_0__inst_mult_30_5_q  & (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_3_q )) # (Xd_0__inst_mult_30_6_q ))))

	.dataa(!Xd_0__inst_mult_30_5_q ),
	.datab(!Xd_0__inst_mult_30_6_q ),
	.datac(!Xd_0__inst_mult_30_7_q ),
	.datad(!Xd_0__inst_mult_30_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_50 ),
	.sharein(Xd_0__inst_mult_30_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_53 ),
	.cout(Xd_0__inst_mult_30_54 ),
	.shareout(Xd_0__inst_mult_30_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_31 (
// Equation(s):
// Xd_0__inst_mult_31_53  = SUM(( !Xd_0__inst_mult_31_5_q  $ (!Xd_0__inst_mult_31_6_q  $ (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_3_q )))) ) + ( Xd_0__inst_mult_31_51  ) + ( Xd_0__inst_mult_31_50  ))
// Xd_0__inst_mult_31_54  = CARRY(( !Xd_0__inst_mult_31_5_q  $ (!Xd_0__inst_mult_31_6_q  $ (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_3_q )))) ) + ( Xd_0__inst_mult_31_51  ) + ( Xd_0__inst_mult_31_50  ))
// Xd_0__inst_mult_31_55  = SHARE((!Xd_0__inst_mult_31_5_q  & (Xd_0__inst_mult_31_6_q  & (Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_3_q ))) # (Xd_0__inst_mult_31_5_q  & (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_3_q )) # (Xd_0__inst_mult_31_6_q ))))

	.dataa(!Xd_0__inst_mult_31_5_q ),
	.datab(!Xd_0__inst_mult_31_6_q ),
	.datac(!Xd_0__inst_mult_31_7_q ),
	.datad(!Xd_0__inst_mult_31_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_50 ),
	.sharein(Xd_0__inst_mult_31_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_53 ),
	.cout(Xd_0__inst_mult_31_54 ),
	.shareout(Xd_0__inst_mult_31_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_30_21 (
// Equation(s):
// Xd_0__inst_mult_30_56  = SUM(( !Xd_0__inst_mult_30_8_q  $ (!Xd_0__inst_mult_30_9_q ) ) + ( Xd_0__inst_mult_30_55  ) + ( Xd_0__inst_mult_30_54  ))
// Xd_0__inst_mult_30_57  = CARRY(( !Xd_0__inst_mult_30_8_q  $ (!Xd_0__inst_mult_30_9_q ) ) + ( Xd_0__inst_mult_30_55  ) + ( Xd_0__inst_mult_30_54  ))
// Xd_0__inst_mult_30_58  = SHARE((Xd_0__inst_mult_30_8_q  & Xd_0__inst_mult_30_9_q ))

	.dataa(!Xd_0__inst_mult_30_8_q ),
	.datab(!Xd_0__inst_mult_30_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_54 ),
	.sharein(Xd_0__inst_mult_30_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_56 ),
	.cout(Xd_0__inst_mult_30_57 ),
	.shareout(Xd_0__inst_mult_30_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_31_21 (
// Equation(s):
// Xd_0__inst_mult_31_56  = SUM(( !Xd_0__inst_mult_31_8_q  $ (!Xd_0__inst_mult_31_9_q ) ) + ( Xd_0__inst_mult_31_55  ) + ( Xd_0__inst_mult_31_54  ))
// Xd_0__inst_mult_31_57  = CARRY(( !Xd_0__inst_mult_31_8_q  $ (!Xd_0__inst_mult_31_9_q ) ) + ( Xd_0__inst_mult_31_55  ) + ( Xd_0__inst_mult_31_54  ))
// Xd_0__inst_mult_31_58  = SHARE((Xd_0__inst_mult_31_8_q  & Xd_0__inst_mult_31_9_q ))

	.dataa(!Xd_0__inst_mult_31_8_q ),
	.datab(!Xd_0__inst_mult_31_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_54 ),
	.sharein(Xd_0__inst_mult_31_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_56 ),
	.cout(Xd_0__inst_mult_31_57 ),
	.shareout(Xd_0__inst_mult_31_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_30_22 (
// Equation(s):
// Xd_0__inst_mult_30_60  = SUM(( !Xd_0__inst_mult_30_10_q  $ (!Xd_0__inst_mult_30_11_q  $ (((Xd_0__inst_mult_30_2_q  & Xd_0__inst_mult_30_1_q )))) ) + ( Xd_0__inst_mult_30_58  ) + ( Xd_0__inst_mult_30_57  ))
// Xd_0__inst_mult_30_61  = CARRY(( !Xd_0__inst_mult_30_10_q  $ (!Xd_0__inst_mult_30_11_q  $ (((Xd_0__inst_mult_30_2_q  & Xd_0__inst_mult_30_1_q )))) ) + ( Xd_0__inst_mult_30_58  ) + ( Xd_0__inst_mult_30_57  ))
// Xd_0__inst_mult_30_62  = SHARE((!Xd_0__inst_mult_30_10_q  & (Xd_0__inst_mult_30_11_q  & (Xd_0__inst_mult_30_2_q  & Xd_0__inst_mult_30_1_q ))) # (Xd_0__inst_mult_30_10_q  & (((Xd_0__inst_mult_30_2_q  & Xd_0__inst_mult_30_1_q )) # (Xd_0__inst_mult_30_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_30_10_q ),
	.datab(!Xd_0__inst_mult_30_11_q ),
	.datac(!Xd_0__inst_mult_30_2_q ),
	.datad(!Xd_0__inst_mult_30_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_57 ),
	.sharein(Xd_0__inst_mult_30_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_60 ),
	.cout(Xd_0__inst_mult_30_61 ),
	.shareout(Xd_0__inst_mult_30_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_31_22 (
// Equation(s):
// Xd_0__inst_mult_31_60  = SUM(( !Xd_0__inst_mult_31_10_q  $ (!Xd_0__inst_mult_31_11_q  $ (((Xd_0__inst_mult_31_2_q  & Xd_0__inst_mult_31_1_q )))) ) + ( Xd_0__inst_mult_31_58  ) + ( Xd_0__inst_mult_31_57  ))
// Xd_0__inst_mult_31_61  = CARRY(( !Xd_0__inst_mult_31_10_q  $ (!Xd_0__inst_mult_31_11_q  $ (((Xd_0__inst_mult_31_2_q  & Xd_0__inst_mult_31_1_q )))) ) + ( Xd_0__inst_mult_31_58  ) + ( Xd_0__inst_mult_31_57  ))
// Xd_0__inst_mult_31_62  = SHARE((!Xd_0__inst_mult_31_10_q  & (Xd_0__inst_mult_31_11_q  & (Xd_0__inst_mult_31_2_q  & Xd_0__inst_mult_31_1_q ))) # (Xd_0__inst_mult_31_10_q  & (((Xd_0__inst_mult_31_2_q  & Xd_0__inst_mult_31_1_q )) # (Xd_0__inst_mult_31_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_31_10_q ),
	.datab(!Xd_0__inst_mult_31_11_q ),
	.datac(!Xd_0__inst_mult_31_2_q ),
	.datad(!Xd_0__inst_mult_31_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_57 ),
	.sharein(Xd_0__inst_mult_31_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_60 ),
	.cout(Xd_0__inst_mult_31_61 ),
	.shareout(Xd_0__inst_mult_31_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_30_23 (
// Equation(s):
// Xd_0__inst_mult_30_64  = SUM(( !Xd_0__inst_mult_30_12_q  $ (!Xd_0__inst_mult_30_13_q ) ) + ( Xd_0__inst_mult_30_62  ) + ( Xd_0__inst_mult_30_61  ))
// Xd_0__inst_mult_30_65  = CARRY(( !Xd_0__inst_mult_30_12_q  $ (!Xd_0__inst_mult_30_13_q ) ) + ( Xd_0__inst_mult_30_62  ) + ( Xd_0__inst_mult_30_61  ))
// Xd_0__inst_mult_30_66  = SHARE((Xd_0__inst_mult_30_12_q  & Xd_0__inst_mult_30_13_q ))

	.dataa(!Xd_0__inst_mult_30_12_q ),
	.datab(!Xd_0__inst_mult_30_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_61 ),
	.sharein(Xd_0__inst_mult_30_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_64 ),
	.cout(Xd_0__inst_mult_30_65 ),
	.shareout(Xd_0__inst_mult_30_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_31_23 (
// Equation(s):
// Xd_0__inst_mult_31_64  = SUM(( !Xd_0__inst_mult_31_12_q  $ (!Xd_0__inst_mult_31_13_q ) ) + ( Xd_0__inst_mult_31_62  ) + ( Xd_0__inst_mult_31_61  ))
// Xd_0__inst_mult_31_65  = CARRY(( !Xd_0__inst_mult_31_12_q  $ (!Xd_0__inst_mult_31_13_q ) ) + ( Xd_0__inst_mult_31_62  ) + ( Xd_0__inst_mult_31_61  ))
// Xd_0__inst_mult_31_66  = SHARE((Xd_0__inst_mult_31_12_q  & Xd_0__inst_mult_31_13_q ))

	.dataa(!Xd_0__inst_mult_31_12_q ),
	.datab(!Xd_0__inst_mult_31_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_61 ),
	.sharein(Xd_0__inst_mult_31_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_64 ),
	.cout(Xd_0__inst_mult_31_65 ),
	.shareout(Xd_0__inst_mult_31_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_30_24 (
// Equation(s):
// Xd_0__inst_mult_30_68  = SUM(( !Xd_0__inst_mult_30_14_q  $ (!Xd_0__inst_mult_30_15_q ) ) + ( Xd_0__inst_mult_30_66  ) + ( Xd_0__inst_mult_30_65  ))
// Xd_0__inst_mult_30_69  = CARRY(( !Xd_0__inst_mult_30_14_q  $ (!Xd_0__inst_mult_30_15_q ) ) + ( Xd_0__inst_mult_30_66  ) + ( Xd_0__inst_mult_30_65  ))
// Xd_0__inst_mult_30_70  = SHARE((Xd_0__inst_mult_30_14_q  & Xd_0__inst_mult_30_15_q ))

	.dataa(!Xd_0__inst_mult_30_14_q ),
	.datab(!Xd_0__inst_mult_30_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_65 ),
	.sharein(Xd_0__inst_mult_30_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_68 ),
	.cout(Xd_0__inst_mult_30_69 ),
	.shareout(Xd_0__inst_mult_30_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_31_24 (
// Equation(s):
// Xd_0__inst_mult_31_68  = SUM(( !Xd_0__inst_mult_31_14_q  $ (!Xd_0__inst_mult_31_15_q ) ) + ( Xd_0__inst_mult_31_66  ) + ( Xd_0__inst_mult_31_65  ))
// Xd_0__inst_mult_31_69  = CARRY(( !Xd_0__inst_mult_31_14_q  $ (!Xd_0__inst_mult_31_15_q ) ) + ( Xd_0__inst_mult_31_66  ) + ( Xd_0__inst_mult_31_65  ))
// Xd_0__inst_mult_31_70  = SHARE((Xd_0__inst_mult_31_14_q  & Xd_0__inst_mult_31_15_q ))

	.dataa(!Xd_0__inst_mult_31_14_q ),
	.datab(!Xd_0__inst_mult_31_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_65 ),
	.sharein(Xd_0__inst_mult_31_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_68 ),
	.cout(Xd_0__inst_mult_31_69 ),
	.shareout(Xd_0__inst_mult_31_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_30_25 (
// Equation(s):
// Xd_0__inst_mult_30_72  = SUM(( !Xd_0__inst_mult_30_16_q  $ (!Xd_0__inst_mult_30_17_q  $ (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_18_q )))) ) + ( Xd_0__inst_mult_30_70  ) + ( Xd_0__inst_mult_30_69  ))
// Xd_0__inst_mult_30_73  = CARRY(( !Xd_0__inst_mult_30_16_q  $ (!Xd_0__inst_mult_30_17_q  $ (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_18_q )))) ) + ( Xd_0__inst_mult_30_70  ) + ( Xd_0__inst_mult_30_69  ))
// Xd_0__inst_mult_30_74  = SHARE((!Xd_0__inst_mult_30_16_q  & (Xd_0__inst_mult_30_17_q  & (Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_18_q ))) # (Xd_0__inst_mult_30_16_q  & (((Xd_0__inst_mult_30_7_q  & Xd_0__inst_mult_30_18_q )) # (Xd_0__inst_mult_30_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_30_16_q ),
	.datab(!Xd_0__inst_mult_30_17_q ),
	.datac(!Xd_0__inst_mult_30_7_q ),
	.datad(!Xd_0__inst_mult_30_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_69 ),
	.sharein(Xd_0__inst_mult_30_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_72 ),
	.cout(Xd_0__inst_mult_30_73 ),
	.shareout(Xd_0__inst_mult_30_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_31_25 (
// Equation(s):
// Xd_0__inst_mult_31_72  = SUM(( !Xd_0__inst_mult_31_16_q  $ (!Xd_0__inst_mult_31_17_q  $ (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_18_q )))) ) + ( Xd_0__inst_mult_31_70  ) + ( Xd_0__inst_mult_31_69  ))
// Xd_0__inst_mult_31_73  = CARRY(( !Xd_0__inst_mult_31_16_q  $ (!Xd_0__inst_mult_31_17_q  $ (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_18_q )))) ) + ( Xd_0__inst_mult_31_70  ) + ( Xd_0__inst_mult_31_69  ))
// Xd_0__inst_mult_31_74  = SHARE((!Xd_0__inst_mult_31_16_q  & (Xd_0__inst_mult_31_17_q  & (Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_18_q ))) # (Xd_0__inst_mult_31_16_q  & (((Xd_0__inst_mult_31_7_q  & Xd_0__inst_mult_31_18_q )) # (Xd_0__inst_mult_31_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_31_16_q ),
	.datab(!Xd_0__inst_mult_31_17_q ),
	.datac(!Xd_0__inst_mult_31_7_q ),
	.datad(!Xd_0__inst_mult_31_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_69 ),
	.sharein(Xd_0__inst_mult_31_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_72 ),
	.cout(Xd_0__inst_mult_31_73 ),
	.shareout(Xd_0__inst_mult_31_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_30_26 (
// Equation(s):
// Xd_0__inst_mult_30_76  = SUM(( !Xd_0__inst_mult_30_20_q  $ (((!Xd_0__inst_mult_30_19_q ) # (!Xd_0__inst_mult_30_18_q ))) ) + ( Xd_0__inst_mult_30_74  ) + ( Xd_0__inst_mult_30_73  ))
// Xd_0__inst_mult_30_77  = CARRY(( !Xd_0__inst_mult_30_20_q  $ (((!Xd_0__inst_mult_30_19_q ) # (!Xd_0__inst_mult_30_18_q ))) ) + ( Xd_0__inst_mult_30_74  ) + ( Xd_0__inst_mult_30_73  ))
// Xd_0__inst_mult_30_78  = SHARE((Xd_0__inst_mult_30_19_q  & (Xd_0__inst_mult_30_18_q  & Xd_0__inst_mult_30_20_q )))

	.dataa(!Xd_0__inst_mult_30_19_q ),
	.datab(!Xd_0__inst_mult_30_18_q ),
	.datac(!Xd_0__inst_mult_30_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_73 ),
	.sharein(Xd_0__inst_mult_30_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_76 ),
	.cout(Xd_0__inst_mult_30_77 ),
	.shareout(Xd_0__inst_mult_30_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_31_26 (
// Equation(s):
// Xd_0__inst_mult_31_76  = SUM(( !Xd_0__inst_mult_31_20_q  $ (((!Xd_0__inst_mult_31_19_q ) # (!Xd_0__inst_mult_31_18_q ))) ) + ( Xd_0__inst_mult_31_74  ) + ( Xd_0__inst_mult_31_73  ))
// Xd_0__inst_mult_31_77  = CARRY(( !Xd_0__inst_mult_31_20_q  $ (((!Xd_0__inst_mult_31_19_q ) # (!Xd_0__inst_mult_31_18_q ))) ) + ( Xd_0__inst_mult_31_74  ) + ( Xd_0__inst_mult_31_73  ))
// Xd_0__inst_mult_31_78  = SHARE((Xd_0__inst_mult_31_19_q  & (Xd_0__inst_mult_31_18_q  & Xd_0__inst_mult_31_20_q )))

	.dataa(!Xd_0__inst_mult_31_19_q ),
	.datab(!Xd_0__inst_mult_31_18_q ),
	.datac(!Xd_0__inst_mult_31_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_73 ),
	.sharein(Xd_0__inst_mult_31_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_76 ),
	.cout(Xd_0__inst_mult_31_77 ),
	.shareout(Xd_0__inst_mult_31_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_27 (
// Equation(s):
// Xd_0__inst_mult_30_80  = SUM(( GND ) + ( Xd_0__inst_mult_30_78  ) + ( Xd_0__inst_mult_30_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_77 ),
	.sharein(Xd_0__inst_mult_30_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_27 (
// Equation(s):
// Xd_0__inst_mult_31_80  = SUM(( GND ) + ( Xd_0__inst_mult_31_78  ) + ( Xd_0__inst_mult_31_77  ))
// Xd_0__inst_mult_31_81  = CARRY(( GND ) + ( Xd_0__inst_mult_31_78  ) + ( Xd_0__inst_mult_31_77  ))
// Xd_0__inst_mult_31_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_77 ),
	.sharein(Xd_0__inst_mult_31_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_80 ),
	.cout(Xd_0__inst_mult_31_81 ),
	.shareout(Xd_0__inst_mult_31_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_89 (
// Equation(s):
// Xd_0__inst_i19_89_sumout  = SUM(( !din_a[181] $ (!din_b[181]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_90  = CARRY(( !din_a[181] $ (!din_b[181]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_91  = SHARE(GND)

	.dataa(!din_a[181]),
	.datab(!din_b[181]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_89_sumout ),
	.cout(Xd_0__inst_i19_90 ),
	.shareout(Xd_0__inst_i19_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_93 (
// Equation(s):
// Xd_0__inst_i19_93_sumout  = SUM(( !din_a[153] $ (!din_b[153]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_94  = CARRY(( !din_a[153] $ (!din_b[153]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_95  = SHARE(GND)

	.dataa(!din_a[153]),
	.datab(!din_b[153]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_93_sumout ),
	.cout(Xd_0__inst_i19_94 ),
	.shareout(Xd_0__inst_i19_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_28 (
// Equation(s):
// Xd_0__inst_mult_30_84  = SUM(( (din_a[210] & din_b[210]) ) + ( Xd_0__inst_mult_25_90  ) + ( Xd_0__inst_mult_25_89  ))
// Xd_0__inst_mult_30_85  = CARRY(( (din_a[210] & din_b[210]) ) + ( Xd_0__inst_mult_25_90  ) + ( Xd_0__inst_mult_25_89  ))
// Xd_0__inst_mult_30_86  = SHARE((din_a[210] & din_b[211]))

	.dataa(!din_a[210]),
	.datab(!din_b[210]),
	.datac(!din_b[211]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_89 ),
	.sharein(Xd_0__inst_mult_25_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_84 ),
	.cout(Xd_0__inst_mult_30_85 ),
	.shareout(Xd_0__inst_mult_30_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_28 (
// Equation(s):
// Xd_0__inst_mult_31_84  = SUM(( (din_a[217] & din_b[217]) ) + ( Xd_0__inst_mult_22_90  ) + ( Xd_0__inst_mult_22_89  ))
// Xd_0__inst_mult_31_85  = CARRY(( (din_a[217] & din_b[217]) ) + ( Xd_0__inst_mult_22_90  ) + ( Xd_0__inst_mult_22_89  ))
// Xd_0__inst_mult_31_86  = SHARE((din_a[217] & din_b[218]))

	.dataa(!din_a[217]),
	.datab(!din_b[217]),
	.datac(!din_b[218]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_89 ),
	.sharein(Xd_0__inst_mult_22_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_84 ),
	.cout(Xd_0__inst_mult_31_85 ),
	.shareout(Xd_0__inst_mult_31_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_97 (
// Equation(s):
// Xd_0__inst_i19_97_sumout  = SUM(( !din_a[13] $ (!din_b[13]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_98  = CARRY(( !din_a[13] $ (!din_b[13]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_99  = SHARE(GND)

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_97_sumout ),
	.cout(Xd_0__inst_i19_98 ),
	.shareout(Xd_0__inst_i19_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_101 (
// Equation(s):
// Xd_0__inst_i19_101_sumout  = SUM(( !din_a[97] $ (!din_b[97]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_102  = CARRY(( !din_a[97] $ (!din_b[97]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_103  = SHARE(GND)

	.dataa(!din_a[97]),
	.datab(!din_b[97]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_101_sumout ),
	.cout(Xd_0__inst_i19_102 ),
	.shareout(Xd_0__inst_i19_103 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_105 (
// Equation(s):
// Xd_0__inst_i19_105_sumout  = SUM(( !din_a[55] $ (!din_b[55]) ) + ( Xd_0__inst_i19_115  ) + ( Xd_0__inst_i19_114  ))
// Xd_0__inst_i19_106  = CARRY(( !din_a[55] $ (!din_b[55]) ) + ( Xd_0__inst_i19_115  ) + ( Xd_0__inst_i19_114  ))
// Xd_0__inst_i19_107  = SHARE(GND)

	.dataa(!din_a[55]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_114 ),
	.sharein(Xd_0__inst_i19_115 ),
	.combout(),
	.sumout(Xd_0__inst_i19_105_sumout ),
	.cout(Xd_0__inst_i19_106 ),
	.shareout(Xd_0__inst_i19_107 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_109 (
// Equation(s):
// Xd_0__inst_i19_109_sumout  = SUM(( !din_a[69] $ (!din_b[69]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_110  = CARRY(( !din_a[69] $ (!din_b[69]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_111  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_109_sumout ),
	.cout(Xd_0__inst_i19_110 ),
	.shareout(Xd_0__inst_i19_111 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_29 (
// Equation(s):
// Xd_0__inst_mult_30_88  = SUM(( (din_a[211] & din_b[210]) ) + ( Xd_0__inst_mult_30_86  ) + ( Xd_0__inst_mult_30_85  ))
// Xd_0__inst_mult_30_89  = CARRY(( (din_a[211] & din_b[210]) ) + ( Xd_0__inst_mult_30_86  ) + ( Xd_0__inst_mult_30_85  ))
// Xd_0__inst_mult_30_90  = SHARE((din_a[210] & din_b[212]))

	.dataa(!din_a[211]),
	.datab(!din_b[210]),
	.datac(!din_a[210]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_85 ),
	.sharein(Xd_0__inst_mult_30_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_88 ),
	.cout(Xd_0__inst_mult_30_89 ),
	.shareout(Xd_0__inst_mult_30_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_29 (
// Equation(s):
// Xd_0__inst_mult_31_88  = SUM(( (din_a[218] & din_b[217]) ) + ( Xd_0__inst_mult_31_86  ) + ( Xd_0__inst_mult_31_85  ))
// Xd_0__inst_mult_31_89  = CARRY(( (din_a[218] & din_b[217]) ) + ( Xd_0__inst_mult_31_86  ) + ( Xd_0__inst_mult_31_85  ))
// Xd_0__inst_mult_31_90  = SHARE((din_a[217] & din_b[219]))

	.dataa(!din_a[218]),
	.datab(!din_b[217]),
	.datac(!din_a[217]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_85 ),
	.sharein(Xd_0__inst_mult_31_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_88 ),
	.cout(Xd_0__inst_mult_31_89 ),
	.shareout(Xd_0__inst_mult_31_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_30 (
// Equation(s):
// Xd_0__inst_mult_30_92  = SUM(( (!din_a[211] & (((din_a[212] & din_b[210])))) # (din_a[211] & (!din_b[211] $ (((!din_a[212]) # (!din_b[210]))))) ) + ( Xd_0__inst_mult_30_90  ) + ( Xd_0__inst_mult_30_89  ))
// Xd_0__inst_mult_30_93  = CARRY(( (!din_a[211] & (((din_a[212] & din_b[210])))) # (din_a[211] & (!din_b[211] $ (((!din_a[212]) # (!din_b[210]))))) ) + ( Xd_0__inst_mult_30_90  ) + ( Xd_0__inst_mult_30_89  ))
// Xd_0__inst_mult_30_94  = SHARE((din_a[211] & (din_b[211] & (din_a[212] & din_b[210]))))

	.dataa(!din_a[211]),
	.datab(!din_b[211]),
	.datac(!din_a[212]),
	.datad(!din_b[210]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_89 ),
	.sharein(Xd_0__inst_mult_30_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_92 ),
	.cout(Xd_0__inst_mult_30_93 ),
	.shareout(Xd_0__inst_mult_30_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_30 (
// Equation(s):
// Xd_0__inst_mult_31_92  = SUM(( (!din_a[218] & (((din_a[219] & din_b[217])))) # (din_a[218] & (!din_b[218] $ (((!din_a[219]) # (!din_b[217]))))) ) + ( Xd_0__inst_mult_31_90  ) + ( Xd_0__inst_mult_31_89  ))
// Xd_0__inst_mult_31_93  = CARRY(( (!din_a[218] & (((din_a[219] & din_b[217])))) # (din_a[218] & (!din_b[218] $ (((!din_a[219]) # (!din_b[217]))))) ) + ( Xd_0__inst_mult_31_90  ) + ( Xd_0__inst_mult_31_89  ))
// Xd_0__inst_mult_31_94  = SHARE((din_a[218] & (din_b[218] & (din_a[219] & din_b[217]))))

	.dataa(!din_a[218]),
	.datab(!din_b[218]),
	.datac(!din_a[219]),
	.datad(!din_b[217]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_89 ),
	.sharein(Xd_0__inst_mult_31_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_92 ),
	.cout(Xd_0__inst_mult_31_93 ),
	.shareout(Xd_0__inst_mult_31_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_28_48 (
// Equation(s):
// Xd_0__inst_mult_28_49  = SUM(( !Xd_0__inst_mult_28_4_q  $ (((!Xd_0__inst_mult_28_2_q ) # (!Xd_0__inst_mult_28_3_q ))) ) + ( Xd_0__inst_mult_28_98  ) + ( Xd_0__inst_mult_28_97  ))
// Xd_0__inst_mult_28_50  = CARRY(( !Xd_0__inst_mult_28_4_q  $ (((!Xd_0__inst_mult_28_2_q ) # (!Xd_0__inst_mult_28_3_q ))) ) + ( Xd_0__inst_mult_28_98  ) + ( Xd_0__inst_mult_28_97  ))
// Xd_0__inst_mult_28_51  = SHARE((Xd_0__inst_mult_28_2_q  & (Xd_0__inst_mult_28_3_q  & Xd_0__inst_mult_28_4_q )))

	.dataa(!Xd_0__inst_mult_28_2_q ),
	.datab(!Xd_0__inst_mult_28_3_q ),
	.datac(!Xd_0__inst_mult_28_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_97 ),
	.sharein(Xd_0__inst_mult_28_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_49 ),
	.cout(Xd_0__inst_mult_28_50 ),
	.shareout(Xd_0__inst_mult_28_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_29_48 (
// Equation(s):
// Xd_0__inst_mult_29_49  = SUM(( !Xd_0__inst_mult_29_4_q  $ (((!Xd_0__inst_mult_29_2_q ) # (!Xd_0__inst_mult_29_3_q ))) ) + ( Xd_0__inst_mult_29_98  ) + ( Xd_0__inst_mult_29_97  ))
// Xd_0__inst_mult_29_50  = CARRY(( !Xd_0__inst_mult_29_4_q  $ (((!Xd_0__inst_mult_29_2_q ) # (!Xd_0__inst_mult_29_3_q ))) ) + ( Xd_0__inst_mult_29_98  ) + ( Xd_0__inst_mult_29_97  ))
// Xd_0__inst_mult_29_51  = SHARE((Xd_0__inst_mult_29_2_q  & (Xd_0__inst_mult_29_3_q  & Xd_0__inst_mult_29_4_q )))

	.dataa(!Xd_0__inst_mult_29_2_q ),
	.datab(!Xd_0__inst_mult_29_3_q ),
	.datac(!Xd_0__inst_mult_29_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_97 ),
	.sharein(Xd_0__inst_mult_29_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_49 ),
	.cout(Xd_0__inst_mult_29_50 ),
	.shareout(Xd_0__inst_mult_29_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_26_48 (
// Equation(s):
// Xd_0__inst_mult_26_49  = SUM(( !Xd_0__inst_mult_26_4_q  $ (((!Xd_0__inst_mult_26_2_q ) # (!Xd_0__inst_mult_26_3_q ))) ) + ( Xd_0__inst_mult_26_98  ) + ( Xd_0__inst_mult_26_97  ))
// Xd_0__inst_mult_26_50  = CARRY(( !Xd_0__inst_mult_26_4_q  $ (((!Xd_0__inst_mult_26_2_q ) # (!Xd_0__inst_mult_26_3_q ))) ) + ( Xd_0__inst_mult_26_98  ) + ( Xd_0__inst_mult_26_97  ))
// Xd_0__inst_mult_26_51  = SHARE((Xd_0__inst_mult_26_2_q  & (Xd_0__inst_mult_26_3_q  & Xd_0__inst_mult_26_4_q )))

	.dataa(!Xd_0__inst_mult_26_2_q ),
	.datab(!Xd_0__inst_mult_26_3_q ),
	.datac(!Xd_0__inst_mult_26_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_97 ),
	.sharein(Xd_0__inst_mult_26_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_49 ),
	.cout(Xd_0__inst_mult_26_50 ),
	.shareout(Xd_0__inst_mult_26_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_27_48 (
// Equation(s):
// Xd_0__inst_mult_27_49  = SUM(( !Xd_0__inst_mult_27_4_q  $ (((!Xd_0__inst_mult_27_2_q ) # (!Xd_0__inst_mult_27_3_q ))) ) + ( Xd_0__inst_mult_27_98  ) + ( Xd_0__inst_mult_27_97  ))
// Xd_0__inst_mult_27_50  = CARRY(( !Xd_0__inst_mult_27_4_q  $ (((!Xd_0__inst_mult_27_2_q ) # (!Xd_0__inst_mult_27_3_q ))) ) + ( Xd_0__inst_mult_27_98  ) + ( Xd_0__inst_mult_27_97  ))
// Xd_0__inst_mult_27_51  = SHARE((Xd_0__inst_mult_27_2_q  & (Xd_0__inst_mult_27_3_q  & Xd_0__inst_mult_27_4_q )))

	.dataa(!Xd_0__inst_mult_27_2_q ),
	.datab(!Xd_0__inst_mult_27_3_q ),
	.datac(!Xd_0__inst_mult_27_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_97 ),
	.sharein(Xd_0__inst_mult_27_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_49 ),
	.cout(Xd_0__inst_mult_27_50 ),
	.shareout(Xd_0__inst_mult_27_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_24_48 (
// Equation(s):
// Xd_0__inst_mult_24_49  = SUM(( !Xd_0__inst_mult_24_4_q  $ (((!Xd_0__inst_mult_24_2_q ) # (!Xd_0__inst_mult_24_3_q ))) ) + ( Xd_0__inst_mult_24_98  ) + ( Xd_0__inst_mult_24_97  ))
// Xd_0__inst_mult_24_50  = CARRY(( !Xd_0__inst_mult_24_4_q  $ (((!Xd_0__inst_mult_24_2_q ) # (!Xd_0__inst_mult_24_3_q ))) ) + ( Xd_0__inst_mult_24_98  ) + ( Xd_0__inst_mult_24_97  ))
// Xd_0__inst_mult_24_51  = SHARE((Xd_0__inst_mult_24_2_q  & (Xd_0__inst_mult_24_3_q  & Xd_0__inst_mult_24_4_q )))

	.dataa(!Xd_0__inst_mult_24_2_q ),
	.datab(!Xd_0__inst_mult_24_3_q ),
	.datac(!Xd_0__inst_mult_24_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_97 ),
	.sharein(Xd_0__inst_mult_24_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_49 ),
	.cout(Xd_0__inst_mult_24_50 ),
	.shareout(Xd_0__inst_mult_24_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_25_48 (
// Equation(s):
// Xd_0__inst_mult_25_49  = SUM(( !Xd_0__inst_mult_25_4_q  $ (((!Xd_0__inst_mult_25_2_q ) # (!Xd_0__inst_mult_25_3_q ))) ) + ( Xd_0__inst_mult_25_102  ) + ( Xd_0__inst_mult_25_101  ))
// Xd_0__inst_mult_25_50  = CARRY(( !Xd_0__inst_mult_25_4_q  $ (((!Xd_0__inst_mult_25_2_q ) # (!Xd_0__inst_mult_25_3_q ))) ) + ( Xd_0__inst_mult_25_102  ) + ( Xd_0__inst_mult_25_101  ))
// Xd_0__inst_mult_25_51  = SHARE((Xd_0__inst_mult_25_2_q  & (Xd_0__inst_mult_25_3_q  & Xd_0__inst_mult_25_4_q )))

	.dataa(!Xd_0__inst_mult_25_2_q ),
	.datab(!Xd_0__inst_mult_25_3_q ),
	.datac(!Xd_0__inst_mult_25_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_101 ),
	.sharein(Xd_0__inst_mult_25_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_49 ),
	.cout(Xd_0__inst_mult_25_50 ),
	.shareout(Xd_0__inst_mult_25_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_22_48 (
// Equation(s):
// Xd_0__inst_mult_22_49  = SUM(( !Xd_0__inst_mult_22_4_q  $ (((!Xd_0__inst_mult_22_2_q ) # (!Xd_0__inst_mult_22_3_q ))) ) + ( Xd_0__inst_mult_22_102  ) + ( Xd_0__inst_mult_22_101  ))
// Xd_0__inst_mult_22_50  = CARRY(( !Xd_0__inst_mult_22_4_q  $ (((!Xd_0__inst_mult_22_2_q ) # (!Xd_0__inst_mult_22_3_q ))) ) + ( Xd_0__inst_mult_22_102  ) + ( Xd_0__inst_mult_22_101  ))
// Xd_0__inst_mult_22_51  = SHARE((Xd_0__inst_mult_22_2_q  & (Xd_0__inst_mult_22_3_q  & Xd_0__inst_mult_22_4_q )))

	.dataa(!Xd_0__inst_mult_22_2_q ),
	.datab(!Xd_0__inst_mult_22_3_q ),
	.datac(!Xd_0__inst_mult_22_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_101 ),
	.sharein(Xd_0__inst_mult_22_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_49 ),
	.cout(Xd_0__inst_mult_22_50 ),
	.shareout(Xd_0__inst_mult_22_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_23_48 (
// Equation(s):
// Xd_0__inst_mult_23_49  = SUM(( !Xd_0__inst_mult_23_4_q  $ (((!Xd_0__inst_mult_23_2_q ) # (!Xd_0__inst_mult_23_3_q ))) ) + ( Xd_0__inst_mult_23_98  ) + ( Xd_0__inst_mult_23_97  ))
// Xd_0__inst_mult_23_50  = CARRY(( !Xd_0__inst_mult_23_4_q  $ (((!Xd_0__inst_mult_23_2_q ) # (!Xd_0__inst_mult_23_3_q ))) ) + ( Xd_0__inst_mult_23_98  ) + ( Xd_0__inst_mult_23_97  ))
// Xd_0__inst_mult_23_51  = SHARE((Xd_0__inst_mult_23_2_q  & (Xd_0__inst_mult_23_3_q  & Xd_0__inst_mult_23_4_q )))

	.dataa(!Xd_0__inst_mult_23_2_q ),
	.datab(!Xd_0__inst_mult_23_3_q ),
	.datac(!Xd_0__inst_mult_23_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_97 ),
	.sharein(Xd_0__inst_mult_23_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_49 ),
	.cout(Xd_0__inst_mult_23_50 ),
	.shareout(Xd_0__inst_mult_23_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_20_48 (
// Equation(s):
// Xd_0__inst_mult_20_49  = SUM(( !Xd_0__inst_mult_20_4_q  $ (((!Xd_0__inst_mult_20_2_q ) # (!Xd_0__inst_mult_20_3_q ))) ) + ( Xd_0__inst_mult_20_98  ) + ( Xd_0__inst_mult_20_97  ))
// Xd_0__inst_mult_20_50  = CARRY(( !Xd_0__inst_mult_20_4_q  $ (((!Xd_0__inst_mult_20_2_q ) # (!Xd_0__inst_mult_20_3_q ))) ) + ( Xd_0__inst_mult_20_98  ) + ( Xd_0__inst_mult_20_97  ))
// Xd_0__inst_mult_20_51  = SHARE((Xd_0__inst_mult_20_2_q  & (Xd_0__inst_mult_20_3_q  & Xd_0__inst_mult_20_4_q )))

	.dataa(!Xd_0__inst_mult_20_2_q ),
	.datab(!Xd_0__inst_mult_20_3_q ),
	.datac(!Xd_0__inst_mult_20_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_97 ),
	.sharein(Xd_0__inst_mult_20_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_49 ),
	.cout(Xd_0__inst_mult_20_50 ),
	.shareout(Xd_0__inst_mult_20_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_21_48 (
// Equation(s):
// Xd_0__inst_mult_21_49  = SUM(( !Xd_0__inst_mult_21_4_q  $ (((!Xd_0__inst_mult_21_2_q ) # (!Xd_0__inst_mult_21_3_q ))) ) + ( Xd_0__inst_mult_21_98  ) + ( Xd_0__inst_mult_21_97  ))
// Xd_0__inst_mult_21_50  = CARRY(( !Xd_0__inst_mult_21_4_q  $ (((!Xd_0__inst_mult_21_2_q ) # (!Xd_0__inst_mult_21_3_q ))) ) + ( Xd_0__inst_mult_21_98  ) + ( Xd_0__inst_mult_21_97  ))
// Xd_0__inst_mult_21_51  = SHARE((Xd_0__inst_mult_21_2_q  & (Xd_0__inst_mult_21_3_q  & Xd_0__inst_mult_21_4_q )))

	.dataa(!Xd_0__inst_mult_21_2_q ),
	.datab(!Xd_0__inst_mult_21_3_q ),
	.datac(!Xd_0__inst_mult_21_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_97 ),
	.sharein(Xd_0__inst_mult_21_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_49 ),
	.cout(Xd_0__inst_mult_21_50 ),
	.shareout(Xd_0__inst_mult_21_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_18_48 (
// Equation(s):
// Xd_0__inst_mult_18_49  = SUM(( !Xd_0__inst_mult_18_4_q  $ (((!Xd_0__inst_mult_18_2_q ) # (!Xd_0__inst_mult_18_3_q ))) ) + ( Xd_0__inst_mult_18_98  ) + ( Xd_0__inst_mult_18_97  ))
// Xd_0__inst_mult_18_50  = CARRY(( !Xd_0__inst_mult_18_4_q  $ (((!Xd_0__inst_mult_18_2_q ) # (!Xd_0__inst_mult_18_3_q ))) ) + ( Xd_0__inst_mult_18_98  ) + ( Xd_0__inst_mult_18_97  ))
// Xd_0__inst_mult_18_51  = SHARE((Xd_0__inst_mult_18_2_q  & (Xd_0__inst_mult_18_3_q  & Xd_0__inst_mult_18_4_q )))

	.dataa(!Xd_0__inst_mult_18_2_q ),
	.datab(!Xd_0__inst_mult_18_3_q ),
	.datac(!Xd_0__inst_mult_18_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_97 ),
	.sharein(Xd_0__inst_mult_18_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_49 ),
	.cout(Xd_0__inst_mult_18_50 ),
	.shareout(Xd_0__inst_mult_18_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_19_48 (
// Equation(s):
// Xd_0__inst_mult_19_49  = SUM(( !Xd_0__inst_mult_19_4_q  $ (((!Xd_0__inst_mult_19_2_q ) # (!Xd_0__inst_mult_19_3_q ))) ) + ( Xd_0__inst_mult_19_98  ) + ( Xd_0__inst_mult_19_97  ))
// Xd_0__inst_mult_19_50  = CARRY(( !Xd_0__inst_mult_19_4_q  $ (((!Xd_0__inst_mult_19_2_q ) # (!Xd_0__inst_mult_19_3_q ))) ) + ( Xd_0__inst_mult_19_98  ) + ( Xd_0__inst_mult_19_97  ))
// Xd_0__inst_mult_19_51  = SHARE((Xd_0__inst_mult_19_2_q  & (Xd_0__inst_mult_19_3_q  & Xd_0__inst_mult_19_4_q )))

	.dataa(!Xd_0__inst_mult_19_2_q ),
	.datab(!Xd_0__inst_mult_19_3_q ),
	.datac(!Xd_0__inst_mult_19_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_97 ),
	.sharein(Xd_0__inst_mult_19_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_49 ),
	.cout(Xd_0__inst_mult_19_50 ),
	.shareout(Xd_0__inst_mult_19_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_31 (
// Equation(s):
// Xd_0__inst_mult_30_97  = CARRY(( GND ) + ( Xd_0__inst_mult_31_82  ) + ( Xd_0__inst_mult_31_81  ))
// Xd_0__inst_mult_30_98  = SHARE((Xd_0__inst_mult_30_0_q  & Xd_0__inst_mult_30_1_q ))

	.dataa(!Xd_0__inst_mult_30_0_q ),
	.datab(!Xd_0__inst_mult_30_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_81 ),
	.sharein(Xd_0__inst_mult_31_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_97 ),
	.shareout(Xd_0__inst_mult_30_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_31 (
// Equation(s):
// Xd_0__inst_mult_31_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_31_98  = SHARE((Xd_0__inst_mult_31_0_q  & Xd_0__inst_mult_31_1_q ))

	.dataa(!Xd_0__inst_mult_31_0_q ),
	.datab(!Xd_0__inst_mult_31_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_97 ),
	.shareout(Xd_0__inst_mult_31_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_16_48 (
// Equation(s):
// Xd_0__inst_mult_16_49  = SUM(( !Xd_0__inst_mult_16_4_q  $ (((!Xd_0__inst_mult_16_2_q ) # (!Xd_0__inst_mult_16_3_q ))) ) + ( Xd_0__inst_mult_16_98  ) + ( Xd_0__inst_mult_16_97  ))
// Xd_0__inst_mult_16_50  = CARRY(( !Xd_0__inst_mult_16_4_q  $ (((!Xd_0__inst_mult_16_2_q ) # (!Xd_0__inst_mult_16_3_q ))) ) + ( Xd_0__inst_mult_16_98  ) + ( Xd_0__inst_mult_16_97  ))
// Xd_0__inst_mult_16_51  = SHARE((Xd_0__inst_mult_16_2_q  & (Xd_0__inst_mult_16_3_q  & Xd_0__inst_mult_16_4_q )))

	.dataa(!Xd_0__inst_mult_16_2_q ),
	.datab(!Xd_0__inst_mult_16_3_q ),
	.datac(!Xd_0__inst_mult_16_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_97 ),
	.sharein(Xd_0__inst_mult_16_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_49 ),
	.cout(Xd_0__inst_mult_16_50 ),
	.shareout(Xd_0__inst_mult_16_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_17_48 (
// Equation(s):
// Xd_0__inst_mult_17_49  = SUM(( !Xd_0__inst_mult_17_4_q  $ (((!Xd_0__inst_mult_17_2_q ) # (!Xd_0__inst_mult_17_3_q ))) ) + ( Xd_0__inst_mult_17_98  ) + ( Xd_0__inst_mult_17_97  ))
// Xd_0__inst_mult_17_50  = CARRY(( !Xd_0__inst_mult_17_4_q  $ (((!Xd_0__inst_mult_17_2_q ) # (!Xd_0__inst_mult_17_3_q ))) ) + ( Xd_0__inst_mult_17_98  ) + ( Xd_0__inst_mult_17_97  ))
// Xd_0__inst_mult_17_51  = SHARE((Xd_0__inst_mult_17_2_q  & (Xd_0__inst_mult_17_3_q  & Xd_0__inst_mult_17_4_q )))

	.dataa(!Xd_0__inst_mult_17_2_q ),
	.datab(!Xd_0__inst_mult_17_3_q ),
	.datac(!Xd_0__inst_mult_17_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_97 ),
	.sharein(Xd_0__inst_mult_17_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_49 ),
	.cout(Xd_0__inst_mult_17_50 ),
	.shareout(Xd_0__inst_mult_17_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_48 (
// Equation(s):
// Xd_0__inst_mult_14_49  = SUM(( !Xd_0__inst_mult_14_4_q  $ (((!Xd_0__inst_mult_14_2_q ) # (!Xd_0__inst_mult_14_3_q ))) ) + ( Xd_0__inst_mult_14_98  ) + ( Xd_0__inst_mult_14_97  ))
// Xd_0__inst_mult_14_50  = CARRY(( !Xd_0__inst_mult_14_4_q  $ (((!Xd_0__inst_mult_14_2_q ) # (!Xd_0__inst_mult_14_3_q ))) ) + ( Xd_0__inst_mult_14_98  ) + ( Xd_0__inst_mult_14_97  ))
// Xd_0__inst_mult_14_51  = SHARE((Xd_0__inst_mult_14_2_q  & (Xd_0__inst_mult_14_3_q  & Xd_0__inst_mult_14_4_q )))

	.dataa(!Xd_0__inst_mult_14_2_q ),
	.datab(!Xd_0__inst_mult_14_3_q ),
	.datac(!Xd_0__inst_mult_14_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_97 ),
	.sharein(Xd_0__inst_mult_14_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_49 ),
	.cout(Xd_0__inst_mult_14_50 ),
	.shareout(Xd_0__inst_mult_14_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_48 (
// Equation(s):
// Xd_0__inst_mult_15_49  = SUM(( !Xd_0__inst_mult_15_4_q  $ (((!Xd_0__inst_mult_15_2_q ) # (!Xd_0__inst_mult_15_3_q ))) ) + ( Xd_0__inst_mult_15_98  ) + ( Xd_0__inst_mult_15_97  ))
// Xd_0__inst_mult_15_50  = CARRY(( !Xd_0__inst_mult_15_4_q  $ (((!Xd_0__inst_mult_15_2_q ) # (!Xd_0__inst_mult_15_3_q ))) ) + ( Xd_0__inst_mult_15_98  ) + ( Xd_0__inst_mult_15_97  ))
// Xd_0__inst_mult_15_51  = SHARE((Xd_0__inst_mult_15_2_q  & (Xd_0__inst_mult_15_3_q  & Xd_0__inst_mult_15_4_q )))

	.dataa(!Xd_0__inst_mult_15_2_q ),
	.datab(!Xd_0__inst_mult_15_3_q ),
	.datac(!Xd_0__inst_mult_15_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_97 ),
	.sharein(Xd_0__inst_mult_15_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_49 ),
	.cout(Xd_0__inst_mult_15_50 ),
	.shareout(Xd_0__inst_mult_15_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_48 (
// Equation(s):
// Xd_0__inst_mult_12_49  = SUM(( !Xd_0__inst_mult_12_4_q  $ (((!Xd_0__inst_mult_12_2_q ) # (!Xd_0__inst_mult_12_3_q ))) ) + ( Xd_0__inst_mult_12_98  ) + ( Xd_0__inst_mult_12_97  ))
// Xd_0__inst_mult_12_50  = CARRY(( !Xd_0__inst_mult_12_4_q  $ (((!Xd_0__inst_mult_12_2_q ) # (!Xd_0__inst_mult_12_3_q ))) ) + ( Xd_0__inst_mult_12_98  ) + ( Xd_0__inst_mult_12_97  ))
// Xd_0__inst_mult_12_51  = SHARE((Xd_0__inst_mult_12_2_q  & (Xd_0__inst_mult_12_3_q  & Xd_0__inst_mult_12_4_q )))

	.dataa(!Xd_0__inst_mult_12_2_q ),
	.datab(!Xd_0__inst_mult_12_3_q ),
	.datac(!Xd_0__inst_mult_12_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_97 ),
	.sharein(Xd_0__inst_mult_12_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_49 ),
	.cout(Xd_0__inst_mult_12_50 ),
	.shareout(Xd_0__inst_mult_12_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_48 (
// Equation(s):
// Xd_0__inst_mult_13_49  = SUM(( !Xd_0__inst_mult_13_4_q  $ (((!Xd_0__inst_mult_13_2_q ) # (!Xd_0__inst_mult_13_3_q ))) ) + ( Xd_0__inst_mult_13_98  ) + ( Xd_0__inst_mult_13_97  ))
// Xd_0__inst_mult_13_50  = CARRY(( !Xd_0__inst_mult_13_4_q  $ (((!Xd_0__inst_mult_13_2_q ) # (!Xd_0__inst_mult_13_3_q ))) ) + ( Xd_0__inst_mult_13_98  ) + ( Xd_0__inst_mult_13_97  ))
// Xd_0__inst_mult_13_51  = SHARE((Xd_0__inst_mult_13_2_q  & (Xd_0__inst_mult_13_3_q  & Xd_0__inst_mult_13_4_q )))

	.dataa(!Xd_0__inst_mult_13_2_q ),
	.datab(!Xd_0__inst_mult_13_3_q ),
	.datac(!Xd_0__inst_mult_13_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_97 ),
	.sharein(Xd_0__inst_mult_13_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_49 ),
	.cout(Xd_0__inst_mult_13_50 ),
	.shareout(Xd_0__inst_mult_13_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_48 (
// Equation(s):
// Xd_0__inst_mult_10_49  = SUM(( !Xd_0__inst_mult_10_4_q  $ (((!Xd_0__inst_mult_10_2_q ) # (!Xd_0__inst_mult_10_3_q ))) ) + ( Xd_0__inst_mult_10_98  ) + ( Xd_0__inst_mult_10_97  ))
// Xd_0__inst_mult_10_50  = CARRY(( !Xd_0__inst_mult_10_4_q  $ (((!Xd_0__inst_mult_10_2_q ) # (!Xd_0__inst_mult_10_3_q ))) ) + ( Xd_0__inst_mult_10_98  ) + ( Xd_0__inst_mult_10_97  ))
// Xd_0__inst_mult_10_51  = SHARE((Xd_0__inst_mult_10_2_q  & (Xd_0__inst_mult_10_3_q  & Xd_0__inst_mult_10_4_q )))

	.dataa(!Xd_0__inst_mult_10_2_q ),
	.datab(!Xd_0__inst_mult_10_3_q ),
	.datac(!Xd_0__inst_mult_10_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_97 ),
	.sharein(Xd_0__inst_mult_10_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_49 ),
	.cout(Xd_0__inst_mult_10_50 ),
	.shareout(Xd_0__inst_mult_10_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_48 (
// Equation(s):
// Xd_0__inst_mult_11_49  = SUM(( !Xd_0__inst_mult_11_4_q  $ (((!Xd_0__inst_mult_11_2_q ) # (!Xd_0__inst_mult_11_3_q ))) ) + ( Xd_0__inst_mult_11_98  ) + ( Xd_0__inst_mult_11_97  ))
// Xd_0__inst_mult_11_50  = CARRY(( !Xd_0__inst_mult_11_4_q  $ (((!Xd_0__inst_mult_11_2_q ) # (!Xd_0__inst_mult_11_3_q ))) ) + ( Xd_0__inst_mult_11_98  ) + ( Xd_0__inst_mult_11_97  ))
// Xd_0__inst_mult_11_51  = SHARE((Xd_0__inst_mult_11_2_q  & (Xd_0__inst_mult_11_3_q  & Xd_0__inst_mult_11_4_q )))

	.dataa(!Xd_0__inst_mult_11_2_q ),
	.datab(!Xd_0__inst_mult_11_3_q ),
	.datac(!Xd_0__inst_mult_11_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_97 ),
	.sharein(Xd_0__inst_mult_11_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_49 ),
	.cout(Xd_0__inst_mult_11_50 ),
	.shareout(Xd_0__inst_mult_11_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_48 (
// Equation(s):
// Xd_0__inst_mult_8_49  = SUM(( !Xd_0__inst_mult_8_4_q  $ (((!Xd_0__inst_mult_8_2_q ) # (!Xd_0__inst_mult_8_3_q ))) ) + ( Xd_0__inst_mult_8_98  ) + ( Xd_0__inst_mult_8_97  ))
// Xd_0__inst_mult_8_50  = CARRY(( !Xd_0__inst_mult_8_4_q  $ (((!Xd_0__inst_mult_8_2_q ) # (!Xd_0__inst_mult_8_3_q ))) ) + ( Xd_0__inst_mult_8_98  ) + ( Xd_0__inst_mult_8_97  ))
// Xd_0__inst_mult_8_51  = SHARE((Xd_0__inst_mult_8_2_q  & (Xd_0__inst_mult_8_3_q  & Xd_0__inst_mult_8_4_q )))

	.dataa(!Xd_0__inst_mult_8_2_q ),
	.datab(!Xd_0__inst_mult_8_3_q ),
	.datac(!Xd_0__inst_mult_8_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_97 ),
	.sharein(Xd_0__inst_mult_8_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_49 ),
	.cout(Xd_0__inst_mult_8_50 ),
	.shareout(Xd_0__inst_mult_8_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_48 (
// Equation(s):
// Xd_0__inst_mult_9_49  = SUM(( !Xd_0__inst_mult_9_4_q  $ (((!Xd_0__inst_mult_9_2_q ) # (!Xd_0__inst_mult_9_3_q ))) ) + ( Xd_0__inst_mult_9_98  ) + ( Xd_0__inst_mult_9_97  ))
// Xd_0__inst_mult_9_50  = CARRY(( !Xd_0__inst_mult_9_4_q  $ (((!Xd_0__inst_mult_9_2_q ) # (!Xd_0__inst_mult_9_3_q ))) ) + ( Xd_0__inst_mult_9_98  ) + ( Xd_0__inst_mult_9_97  ))
// Xd_0__inst_mult_9_51  = SHARE((Xd_0__inst_mult_9_2_q  & (Xd_0__inst_mult_9_3_q  & Xd_0__inst_mult_9_4_q )))

	.dataa(!Xd_0__inst_mult_9_2_q ),
	.datab(!Xd_0__inst_mult_9_3_q ),
	.datac(!Xd_0__inst_mult_9_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_97 ),
	.sharein(Xd_0__inst_mult_9_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_49 ),
	.cout(Xd_0__inst_mult_9_50 ),
	.shareout(Xd_0__inst_mult_9_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_48 (
// Equation(s):
// Xd_0__inst_mult_6_49  = SUM(( !Xd_0__inst_mult_6_4_q  $ (((!Xd_0__inst_mult_6_2_q ) # (!Xd_0__inst_mult_6_3_q ))) ) + ( Xd_0__inst_mult_6_98  ) + ( Xd_0__inst_mult_6_97  ))
// Xd_0__inst_mult_6_50  = CARRY(( !Xd_0__inst_mult_6_4_q  $ (((!Xd_0__inst_mult_6_2_q ) # (!Xd_0__inst_mult_6_3_q ))) ) + ( Xd_0__inst_mult_6_98  ) + ( Xd_0__inst_mult_6_97  ))
// Xd_0__inst_mult_6_51  = SHARE((Xd_0__inst_mult_6_2_q  & (Xd_0__inst_mult_6_3_q  & Xd_0__inst_mult_6_4_q )))

	.dataa(!Xd_0__inst_mult_6_2_q ),
	.datab(!Xd_0__inst_mult_6_3_q ),
	.datac(!Xd_0__inst_mult_6_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_97 ),
	.sharein(Xd_0__inst_mult_6_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_49 ),
	.cout(Xd_0__inst_mult_6_50 ),
	.shareout(Xd_0__inst_mult_6_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_48 (
// Equation(s):
// Xd_0__inst_mult_7_49  = SUM(( !Xd_0__inst_mult_7_4_q  $ (((!Xd_0__inst_mult_7_2_q ) # (!Xd_0__inst_mult_7_3_q ))) ) + ( Xd_0__inst_mult_7_98  ) + ( Xd_0__inst_mult_7_97  ))
// Xd_0__inst_mult_7_50  = CARRY(( !Xd_0__inst_mult_7_4_q  $ (((!Xd_0__inst_mult_7_2_q ) # (!Xd_0__inst_mult_7_3_q ))) ) + ( Xd_0__inst_mult_7_98  ) + ( Xd_0__inst_mult_7_97  ))
// Xd_0__inst_mult_7_51  = SHARE((Xd_0__inst_mult_7_2_q  & (Xd_0__inst_mult_7_3_q  & Xd_0__inst_mult_7_4_q )))

	.dataa(!Xd_0__inst_mult_7_2_q ),
	.datab(!Xd_0__inst_mult_7_3_q ),
	.datac(!Xd_0__inst_mult_7_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_97 ),
	.sharein(Xd_0__inst_mult_7_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_49 ),
	.cout(Xd_0__inst_mult_7_50 ),
	.shareout(Xd_0__inst_mult_7_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_48 (
// Equation(s):
// Xd_0__inst_mult_4_49  = SUM(( !Xd_0__inst_mult_4_4_q  $ (((!Xd_0__inst_mult_4_2_q ) # (!Xd_0__inst_mult_4_3_q ))) ) + ( Xd_0__inst_mult_4_98  ) + ( Xd_0__inst_mult_4_97  ))
// Xd_0__inst_mult_4_50  = CARRY(( !Xd_0__inst_mult_4_4_q  $ (((!Xd_0__inst_mult_4_2_q ) # (!Xd_0__inst_mult_4_3_q ))) ) + ( Xd_0__inst_mult_4_98  ) + ( Xd_0__inst_mult_4_97  ))
// Xd_0__inst_mult_4_51  = SHARE((Xd_0__inst_mult_4_2_q  & (Xd_0__inst_mult_4_3_q  & Xd_0__inst_mult_4_4_q )))

	.dataa(!Xd_0__inst_mult_4_2_q ),
	.datab(!Xd_0__inst_mult_4_3_q ),
	.datac(!Xd_0__inst_mult_4_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_97 ),
	.sharein(Xd_0__inst_mult_4_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_49 ),
	.cout(Xd_0__inst_mult_4_50 ),
	.shareout(Xd_0__inst_mult_4_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_48 (
// Equation(s):
// Xd_0__inst_mult_5_49  = SUM(( !Xd_0__inst_mult_5_4_q  $ (((!Xd_0__inst_mult_5_2_q ) # (!Xd_0__inst_mult_5_3_q ))) ) + ( Xd_0__inst_mult_5_98  ) + ( Xd_0__inst_mult_5_97  ))
// Xd_0__inst_mult_5_50  = CARRY(( !Xd_0__inst_mult_5_4_q  $ (((!Xd_0__inst_mult_5_2_q ) # (!Xd_0__inst_mult_5_3_q ))) ) + ( Xd_0__inst_mult_5_98  ) + ( Xd_0__inst_mult_5_97  ))
// Xd_0__inst_mult_5_51  = SHARE((Xd_0__inst_mult_5_2_q  & (Xd_0__inst_mult_5_3_q  & Xd_0__inst_mult_5_4_q )))

	.dataa(!Xd_0__inst_mult_5_2_q ),
	.datab(!Xd_0__inst_mult_5_3_q ),
	.datac(!Xd_0__inst_mult_5_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_97 ),
	.sharein(Xd_0__inst_mult_5_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_49 ),
	.cout(Xd_0__inst_mult_5_50 ),
	.shareout(Xd_0__inst_mult_5_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_48 (
// Equation(s):
// Xd_0__inst_mult_2_49  = SUM(( !Xd_0__inst_mult_2_4_q  $ (((!Xd_0__inst_mult_2_2_q ) # (!Xd_0__inst_mult_2_3_q ))) ) + ( Xd_0__inst_mult_2_98  ) + ( Xd_0__inst_mult_2_97  ))
// Xd_0__inst_mult_2_50  = CARRY(( !Xd_0__inst_mult_2_4_q  $ (((!Xd_0__inst_mult_2_2_q ) # (!Xd_0__inst_mult_2_3_q ))) ) + ( Xd_0__inst_mult_2_98  ) + ( Xd_0__inst_mult_2_97  ))
// Xd_0__inst_mult_2_51  = SHARE((Xd_0__inst_mult_2_2_q  & (Xd_0__inst_mult_2_3_q  & Xd_0__inst_mult_2_4_q )))

	.dataa(!Xd_0__inst_mult_2_2_q ),
	.datab(!Xd_0__inst_mult_2_3_q ),
	.datac(!Xd_0__inst_mult_2_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_97 ),
	.sharein(Xd_0__inst_mult_2_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_49 ),
	.cout(Xd_0__inst_mult_2_50 ),
	.shareout(Xd_0__inst_mult_2_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_48 (
// Equation(s):
// Xd_0__inst_mult_3_49  = SUM(( !Xd_0__inst_mult_3_4_q  $ (((!Xd_0__inst_mult_3_2_q ) # (!Xd_0__inst_mult_3_3_q ))) ) + ( Xd_0__inst_mult_3_98  ) + ( Xd_0__inst_mult_3_97  ))
// Xd_0__inst_mult_3_50  = CARRY(( !Xd_0__inst_mult_3_4_q  $ (((!Xd_0__inst_mult_3_2_q ) # (!Xd_0__inst_mult_3_3_q ))) ) + ( Xd_0__inst_mult_3_98  ) + ( Xd_0__inst_mult_3_97  ))
// Xd_0__inst_mult_3_51  = SHARE((Xd_0__inst_mult_3_2_q  & (Xd_0__inst_mult_3_3_q  & Xd_0__inst_mult_3_4_q )))

	.dataa(!Xd_0__inst_mult_3_2_q ),
	.datab(!Xd_0__inst_mult_3_3_q ),
	.datac(!Xd_0__inst_mult_3_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_97 ),
	.sharein(Xd_0__inst_mult_3_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_49 ),
	.cout(Xd_0__inst_mult_3_50 ),
	.shareout(Xd_0__inst_mult_3_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_48 (
// Equation(s):
// Xd_0__inst_mult_0_49  = SUM(( !Xd_0__inst_mult_0_4_q  $ (((!Xd_0__inst_mult_0_2_q ) # (!Xd_0__inst_mult_0_3_q ))) ) + ( Xd_0__inst_mult_0_98  ) + ( Xd_0__inst_mult_0_97  ))
// Xd_0__inst_mult_0_50  = CARRY(( !Xd_0__inst_mult_0_4_q  $ (((!Xd_0__inst_mult_0_2_q ) # (!Xd_0__inst_mult_0_3_q ))) ) + ( Xd_0__inst_mult_0_98  ) + ( Xd_0__inst_mult_0_97  ))
// Xd_0__inst_mult_0_51  = SHARE((Xd_0__inst_mult_0_2_q  & (Xd_0__inst_mult_0_3_q  & Xd_0__inst_mult_0_4_q )))

	.dataa(!Xd_0__inst_mult_0_2_q ),
	.datab(!Xd_0__inst_mult_0_3_q ),
	.datac(!Xd_0__inst_mult_0_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_97 ),
	.sharein(Xd_0__inst_mult_0_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_49 ),
	.cout(Xd_0__inst_mult_0_50 ),
	.shareout(Xd_0__inst_mult_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_48 (
// Equation(s):
// Xd_0__inst_mult_1_49  = SUM(( !Xd_0__inst_mult_1_4_q  $ (((!Xd_0__inst_mult_1_2_q ) # (!Xd_0__inst_mult_1_3_q ))) ) + ( Xd_0__inst_mult_1_98  ) + ( Xd_0__inst_mult_1_97  ))
// Xd_0__inst_mult_1_50  = CARRY(( !Xd_0__inst_mult_1_4_q  $ (((!Xd_0__inst_mult_1_2_q ) # (!Xd_0__inst_mult_1_3_q ))) ) + ( Xd_0__inst_mult_1_98  ) + ( Xd_0__inst_mult_1_97  ))
// Xd_0__inst_mult_1_51  = SHARE((Xd_0__inst_mult_1_2_q  & (Xd_0__inst_mult_1_3_q  & Xd_0__inst_mult_1_4_q )))

	.dataa(!Xd_0__inst_mult_1_2_q ),
	.datab(!Xd_0__inst_mult_1_3_q ),
	.datac(!Xd_0__inst_mult_1_4_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_97 ),
	.sharein(Xd_0__inst_mult_1_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_49 ),
	.cout(Xd_0__inst_mult_1_50 ),
	.shareout(Xd_0__inst_mult_1_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_28 (
// Equation(s):
// Xd_0__inst_mult_28_53  = SUM(( !Xd_0__inst_mult_28_5_q  $ (!Xd_0__inst_mult_28_6_q  $ (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_3_q )))) ) + ( Xd_0__inst_mult_28_51  ) + ( Xd_0__inst_mult_28_50  ))
// Xd_0__inst_mult_28_54  = CARRY(( !Xd_0__inst_mult_28_5_q  $ (!Xd_0__inst_mult_28_6_q  $ (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_3_q )))) ) + ( Xd_0__inst_mult_28_51  ) + ( Xd_0__inst_mult_28_50  ))
// Xd_0__inst_mult_28_55  = SHARE((!Xd_0__inst_mult_28_5_q  & (Xd_0__inst_mult_28_6_q  & (Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_3_q ))) # (Xd_0__inst_mult_28_5_q  & (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_3_q )) # (Xd_0__inst_mult_28_6_q ))))

	.dataa(!Xd_0__inst_mult_28_5_q ),
	.datab(!Xd_0__inst_mult_28_6_q ),
	.datac(!Xd_0__inst_mult_28_7_q ),
	.datad(!Xd_0__inst_mult_28_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_50 ),
	.sharein(Xd_0__inst_mult_28_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_53 ),
	.cout(Xd_0__inst_mult_28_54 ),
	.shareout(Xd_0__inst_mult_28_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_29 (
// Equation(s):
// Xd_0__inst_mult_29_53  = SUM(( !Xd_0__inst_mult_29_5_q  $ (!Xd_0__inst_mult_29_6_q  $ (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_3_q )))) ) + ( Xd_0__inst_mult_29_51  ) + ( Xd_0__inst_mult_29_50  ))
// Xd_0__inst_mult_29_54  = CARRY(( !Xd_0__inst_mult_29_5_q  $ (!Xd_0__inst_mult_29_6_q  $ (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_3_q )))) ) + ( Xd_0__inst_mult_29_51  ) + ( Xd_0__inst_mult_29_50  ))
// Xd_0__inst_mult_29_55  = SHARE((!Xd_0__inst_mult_29_5_q  & (Xd_0__inst_mult_29_6_q  & (Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_3_q ))) # (Xd_0__inst_mult_29_5_q  & (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_3_q )) # (Xd_0__inst_mult_29_6_q ))))

	.dataa(!Xd_0__inst_mult_29_5_q ),
	.datab(!Xd_0__inst_mult_29_6_q ),
	.datac(!Xd_0__inst_mult_29_7_q ),
	.datad(!Xd_0__inst_mult_29_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_50 ),
	.sharein(Xd_0__inst_mult_29_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_53 ),
	.cout(Xd_0__inst_mult_29_54 ),
	.shareout(Xd_0__inst_mult_29_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_26 (
// Equation(s):
// Xd_0__inst_mult_26_53  = SUM(( !Xd_0__inst_mult_26_5_q  $ (!Xd_0__inst_mult_26_6_q  $ (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_3_q )))) ) + ( Xd_0__inst_mult_26_51  ) + ( Xd_0__inst_mult_26_50  ))
// Xd_0__inst_mult_26_54  = CARRY(( !Xd_0__inst_mult_26_5_q  $ (!Xd_0__inst_mult_26_6_q  $ (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_3_q )))) ) + ( Xd_0__inst_mult_26_51  ) + ( Xd_0__inst_mult_26_50  ))
// Xd_0__inst_mult_26_55  = SHARE((!Xd_0__inst_mult_26_5_q  & (Xd_0__inst_mult_26_6_q  & (Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_3_q ))) # (Xd_0__inst_mult_26_5_q  & (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_3_q )) # (Xd_0__inst_mult_26_6_q ))))

	.dataa(!Xd_0__inst_mult_26_5_q ),
	.datab(!Xd_0__inst_mult_26_6_q ),
	.datac(!Xd_0__inst_mult_26_7_q ),
	.datad(!Xd_0__inst_mult_26_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_50 ),
	.sharein(Xd_0__inst_mult_26_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_53 ),
	.cout(Xd_0__inst_mult_26_54 ),
	.shareout(Xd_0__inst_mult_26_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_27 (
// Equation(s):
// Xd_0__inst_mult_27_53  = SUM(( !Xd_0__inst_mult_27_5_q  $ (!Xd_0__inst_mult_27_6_q  $ (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_3_q )))) ) + ( Xd_0__inst_mult_27_51  ) + ( Xd_0__inst_mult_27_50  ))
// Xd_0__inst_mult_27_54  = CARRY(( !Xd_0__inst_mult_27_5_q  $ (!Xd_0__inst_mult_27_6_q  $ (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_3_q )))) ) + ( Xd_0__inst_mult_27_51  ) + ( Xd_0__inst_mult_27_50  ))
// Xd_0__inst_mult_27_55  = SHARE((!Xd_0__inst_mult_27_5_q  & (Xd_0__inst_mult_27_6_q  & (Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_3_q ))) # (Xd_0__inst_mult_27_5_q  & (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_3_q )) # (Xd_0__inst_mult_27_6_q ))))

	.dataa(!Xd_0__inst_mult_27_5_q ),
	.datab(!Xd_0__inst_mult_27_6_q ),
	.datac(!Xd_0__inst_mult_27_7_q ),
	.datad(!Xd_0__inst_mult_27_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_50 ),
	.sharein(Xd_0__inst_mult_27_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_53 ),
	.cout(Xd_0__inst_mult_27_54 ),
	.shareout(Xd_0__inst_mult_27_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_24 (
// Equation(s):
// Xd_0__inst_mult_24_53  = SUM(( !Xd_0__inst_mult_24_5_q  $ (!Xd_0__inst_mult_24_6_q  $ (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_3_q )))) ) + ( Xd_0__inst_mult_24_51  ) + ( Xd_0__inst_mult_24_50  ))
// Xd_0__inst_mult_24_54  = CARRY(( !Xd_0__inst_mult_24_5_q  $ (!Xd_0__inst_mult_24_6_q  $ (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_3_q )))) ) + ( Xd_0__inst_mult_24_51  ) + ( Xd_0__inst_mult_24_50  ))
// Xd_0__inst_mult_24_55  = SHARE((!Xd_0__inst_mult_24_5_q  & (Xd_0__inst_mult_24_6_q  & (Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_3_q ))) # (Xd_0__inst_mult_24_5_q  & (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_3_q )) # (Xd_0__inst_mult_24_6_q ))))

	.dataa(!Xd_0__inst_mult_24_5_q ),
	.datab(!Xd_0__inst_mult_24_6_q ),
	.datac(!Xd_0__inst_mult_24_7_q ),
	.datad(!Xd_0__inst_mult_24_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_50 ),
	.sharein(Xd_0__inst_mult_24_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_53 ),
	.cout(Xd_0__inst_mult_24_54 ),
	.shareout(Xd_0__inst_mult_24_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_25 (
// Equation(s):
// Xd_0__inst_mult_25_53  = SUM(( !Xd_0__inst_mult_25_5_q  $ (!Xd_0__inst_mult_25_6_q  $ (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_3_q )))) ) + ( Xd_0__inst_mult_25_51  ) + ( Xd_0__inst_mult_25_50  ))
// Xd_0__inst_mult_25_54  = CARRY(( !Xd_0__inst_mult_25_5_q  $ (!Xd_0__inst_mult_25_6_q  $ (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_3_q )))) ) + ( Xd_0__inst_mult_25_51  ) + ( Xd_0__inst_mult_25_50  ))
// Xd_0__inst_mult_25_55  = SHARE((!Xd_0__inst_mult_25_5_q  & (Xd_0__inst_mult_25_6_q  & (Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_3_q ))) # (Xd_0__inst_mult_25_5_q  & (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_3_q )) # (Xd_0__inst_mult_25_6_q ))))

	.dataa(!Xd_0__inst_mult_25_5_q ),
	.datab(!Xd_0__inst_mult_25_6_q ),
	.datac(!Xd_0__inst_mult_25_7_q ),
	.datad(!Xd_0__inst_mult_25_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_50 ),
	.sharein(Xd_0__inst_mult_25_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_53 ),
	.cout(Xd_0__inst_mult_25_54 ),
	.shareout(Xd_0__inst_mult_25_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_22 (
// Equation(s):
// Xd_0__inst_mult_22_53  = SUM(( !Xd_0__inst_mult_22_5_q  $ (!Xd_0__inst_mult_22_6_q  $ (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_3_q )))) ) + ( Xd_0__inst_mult_22_51  ) + ( Xd_0__inst_mult_22_50  ))
// Xd_0__inst_mult_22_54  = CARRY(( !Xd_0__inst_mult_22_5_q  $ (!Xd_0__inst_mult_22_6_q  $ (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_3_q )))) ) + ( Xd_0__inst_mult_22_51  ) + ( Xd_0__inst_mult_22_50  ))
// Xd_0__inst_mult_22_55  = SHARE((!Xd_0__inst_mult_22_5_q  & (Xd_0__inst_mult_22_6_q  & (Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_3_q ))) # (Xd_0__inst_mult_22_5_q  & (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_3_q )) # (Xd_0__inst_mult_22_6_q ))))

	.dataa(!Xd_0__inst_mult_22_5_q ),
	.datab(!Xd_0__inst_mult_22_6_q ),
	.datac(!Xd_0__inst_mult_22_7_q ),
	.datad(!Xd_0__inst_mult_22_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_50 ),
	.sharein(Xd_0__inst_mult_22_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_53 ),
	.cout(Xd_0__inst_mult_22_54 ),
	.shareout(Xd_0__inst_mult_22_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_23 (
// Equation(s):
// Xd_0__inst_mult_23_53  = SUM(( !Xd_0__inst_mult_23_5_q  $ (!Xd_0__inst_mult_23_6_q  $ (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_3_q )))) ) + ( Xd_0__inst_mult_23_51  ) + ( Xd_0__inst_mult_23_50  ))
// Xd_0__inst_mult_23_54  = CARRY(( !Xd_0__inst_mult_23_5_q  $ (!Xd_0__inst_mult_23_6_q  $ (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_3_q )))) ) + ( Xd_0__inst_mult_23_51  ) + ( Xd_0__inst_mult_23_50  ))
// Xd_0__inst_mult_23_55  = SHARE((!Xd_0__inst_mult_23_5_q  & (Xd_0__inst_mult_23_6_q  & (Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_3_q ))) # (Xd_0__inst_mult_23_5_q  & (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_3_q )) # (Xd_0__inst_mult_23_6_q ))))

	.dataa(!Xd_0__inst_mult_23_5_q ),
	.datab(!Xd_0__inst_mult_23_6_q ),
	.datac(!Xd_0__inst_mult_23_7_q ),
	.datad(!Xd_0__inst_mult_23_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_50 ),
	.sharein(Xd_0__inst_mult_23_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_53 ),
	.cout(Xd_0__inst_mult_23_54 ),
	.shareout(Xd_0__inst_mult_23_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_20 (
// Equation(s):
// Xd_0__inst_mult_20_53  = SUM(( !Xd_0__inst_mult_20_5_q  $ (!Xd_0__inst_mult_20_6_q  $ (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_3_q )))) ) + ( Xd_0__inst_mult_20_51  ) + ( Xd_0__inst_mult_20_50  ))
// Xd_0__inst_mult_20_54  = CARRY(( !Xd_0__inst_mult_20_5_q  $ (!Xd_0__inst_mult_20_6_q  $ (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_3_q )))) ) + ( Xd_0__inst_mult_20_51  ) + ( Xd_0__inst_mult_20_50  ))
// Xd_0__inst_mult_20_55  = SHARE((!Xd_0__inst_mult_20_5_q  & (Xd_0__inst_mult_20_6_q  & (Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_3_q ))) # (Xd_0__inst_mult_20_5_q  & (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_3_q )) # (Xd_0__inst_mult_20_6_q ))))

	.dataa(!Xd_0__inst_mult_20_5_q ),
	.datab(!Xd_0__inst_mult_20_6_q ),
	.datac(!Xd_0__inst_mult_20_7_q ),
	.datad(!Xd_0__inst_mult_20_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_50 ),
	.sharein(Xd_0__inst_mult_20_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_53 ),
	.cout(Xd_0__inst_mult_20_54 ),
	.shareout(Xd_0__inst_mult_20_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_21 (
// Equation(s):
// Xd_0__inst_mult_21_53  = SUM(( !Xd_0__inst_mult_21_5_q  $ (!Xd_0__inst_mult_21_6_q  $ (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_3_q )))) ) + ( Xd_0__inst_mult_21_51  ) + ( Xd_0__inst_mult_21_50  ))
// Xd_0__inst_mult_21_54  = CARRY(( !Xd_0__inst_mult_21_5_q  $ (!Xd_0__inst_mult_21_6_q  $ (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_3_q )))) ) + ( Xd_0__inst_mult_21_51  ) + ( Xd_0__inst_mult_21_50  ))
// Xd_0__inst_mult_21_55  = SHARE((!Xd_0__inst_mult_21_5_q  & (Xd_0__inst_mult_21_6_q  & (Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_3_q ))) # (Xd_0__inst_mult_21_5_q  & (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_3_q )) # (Xd_0__inst_mult_21_6_q ))))

	.dataa(!Xd_0__inst_mult_21_5_q ),
	.datab(!Xd_0__inst_mult_21_6_q ),
	.datac(!Xd_0__inst_mult_21_7_q ),
	.datad(!Xd_0__inst_mult_21_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_50 ),
	.sharein(Xd_0__inst_mult_21_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_53 ),
	.cout(Xd_0__inst_mult_21_54 ),
	.shareout(Xd_0__inst_mult_21_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_18 (
// Equation(s):
// Xd_0__inst_mult_18_53  = SUM(( !Xd_0__inst_mult_18_5_q  $ (!Xd_0__inst_mult_18_6_q  $ (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_3_q )))) ) + ( Xd_0__inst_mult_18_51  ) + ( Xd_0__inst_mult_18_50  ))
// Xd_0__inst_mult_18_54  = CARRY(( !Xd_0__inst_mult_18_5_q  $ (!Xd_0__inst_mult_18_6_q  $ (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_3_q )))) ) + ( Xd_0__inst_mult_18_51  ) + ( Xd_0__inst_mult_18_50  ))
// Xd_0__inst_mult_18_55  = SHARE((!Xd_0__inst_mult_18_5_q  & (Xd_0__inst_mult_18_6_q  & (Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_3_q ))) # (Xd_0__inst_mult_18_5_q  & (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_3_q )) # (Xd_0__inst_mult_18_6_q ))))

	.dataa(!Xd_0__inst_mult_18_5_q ),
	.datab(!Xd_0__inst_mult_18_6_q ),
	.datac(!Xd_0__inst_mult_18_7_q ),
	.datad(!Xd_0__inst_mult_18_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_50 ),
	.sharein(Xd_0__inst_mult_18_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_53 ),
	.cout(Xd_0__inst_mult_18_54 ),
	.shareout(Xd_0__inst_mult_18_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_19 (
// Equation(s):
// Xd_0__inst_mult_19_53  = SUM(( !Xd_0__inst_mult_19_5_q  $ (!Xd_0__inst_mult_19_6_q  $ (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_3_q )))) ) + ( Xd_0__inst_mult_19_51  ) + ( Xd_0__inst_mult_19_50  ))
// Xd_0__inst_mult_19_54  = CARRY(( !Xd_0__inst_mult_19_5_q  $ (!Xd_0__inst_mult_19_6_q  $ (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_3_q )))) ) + ( Xd_0__inst_mult_19_51  ) + ( Xd_0__inst_mult_19_50  ))
// Xd_0__inst_mult_19_55  = SHARE((!Xd_0__inst_mult_19_5_q  & (Xd_0__inst_mult_19_6_q  & (Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_3_q ))) # (Xd_0__inst_mult_19_5_q  & (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_3_q )) # (Xd_0__inst_mult_19_6_q ))))

	.dataa(!Xd_0__inst_mult_19_5_q ),
	.datab(!Xd_0__inst_mult_19_6_q ),
	.datac(!Xd_0__inst_mult_19_7_q ),
	.datad(!Xd_0__inst_mult_19_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_50 ),
	.sharein(Xd_0__inst_mult_19_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_53 ),
	.cout(Xd_0__inst_mult_19_54 ),
	.shareout(Xd_0__inst_mult_19_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_16 (
// Equation(s):
// Xd_0__inst_mult_16_53  = SUM(( !Xd_0__inst_mult_16_5_q  $ (!Xd_0__inst_mult_16_6_q  $ (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_3_q )))) ) + ( Xd_0__inst_mult_16_51  ) + ( Xd_0__inst_mult_16_50  ))
// Xd_0__inst_mult_16_54  = CARRY(( !Xd_0__inst_mult_16_5_q  $ (!Xd_0__inst_mult_16_6_q  $ (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_3_q )))) ) + ( Xd_0__inst_mult_16_51  ) + ( Xd_0__inst_mult_16_50  ))
// Xd_0__inst_mult_16_55  = SHARE((!Xd_0__inst_mult_16_5_q  & (Xd_0__inst_mult_16_6_q  & (Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_3_q ))) # (Xd_0__inst_mult_16_5_q  & (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_3_q )) # (Xd_0__inst_mult_16_6_q ))))

	.dataa(!Xd_0__inst_mult_16_5_q ),
	.datab(!Xd_0__inst_mult_16_6_q ),
	.datac(!Xd_0__inst_mult_16_7_q ),
	.datad(!Xd_0__inst_mult_16_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_50 ),
	.sharein(Xd_0__inst_mult_16_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_53 ),
	.cout(Xd_0__inst_mult_16_54 ),
	.shareout(Xd_0__inst_mult_16_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_17 (
// Equation(s):
// Xd_0__inst_mult_17_53  = SUM(( !Xd_0__inst_mult_17_5_q  $ (!Xd_0__inst_mult_17_6_q  $ (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_3_q )))) ) + ( Xd_0__inst_mult_17_51  ) + ( Xd_0__inst_mult_17_50  ))
// Xd_0__inst_mult_17_54  = CARRY(( !Xd_0__inst_mult_17_5_q  $ (!Xd_0__inst_mult_17_6_q  $ (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_3_q )))) ) + ( Xd_0__inst_mult_17_51  ) + ( Xd_0__inst_mult_17_50  ))
// Xd_0__inst_mult_17_55  = SHARE((!Xd_0__inst_mult_17_5_q  & (Xd_0__inst_mult_17_6_q  & (Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_3_q ))) # (Xd_0__inst_mult_17_5_q  & (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_3_q )) # (Xd_0__inst_mult_17_6_q ))))

	.dataa(!Xd_0__inst_mult_17_5_q ),
	.datab(!Xd_0__inst_mult_17_6_q ),
	.datac(!Xd_0__inst_mult_17_7_q ),
	.datad(!Xd_0__inst_mult_17_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_50 ),
	.sharein(Xd_0__inst_mult_17_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_53 ),
	.cout(Xd_0__inst_mult_17_54 ),
	.shareout(Xd_0__inst_mult_17_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14 (
// Equation(s):
// Xd_0__inst_mult_14_53  = SUM(( !Xd_0__inst_mult_14_5_q  $ (!Xd_0__inst_mult_14_6_q  $ (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_3_q )))) ) + ( Xd_0__inst_mult_14_51  ) + ( Xd_0__inst_mult_14_50  ))
// Xd_0__inst_mult_14_54  = CARRY(( !Xd_0__inst_mult_14_5_q  $ (!Xd_0__inst_mult_14_6_q  $ (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_3_q )))) ) + ( Xd_0__inst_mult_14_51  ) + ( Xd_0__inst_mult_14_50  ))
// Xd_0__inst_mult_14_55  = SHARE((!Xd_0__inst_mult_14_5_q  & (Xd_0__inst_mult_14_6_q  & (Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_3_q ))) # (Xd_0__inst_mult_14_5_q  & (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_3_q )) # (Xd_0__inst_mult_14_6_q ))))

	.dataa(!Xd_0__inst_mult_14_5_q ),
	.datab(!Xd_0__inst_mult_14_6_q ),
	.datac(!Xd_0__inst_mult_14_7_q ),
	.datad(!Xd_0__inst_mult_14_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_50 ),
	.sharein(Xd_0__inst_mult_14_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_53 ),
	.cout(Xd_0__inst_mult_14_54 ),
	.shareout(Xd_0__inst_mult_14_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15 (
// Equation(s):
// Xd_0__inst_mult_15_53  = SUM(( !Xd_0__inst_mult_15_5_q  $ (!Xd_0__inst_mult_15_6_q  $ (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_3_q )))) ) + ( Xd_0__inst_mult_15_51  ) + ( Xd_0__inst_mult_15_50  ))
// Xd_0__inst_mult_15_54  = CARRY(( !Xd_0__inst_mult_15_5_q  $ (!Xd_0__inst_mult_15_6_q  $ (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_3_q )))) ) + ( Xd_0__inst_mult_15_51  ) + ( Xd_0__inst_mult_15_50  ))
// Xd_0__inst_mult_15_55  = SHARE((!Xd_0__inst_mult_15_5_q  & (Xd_0__inst_mult_15_6_q  & (Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_3_q ))) # (Xd_0__inst_mult_15_5_q  & (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_3_q )) # (Xd_0__inst_mult_15_6_q ))))

	.dataa(!Xd_0__inst_mult_15_5_q ),
	.datab(!Xd_0__inst_mult_15_6_q ),
	.datac(!Xd_0__inst_mult_15_7_q ),
	.datad(!Xd_0__inst_mult_15_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_50 ),
	.sharein(Xd_0__inst_mult_15_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_53 ),
	.cout(Xd_0__inst_mult_15_54 ),
	.shareout(Xd_0__inst_mult_15_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12 (
// Equation(s):
// Xd_0__inst_mult_12_53  = SUM(( !Xd_0__inst_mult_12_5_q  $ (!Xd_0__inst_mult_12_6_q  $ (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_3_q )))) ) + ( Xd_0__inst_mult_12_51  ) + ( Xd_0__inst_mult_12_50  ))
// Xd_0__inst_mult_12_54  = CARRY(( !Xd_0__inst_mult_12_5_q  $ (!Xd_0__inst_mult_12_6_q  $ (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_3_q )))) ) + ( Xd_0__inst_mult_12_51  ) + ( Xd_0__inst_mult_12_50  ))
// Xd_0__inst_mult_12_55  = SHARE((!Xd_0__inst_mult_12_5_q  & (Xd_0__inst_mult_12_6_q  & (Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_3_q ))) # (Xd_0__inst_mult_12_5_q  & (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_3_q )) # (Xd_0__inst_mult_12_6_q ))))

	.dataa(!Xd_0__inst_mult_12_5_q ),
	.datab(!Xd_0__inst_mult_12_6_q ),
	.datac(!Xd_0__inst_mult_12_7_q ),
	.datad(!Xd_0__inst_mult_12_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_50 ),
	.sharein(Xd_0__inst_mult_12_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_53 ),
	.cout(Xd_0__inst_mult_12_54 ),
	.shareout(Xd_0__inst_mult_12_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13 (
// Equation(s):
// Xd_0__inst_mult_13_53  = SUM(( !Xd_0__inst_mult_13_5_q  $ (!Xd_0__inst_mult_13_6_q  $ (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_3_q )))) ) + ( Xd_0__inst_mult_13_51  ) + ( Xd_0__inst_mult_13_50  ))
// Xd_0__inst_mult_13_54  = CARRY(( !Xd_0__inst_mult_13_5_q  $ (!Xd_0__inst_mult_13_6_q  $ (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_3_q )))) ) + ( Xd_0__inst_mult_13_51  ) + ( Xd_0__inst_mult_13_50  ))
// Xd_0__inst_mult_13_55  = SHARE((!Xd_0__inst_mult_13_5_q  & (Xd_0__inst_mult_13_6_q  & (Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_3_q ))) # (Xd_0__inst_mult_13_5_q  & (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_3_q )) # (Xd_0__inst_mult_13_6_q ))))

	.dataa(!Xd_0__inst_mult_13_5_q ),
	.datab(!Xd_0__inst_mult_13_6_q ),
	.datac(!Xd_0__inst_mult_13_7_q ),
	.datad(!Xd_0__inst_mult_13_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_50 ),
	.sharein(Xd_0__inst_mult_13_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_53 ),
	.cout(Xd_0__inst_mult_13_54 ),
	.shareout(Xd_0__inst_mult_13_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10 (
// Equation(s):
// Xd_0__inst_mult_10_53  = SUM(( !Xd_0__inst_mult_10_5_q  $ (!Xd_0__inst_mult_10_6_q  $ (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_3_q )))) ) + ( Xd_0__inst_mult_10_51  ) + ( Xd_0__inst_mult_10_50  ))
// Xd_0__inst_mult_10_54  = CARRY(( !Xd_0__inst_mult_10_5_q  $ (!Xd_0__inst_mult_10_6_q  $ (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_3_q )))) ) + ( Xd_0__inst_mult_10_51  ) + ( Xd_0__inst_mult_10_50  ))
// Xd_0__inst_mult_10_55  = SHARE((!Xd_0__inst_mult_10_5_q  & (Xd_0__inst_mult_10_6_q  & (Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_3_q ))) # (Xd_0__inst_mult_10_5_q  & (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_3_q )) # (Xd_0__inst_mult_10_6_q ))))

	.dataa(!Xd_0__inst_mult_10_5_q ),
	.datab(!Xd_0__inst_mult_10_6_q ),
	.datac(!Xd_0__inst_mult_10_7_q ),
	.datad(!Xd_0__inst_mult_10_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_50 ),
	.sharein(Xd_0__inst_mult_10_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_53 ),
	.cout(Xd_0__inst_mult_10_54 ),
	.shareout(Xd_0__inst_mult_10_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11 (
// Equation(s):
// Xd_0__inst_mult_11_53  = SUM(( !Xd_0__inst_mult_11_5_q  $ (!Xd_0__inst_mult_11_6_q  $ (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_3_q )))) ) + ( Xd_0__inst_mult_11_51  ) + ( Xd_0__inst_mult_11_50  ))
// Xd_0__inst_mult_11_54  = CARRY(( !Xd_0__inst_mult_11_5_q  $ (!Xd_0__inst_mult_11_6_q  $ (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_3_q )))) ) + ( Xd_0__inst_mult_11_51  ) + ( Xd_0__inst_mult_11_50  ))
// Xd_0__inst_mult_11_55  = SHARE((!Xd_0__inst_mult_11_5_q  & (Xd_0__inst_mult_11_6_q  & (Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_3_q ))) # (Xd_0__inst_mult_11_5_q  & (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_3_q )) # (Xd_0__inst_mult_11_6_q ))))

	.dataa(!Xd_0__inst_mult_11_5_q ),
	.datab(!Xd_0__inst_mult_11_6_q ),
	.datac(!Xd_0__inst_mult_11_7_q ),
	.datad(!Xd_0__inst_mult_11_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_50 ),
	.sharein(Xd_0__inst_mult_11_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_53 ),
	.cout(Xd_0__inst_mult_11_54 ),
	.shareout(Xd_0__inst_mult_11_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8 (
// Equation(s):
// Xd_0__inst_mult_8_53  = SUM(( !Xd_0__inst_mult_8_5_q  $ (!Xd_0__inst_mult_8_6_q  $ (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_3_q )))) ) + ( Xd_0__inst_mult_8_51  ) + ( Xd_0__inst_mult_8_50  ))
// Xd_0__inst_mult_8_54  = CARRY(( !Xd_0__inst_mult_8_5_q  $ (!Xd_0__inst_mult_8_6_q  $ (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_3_q )))) ) + ( Xd_0__inst_mult_8_51  ) + ( Xd_0__inst_mult_8_50  ))
// Xd_0__inst_mult_8_55  = SHARE((!Xd_0__inst_mult_8_5_q  & (Xd_0__inst_mult_8_6_q  & (Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_3_q ))) # (Xd_0__inst_mult_8_5_q  & (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_3_q )) # (Xd_0__inst_mult_8_6_q ))))

	.dataa(!Xd_0__inst_mult_8_5_q ),
	.datab(!Xd_0__inst_mult_8_6_q ),
	.datac(!Xd_0__inst_mult_8_7_q ),
	.datad(!Xd_0__inst_mult_8_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_50 ),
	.sharein(Xd_0__inst_mult_8_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_53 ),
	.cout(Xd_0__inst_mult_8_54 ),
	.shareout(Xd_0__inst_mult_8_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9 (
// Equation(s):
// Xd_0__inst_mult_9_53  = SUM(( !Xd_0__inst_mult_9_5_q  $ (!Xd_0__inst_mult_9_6_q  $ (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_3_q )))) ) + ( Xd_0__inst_mult_9_51  ) + ( Xd_0__inst_mult_9_50  ))
// Xd_0__inst_mult_9_54  = CARRY(( !Xd_0__inst_mult_9_5_q  $ (!Xd_0__inst_mult_9_6_q  $ (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_3_q )))) ) + ( Xd_0__inst_mult_9_51  ) + ( Xd_0__inst_mult_9_50  ))
// Xd_0__inst_mult_9_55  = SHARE((!Xd_0__inst_mult_9_5_q  & (Xd_0__inst_mult_9_6_q  & (Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_3_q ))) # (Xd_0__inst_mult_9_5_q  & (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_3_q )) # (Xd_0__inst_mult_9_6_q ))))

	.dataa(!Xd_0__inst_mult_9_5_q ),
	.datab(!Xd_0__inst_mult_9_6_q ),
	.datac(!Xd_0__inst_mult_9_7_q ),
	.datad(!Xd_0__inst_mult_9_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_50 ),
	.sharein(Xd_0__inst_mult_9_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_53 ),
	.cout(Xd_0__inst_mult_9_54 ),
	.shareout(Xd_0__inst_mult_9_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6 (
// Equation(s):
// Xd_0__inst_mult_6_53  = SUM(( !Xd_0__inst_mult_6_5_q  $ (!Xd_0__inst_mult_6_6_q  $ (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_3_q )))) ) + ( Xd_0__inst_mult_6_51  ) + ( Xd_0__inst_mult_6_50  ))
// Xd_0__inst_mult_6_54  = CARRY(( !Xd_0__inst_mult_6_5_q  $ (!Xd_0__inst_mult_6_6_q  $ (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_3_q )))) ) + ( Xd_0__inst_mult_6_51  ) + ( Xd_0__inst_mult_6_50  ))
// Xd_0__inst_mult_6_55  = SHARE((!Xd_0__inst_mult_6_5_q  & (Xd_0__inst_mult_6_6_q  & (Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_3_q ))) # (Xd_0__inst_mult_6_5_q  & (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_3_q )) # (Xd_0__inst_mult_6_6_q ))))

	.dataa(!Xd_0__inst_mult_6_5_q ),
	.datab(!Xd_0__inst_mult_6_6_q ),
	.datac(!Xd_0__inst_mult_6_7_q ),
	.datad(!Xd_0__inst_mult_6_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_50 ),
	.sharein(Xd_0__inst_mult_6_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_53 ),
	.cout(Xd_0__inst_mult_6_54 ),
	.shareout(Xd_0__inst_mult_6_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7 (
// Equation(s):
// Xd_0__inst_mult_7_53  = SUM(( !Xd_0__inst_mult_7_5_q  $ (!Xd_0__inst_mult_7_6_q  $ (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_3_q )))) ) + ( Xd_0__inst_mult_7_51  ) + ( Xd_0__inst_mult_7_50  ))
// Xd_0__inst_mult_7_54  = CARRY(( !Xd_0__inst_mult_7_5_q  $ (!Xd_0__inst_mult_7_6_q  $ (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_3_q )))) ) + ( Xd_0__inst_mult_7_51  ) + ( Xd_0__inst_mult_7_50  ))
// Xd_0__inst_mult_7_55  = SHARE((!Xd_0__inst_mult_7_5_q  & (Xd_0__inst_mult_7_6_q  & (Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_3_q ))) # (Xd_0__inst_mult_7_5_q  & (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_3_q )) # (Xd_0__inst_mult_7_6_q ))))

	.dataa(!Xd_0__inst_mult_7_5_q ),
	.datab(!Xd_0__inst_mult_7_6_q ),
	.datac(!Xd_0__inst_mult_7_7_q ),
	.datad(!Xd_0__inst_mult_7_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_50 ),
	.sharein(Xd_0__inst_mult_7_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_53 ),
	.cout(Xd_0__inst_mult_7_54 ),
	.shareout(Xd_0__inst_mult_7_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4 (
// Equation(s):
// Xd_0__inst_mult_4_53  = SUM(( !Xd_0__inst_mult_4_5_q  $ (!Xd_0__inst_mult_4_6_q  $ (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_3_q )))) ) + ( Xd_0__inst_mult_4_51  ) + ( Xd_0__inst_mult_4_50  ))
// Xd_0__inst_mult_4_54  = CARRY(( !Xd_0__inst_mult_4_5_q  $ (!Xd_0__inst_mult_4_6_q  $ (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_3_q )))) ) + ( Xd_0__inst_mult_4_51  ) + ( Xd_0__inst_mult_4_50  ))
// Xd_0__inst_mult_4_55  = SHARE((!Xd_0__inst_mult_4_5_q  & (Xd_0__inst_mult_4_6_q  & (Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_3_q ))) # (Xd_0__inst_mult_4_5_q  & (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_3_q )) # (Xd_0__inst_mult_4_6_q ))))

	.dataa(!Xd_0__inst_mult_4_5_q ),
	.datab(!Xd_0__inst_mult_4_6_q ),
	.datac(!Xd_0__inst_mult_4_7_q ),
	.datad(!Xd_0__inst_mult_4_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_50 ),
	.sharein(Xd_0__inst_mult_4_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_53 ),
	.cout(Xd_0__inst_mult_4_54 ),
	.shareout(Xd_0__inst_mult_4_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5 (
// Equation(s):
// Xd_0__inst_mult_5_53  = SUM(( !Xd_0__inst_mult_5_5_q  $ (!Xd_0__inst_mult_5_6_q  $ (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_3_q )))) ) + ( Xd_0__inst_mult_5_51  ) + ( Xd_0__inst_mult_5_50  ))
// Xd_0__inst_mult_5_54  = CARRY(( !Xd_0__inst_mult_5_5_q  $ (!Xd_0__inst_mult_5_6_q  $ (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_3_q )))) ) + ( Xd_0__inst_mult_5_51  ) + ( Xd_0__inst_mult_5_50  ))
// Xd_0__inst_mult_5_55  = SHARE((!Xd_0__inst_mult_5_5_q  & (Xd_0__inst_mult_5_6_q  & (Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_3_q ))) # (Xd_0__inst_mult_5_5_q  & (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_3_q )) # (Xd_0__inst_mult_5_6_q ))))

	.dataa(!Xd_0__inst_mult_5_5_q ),
	.datab(!Xd_0__inst_mult_5_6_q ),
	.datac(!Xd_0__inst_mult_5_7_q ),
	.datad(!Xd_0__inst_mult_5_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_50 ),
	.sharein(Xd_0__inst_mult_5_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_53 ),
	.cout(Xd_0__inst_mult_5_54 ),
	.shareout(Xd_0__inst_mult_5_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2 (
// Equation(s):
// Xd_0__inst_mult_2_53  = SUM(( !Xd_0__inst_mult_2_5_q  $ (!Xd_0__inst_mult_2_6_q  $ (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_3_q )))) ) + ( Xd_0__inst_mult_2_51  ) + ( Xd_0__inst_mult_2_50  ))
// Xd_0__inst_mult_2_54  = CARRY(( !Xd_0__inst_mult_2_5_q  $ (!Xd_0__inst_mult_2_6_q  $ (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_3_q )))) ) + ( Xd_0__inst_mult_2_51  ) + ( Xd_0__inst_mult_2_50  ))
// Xd_0__inst_mult_2_55  = SHARE((!Xd_0__inst_mult_2_5_q  & (Xd_0__inst_mult_2_6_q  & (Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_3_q ))) # (Xd_0__inst_mult_2_5_q  & (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_3_q )) # (Xd_0__inst_mult_2_6_q ))))

	.dataa(!Xd_0__inst_mult_2_5_q ),
	.datab(!Xd_0__inst_mult_2_6_q ),
	.datac(!Xd_0__inst_mult_2_7_q ),
	.datad(!Xd_0__inst_mult_2_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_50 ),
	.sharein(Xd_0__inst_mult_2_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_53 ),
	.cout(Xd_0__inst_mult_2_54 ),
	.shareout(Xd_0__inst_mult_2_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3 (
// Equation(s):
// Xd_0__inst_mult_3_53  = SUM(( !Xd_0__inst_mult_3_5_q  $ (!Xd_0__inst_mult_3_6_q  $ (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_3_q )))) ) + ( Xd_0__inst_mult_3_51  ) + ( Xd_0__inst_mult_3_50  ))
// Xd_0__inst_mult_3_54  = CARRY(( !Xd_0__inst_mult_3_5_q  $ (!Xd_0__inst_mult_3_6_q  $ (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_3_q )))) ) + ( Xd_0__inst_mult_3_51  ) + ( Xd_0__inst_mult_3_50  ))
// Xd_0__inst_mult_3_55  = SHARE((!Xd_0__inst_mult_3_5_q  & (Xd_0__inst_mult_3_6_q  & (Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_3_q ))) # (Xd_0__inst_mult_3_5_q  & (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_3_q )) # (Xd_0__inst_mult_3_6_q ))))

	.dataa(!Xd_0__inst_mult_3_5_q ),
	.datab(!Xd_0__inst_mult_3_6_q ),
	.datac(!Xd_0__inst_mult_3_7_q ),
	.datad(!Xd_0__inst_mult_3_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_50 ),
	.sharein(Xd_0__inst_mult_3_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_53 ),
	.cout(Xd_0__inst_mult_3_54 ),
	.shareout(Xd_0__inst_mult_3_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0 (
// Equation(s):
// Xd_0__inst_mult_0_53  = SUM(( !Xd_0__inst_mult_0_5_q  $ (!Xd_0__inst_mult_0_6_q  $ (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_3_q )))) ) + ( Xd_0__inst_mult_0_51  ) + ( Xd_0__inst_mult_0_50  ))
// Xd_0__inst_mult_0_54  = CARRY(( !Xd_0__inst_mult_0_5_q  $ (!Xd_0__inst_mult_0_6_q  $ (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_3_q )))) ) + ( Xd_0__inst_mult_0_51  ) + ( Xd_0__inst_mult_0_50  ))
// Xd_0__inst_mult_0_55  = SHARE((!Xd_0__inst_mult_0_5_q  & (Xd_0__inst_mult_0_6_q  & (Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_3_q ))) # (Xd_0__inst_mult_0_5_q  & (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_3_q )) # (Xd_0__inst_mult_0_6_q ))))

	.dataa(!Xd_0__inst_mult_0_5_q ),
	.datab(!Xd_0__inst_mult_0_6_q ),
	.datac(!Xd_0__inst_mult_0_7_q ),
	.datad(!Xd_0__inst_mult_0_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_50 ),
	.sharein(Xd_0__inst_mult_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_53 ),
	.cout(Xd_0__inst_mult_0_54 ),
	.shareout(Xd_0__inst_mult_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1 (
// Equation(s):
// Xd_0__inst_mult_1_53  = SUM(( !Xd_0__inst_mult_1_5_q  $ (!Xd_0__inst_mult_1_6_q  $ (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_3_q )))) ) + ( Xd_0__inst_mult_1_51  ) + ( Xd_0__inst_mult_1_50  ))
// Xd_0__inst_mult_1_54  = CARRY(( !Xd_0__inst_mult_1_5_q  $ (!Xd_0__inst_mult_1_6_q  $ (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_3_q )))) ) + ( Xd_0__inst_mult_1_51  ) + ( Xd_0__inst_mult_1_50  ))
// Xd_0__inst_mult_1_55  = SHARE((!Xd_0__inst_mult_1_5_q  & (Xd_0__inst_mult_1_6_q  & (Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_3_q ))) # (Xd_0__inst_mult_1_5_q  & (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_3_q )) # (Xd_0__inst_mult_1_6_q ))))

	.dataa(!Xd_0__inst_mult_1_5_q ),
	.datab(!Xd_0__inst_mult_1_6_q ),
	.datac(!Xd_0__inst_mult_1_7_q ),
	.datad(!Xd_0__inst_mult_1_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_50 ),
	.sharein(Xd_0__inst_mult_1_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_53 ),
	.cout(Xd_0__inst_mult_1_54 ),
	.shareout(Xd_0__inst_mult_1_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_28_21 (
// Equation(s):
// Xd_0__inst_mult_28_56  = SUM(( !Xd_0__inst_mult_28_8_q  $ (!Xd_0__inst_mult_28_9_q ) ) + ( Xd_0__inst_mult_28_55  ) + ( Xd_0__inst_mult_28_54  ))
// Xd_0__inst_mult_28_57  = CARRY(( !Xd_0__inst_mult_28_8_q  $ (!Xd_0__inst_mult_28_9_q ) ) + ( Xd_0__inst_mult_28_55  ) + ( Xd_0__inst_mult_28_54  ))
// Xd_0__inst_mult_28_58  = SHARE((Xd_0__inst_mult_28_8_q  & Xd_0__inst_mult_28_9_q ))

	.dataa(!Xd_0__inst_mult_28_8_q ),
	.datab(!Xd_0__inst_mult_28_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_54 ),
	.sharein(Xd_0__inst_mult_28_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_56 ),
	.cout(Xd_0__inst_mult_28_57 ),
	.shareout(Xd_0__inst_mult_28_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_29_21 (
// Equation(s):
// Xd_0__inst_mult_29_56  = SUM(( !Xd_0__inst_mult_29_8_q  $ (!Xd_0__inst_mult_29_9_q ) ) + ( Xd_0__inst_mult_29_55  ) + ( Xd_0__inst_mult_29_54  ))
// Xd_0__inst_mult_29_57  = CARRY(( !Xd_0__inst_mult_29_8_q  $ (!Xd_0__inst_mult_29_9_q ) ) + ( Xd_0__inst_mult_29_55  ) + ( Xd_0__inst_mult_29_54  ))
// Xd_0__inst_mult_29_58  = SHARE((Xd_0__inst_mult_29_8_q  & Xd_0__inst_mult_29_9_q ))

	.dataa(!Xd_0__inst_mult_29_8_q ),
	.datab(!Xd_0__inst_mult_29_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_54 ),
	.sharein(Xd_0__inst_mult_29_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_56 ),
	.cout(Xd_0__inst_mult_29_57 ),
	.shareout(Xd_0__inst_mult_29_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_26_21 (
// Equation(s):
// Xd_0__inst_mult_26_56  = SUM(( !Xd_0__inst_mult_26_8_q  $ (!Xd_0__inst_mult_26_9_q ) ) + ( Xd_0__inst_mult_26_55  ) + ( Xd_0__inst_mult_26_54  ))
// Xd_0__inst_mult_26_57  = CARRY(( !Xd_0__inst_mult_26_8_q  $ (!Xd_0__inst_mult_26_9_q ) ) + ( Xd_0__inst_mult_26_55  ) + ( Xd_0__inst_mult_26_54  ))
// Xd_0__inst_mult_26_58  = SHARE((Xd_0__inst_mult_26_8_q  & Xd_0__inst_mult_26_9_q ))

	.dataa(!Xd_0__inst_mult_26_8_q ),
	.datab(!Xd_0__inst_mult_26_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_54 ),
	.sharein(Xd_0__inst_mult_26_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_56 ),
	.cout(Xd_0__inst_mult_26_57 ),
	.shareout(Xd_0__inst_mult_26_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_27_21 (
// Equation(s):
// Xd_0__inst_mult_27_56  = SUM(( !Xd_0__inst_mult_27_8_q  $ (!Xd_0__inst_mult_27_9_q ) ) + ( Xd_0__inst_mult_27_55  ) + ( Xd_0__inst_mult_27_54  ))
// Xd_0__inst_mult_27_57  = CARRY(( !Xd_0__inst_mult_27_8_q  $ (!Xd_0__inst_mult_27_9_q ) ) + ( Xd_0__inst_mult_27_55  ) + ( Xd_0__inst_mult_27_54  ))
// Xd_0__inst_mult_27_58  = SHARE((Xd_0__inst_mult_27_8_q  & Xd_0__inst_mult_27_9_q ))

	.dataa(!Xd_0__inst_mult_27_8_q ),
	.datab(!Xd_0__inst_mult_27_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_54 ),
	.sharein(Xd_0__inst_mult_27_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_56 ),
	.cout(Xd_0__inst_mult_27_57 ),
	.shareout(Xd_0__inst_mult_27_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_24_21 (
// Equation(s):
// Xd_0__inst_mult_24_56  = SUM(( !Xd_0__inst_mult_24_8_q  $ (!Xd_0__inst_mult_24_9_q ) ) + ( Xd_0__inst_mult_24_55  ) + ( Xd_0__inst_mult_24_54  ))
// Xd_0__inst_mult_24_57  = CARRY(( !Xd_0__inst_mult_24_8_q  $ (!Xd_0__inst_mult_24_9_q ) ) + ( Xd_0__inst_mult_24_55  ) + ( Xd_0__inst_mult_24_54  ))
// Xd_0__inst_mult_24_58  = SHARE((Xd_0__inst_mult_24_8_q  & Xd_0__inst_mult_24_9_q ))

	.dataa(!Xd_0__inst_mult_24_8_q ),
	.datab(!Xd_0__inst_mult_24_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_54 ),
	.sharein(Xd_0__inst_mult_24_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_56 ),
	.cout(Xd_0__inst_mult_24_57 ),
	.shareout(Xd_0__inst_mult_24_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_25_21 (
// Equation(s):
// Xd_0__inst_mult_25_56  = SUM(( !Xd_0__inst_mult_25_8_q  $ (!Xd_0__inst_mult_25_9_q ) ) + ( Xd_0__inst_mult_25_55  ) + ( Xd_0__inst_mult_25_54  ))
// Xd_0__inst_mult_25_57  = CARRY(( !Xd_0__inst_mult_25_8_q  $ (!Xd_0__inst_mult_25_9_q ) ) + ( Xd_0__inst_mult_25_55  ) + ( Xd_0__inst_mult_25_54  ))
// Xd_0__inst_mult_25_58  = SHARE((Xd_0__inst_mult_25_8_q  & Xd_0__inst_mult_25_9_q ))

	.dataa(!Xd_0__inst_mult_25_8_q ),
	.datab(!Xd_0__inst_mult_25_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_54 ),
	.sharein(Xd_0__inst_mult_25_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_56 ),
	.cout(Xd_0__inst_mult_25_57 ),
	.shareout(Xd_0__inst_mult_25_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_22_21 (
// Equation(s):
// Xd_0__inst_mult_22_56  = SUM(( !Xd_0__inst_mult_22_8_q  $ (!Xd_0__inst_mult_22_9_q ) ) + ( Xd_0__inst_mult_22_55  ) + ( Xd_0__inst_mult_22_54  ))
// Xd_0__inst_mult_22_57  = CARRY(( !Xd_0__inst_mult_22_8_q  $ (!Xd_0__inst_mult_22_9_q ) ) + ( Xd_0__inst_mult_22_55  ) + ( Xd_0__inst_mult_22_54  ))
// Xd_0__inst_mult_22_58  = SHARE((Xd_0__inst_mult_22_8_q  & Xd_0__inst_mult_22_9_q ))

	.dataa(!Xd_0__inst_mult_22_8_q ),
	.datab(!Xd_0__inst_mult_22_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_54 ),
	.sharein(Xd_0__inst_mult_22_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_56 ),
	.cout(Xd_0__inst_mult_22_57 ),
	.shareout(Xd_0__inst_mult_22_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_23_21 (
// Equation(s):
// Xd_0__inst_mult_23_56  = SUM(( !Xd_0__inst_mult_23_8_q  $ (!Xd_0__inst_mult_23_9_q ) ) + ( Xd_0__inst_mult_23_55  ) + ( Xd_0__inst_mult_23_54  ))
// Xd_0__inst_mult_23_57  = CARRY(( !Xd_0__inst_mult_23_8_q  $ (!Xd_0__inst_mult_23_9_q ) ) + ( Xd_0__inst_mult_23_55  ) + ( Xd_0__inst_mult_23_54  ))
// Xd_0__inst_mult_23_58  = SHARE((Xd_0__inst_mult_23_8_q  & Xd_0__inst_mult_23_9_q ))

	.dataa(!Xd_0__inst_mult_23_8_q ),
	.datab(!Xd_0__inst_mult_23_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_54 ),
	.sharein(Xd_0__inst_mult_23_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_56 ),
	.cout(Xd_0__inst_mult_23_57 ),
	.shareout(Xd_0__inst_mult_23_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_20_21 (
// Equation(s):
// Xd_0__inst_mult_20_56  = SUM(( !Xd_0__inst_mult_20_8_q  $ (!Xd_0__inst_mult_20_9_q ) ) + ( Xd_0__inst_mult_20_55  ) + ( Xd_0__inst_mult_20_54  ))
// Xd_0__inst_mult_20_57  = CARRY(( !Xd_0__inst_mult_20_8_q  $ (!Xd_0__inst_mult_20_9_q ) ) + ( Xd_0__inst_mult_20_55  ) + ( Xd_0__inst_mult_20_54  ))
// Xd_0__inst_mult_20_58  = SHARE((Xd_0__inst_mult_20_8_q  & Xd_0__inst_mult_20_9_q ))

	.dataa(!Xd_0__inst_mult_20_8_q ),
	.datab(!Xd_0__inst_mult_20_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_54 ),
	.sharein(Xd_0__inst_mult_20_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_56 ),
	.cout(Xd_0__inst_mult_20_57 ),
	.shareout(Xd_0__inst_mult_20_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_21_21 (
// Equation(s):
// Xd_0__inst_mult_21_56  = SUM(( !Xd_0__inst_mult_21_8_q  $ (!Xd_0__inst_mult_21_9_q ) ) + ( Xd_0__inst_mult_21_55  ) + ( Xd_0__inst_mult_21_54  ))
// Xd_0__inst_mult_21_57  = CARRY(( !Xd_0__inst_mult_21_8_q  $ (!Xd_0__inst_mult_21_9_q ) ) + ( Xd_0__inst_mult_21_55  ) + ( Xd_0__inst_mult_21_54  ))
// Xd_0__inst_mult_21_58  = SHARE((Xd_0__inst_mult_21_8_q  & Xd_0__inst_mult_21_9_q ))

	.dataa(!Xd_0__inst_mult_21_8_q ),
	.datab(!Xd_0__inst_mult_21_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_54 ),
	.sharein(Xd_0__inst_mult_21_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_56 ),
	.cout(Xd_0__inst_mult_21_57 ),
	.shareout(Xd_0__inst_mult_21_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_18_21 (
// Equation(s):
// Xd_0__inst_mult_18_56  = SUM(( !Xd_0__inst_mult_18_8_q  $ (!Xd_0__inst_mult_18_9_q ) ) + ( Xd_0__inst_mult_18_55  ) + ( Xd_0__inst_mult_18_54  ))
// Xd_0__inst_mult_18_57  = CARRY(( !Xd_0__inst_mult_18_8_q  $ (!Xd_0__inst_mult_18_9_q ) ) + ( Xd_0__inst_mult_18_55  ) + ( Xd_0__inst_mult_18_54  ))
// Xd_0__inst_mult_18_58  = SHARE((Xd_0__inst_mult_18_8_q  & Xd_0__inst_mult_18_9_q ))

	.dataa(!Xd_0__inst_mult_18_8_q ),
	.datab(!Xd_0__inst_mult_18_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_54 ),
	.sharein(Xd_0__inst_mult_18_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_56 ),
	.cout(Xd_0__inst_mult_18_57 ),
	.shareout(Xd_0__inst_mult_18_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_19_21 (
// Equation(s):
// Xd_0__inst_mult_19_56  = SUM(( !Xd_0__inst_mult_19_8_q  $ (!Xd_0__inst_mult_19_9_q ) ) + ( Xd_0__inst_mult_19_55  ) + ( Xd_0__inst_mult_19_54  ))
// Xd_0__inst_mult_19_57  = CARRY(( !Xd_0__inst_mult_19_8_q  $ (!Xd_0__inst_mult_19_9_q ) ) + ( Xd_0__inst_mult_19_55  ) + ( Xd_0__inst_mult_19_54  ))
// Xd_0__inst_mult_19_58  = SHARE((Xd_0__inst_mult_19_8_q  & Xd_0__inst_mult_19_9_q ))

	.dataa(!Xd_0__inst_mult_19_8_q ),
	.datab(!Xd_0__inst_mult_19_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_54 ),
	.sharein(Xd_0__inst_mult_19_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_56 ),
	.cout(Xd_0__inst_mult_19_57 ),
	.shareout(Xd_0__inst_mult_19_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_16_21 (
// Equation(s):
// Xd_0__inst_mult_16_56  = SUM(( !Xd_0__inst_mult_16_8_q  $ (!Xd_0__inst_mult_16_9_q ) ) + ( Xd_0__inst_mult_16_55  ) + ( Xd_0__inst_mult_16_54  ))
// Xd_0__inst_mult_16_57  = CARRY(( !Xd_0__inst_mult_16_8_q  $ (!Xd_0__inst_mult_16_9_q ) ) + ( Xd_0__inst_mult_16_55  ) + ( Xd_0__inst_mult_16_54  ))
// Xd_0__inst_mult_16_58  = SHARE((Xd_0__inst_mult_16_8_q  & Xd_0__inst_mult_16_9_q ))

	.dataa(!Xd_0__inst_mult_16_8_q ),
	.datab(!Xd_0__inst_mult_16_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_54 ),
	.sharein(Xd_0__inst_mult_16_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_56 ),
	.cout(Xd_0__inst_mult_16_57 ),
	.shareout(Xd_0__inst_mult_16_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_17_21 (
// Equation(s):
// Xd_0__inst_mult_17_56  = SUM(( !Xd_0__inst_mult_17_8_q  $ (!Xd_0__inst_mult_17_9_q ) ) + ( Xd_0__inst_mult_17_55  ) + ( Xd_0__inst_mult_17_54  ))
// Xd_0__inst_mult_17_57  = CARRY(( !Xd_0__inst_mult_17_8_q  $ (!Xd_0__inst_mult_17_9_q ) ) + ( Xd_0__inst_mult_17_55  ) + ( Xd_0__inst_mult_17_54  ))
// Xd_0__inst_mult_17_58  = SHARE((Xd_0__inst_mult_17_8_q  & Xd_0__inst_mult_17_9_q ))

	.dataa(!Xd_0__inst_mult_17_8_q ),
	.datab(!Xd_0__inst_mult_17_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_54 ),
	.sharein(Xd_0__inst_mult_17_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_56 ),
	.cout(Xd_0__inst_mult_17_57 ),
	.shareout(Xd_0__inst_mult_17_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_21 (
// Equation(s):
// Xd_0__inst_mult_14_56  = SUM(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q ) ) + ( Xd_0__inst_mult_14_55  ) + ( Xd_0__inst_mult_14_54  ))
// Xd_0__inst_mult_14_57  = CARRY(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q ) ) + ( Xd_0__inst_mult_14_55  ) + ( Xd_0__inst_mult_14_54  ))
// Xd_0__inst_mult_14_58  = SHARE((Xd_0__inst_mult_14_8_q  & Xd_0__inst_mult_14_9_q ))

	.dataa(!Xd_0__inst_mult_14_8_q ),
	.datab(!Xd_0__inst_mult_14_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_54 ),
	.sharein(Xd_0__inst_mult_14_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_56 ),
	.cout(Xd_0__inst_mult_14_57 ),
	.shareout(Xd_0__inst_mult_14_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_21 (
// Equation(s):
// Xd_0__inst_mult_15_56  = SUM(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q ) ) + ( Xd_0__inst_mult_15_55  ) + ( Xd_0__inst_mult_15_54  ))
// Xd_0__inst_mult_15_57  = CARRY(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q ) ) + ( Xd_0__inst_mult_15_55  ) + ( Xd_0__inst_mult_15_54  ))
// Xd_0__inst_mult_15_58  = SHARE((Xd_0__inst_mult_15_8_q  & Xd_0__inst_mult_15_9_q ))

	.dataa(!Xd_0__inst_mult_15_8_q ),
	.datab(!Xd_0__inst_mult_15_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_54 ),
	.sharein(Xd_0__inst_mult_15_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_56 ),
	.cout(Xd_0__inst_mult_15_57 ),
	.shareout(Xd_0__inst_mult_15_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_21 (
// Equation(s):
// Xd_0__inst_mult_12_56  = SUM(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q ) ) + ( Xd_0__inst_mult_12_55  ) + ( Xd_0__inst_mult_12_54  ))
// Xd_0__inst_mult_12_57  = CARRY(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q ) ) + ( Xd_0__inst_mult_12_55  ) + ( Xd_0__inst_mult_12_54  ))
// Xd_0__inst_mult_12_58  = SHARE((Xd_0__inst_mult_12_8_q  & Xd_0__inst_mult_12_9_q ))

	.dataa(!Xd_0__inst_mult_12_8_q ),
	.datab(!Xd_0__inst_mult_12_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_54 ),
	.sharein(Xd_0__inst_mult_12_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_56 ),
	.cout(Xd_0__inst_mult_12_57 ),
	.shareout(Xd_0__inst_mult_12_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_21 (
// Equation(s):
// Xd_0__inst_mult_13_56  = SUM(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q ) ) + ( Xd_0__inst_mult_13_55  ) + ( Xd_0__inst_mult_13_54  ))
// Xd_0__inst_mult_13_57  = CARRY(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q ) ) + ( Xd_0__inst_mult_13_55  ) + ( Xd_0__inst_mult_13_54  ))
// Xd_0__inst_mult_13_58  = SHARE((Xd_0__inst_mult_13_8_q  & Xd_0__inst_mult_13_9_q ))

	.dataa(!Xd_0__inst_mult_13_8_q ),
	.datab(!Xd_0__inst_mult_13_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_54 ),
	.sharein(Xd_0__inst_mult_13_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_56 ),
	.cout(Xd_0__inst_mult_13_57 ),
	.shareout(Xd_0__inst_mult_13_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_21 (
// Equation(s):
// Xd_0__inst_mult_10_56  = SUM(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q ) ) + ( Xd_0__inst_mult_10_55  ) + ( Xd_0__inst_mult_10_54  ))
// Xd_0__inst_mult_10_57  = CARRY(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q ) ) + ( Xd_0__inst_mult_10_55  ) + ( Xd_0__inst_mult_10_54  ))
// Xd_0__inst_mult_10_58  = SHARE((Xd_0__inst_mult_10_8_q  & Xd_0__inst_mult_10_9_q ))

	.dataa(!Xd_0__inst_mult_10_8_q ),
	.datab(!Xd_0__inst_mult_10_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_54 ),
	.sharein(Xd_0__inst_mult_10_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_56 ),
	.cout(Xd_0__inst_mult_10_57 ),
	.shareout(Xd_0__inst_mult_10_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_21 (
// Equation(s):
// Xd_0__inst_mult_11_56  = SUM(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q ) ) + ( Xd_0__inst_mult_11_55  ) + ( Xd_0__inst_mult_11_54  ))
// Xd_0__inst_mult_11_57  = CARRY(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q ) ) + ( Xd_0__inst_mult_11_55  ) + ( Xd_0__inst_mult_11_54  ))
// Xd_0__inst_mult_11_58  = SHARE((Xd_0__inst_mult_11_8_q  & Xd_0__inst_mult_11_9_q ))

	.dataa(!Xd_0__inst_mult_11_8_q ),
	.datab(!Xd_0__inst_mult_11_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_54 ),
	.sharein(Xd_0__inst_mult_11_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_56 ),
	.cout(Xd_0__inst_mult_11_57 ),
	.shareout(Xd_0__inst_mult_11_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_21 (
// Equation(s):
// Xd_0__inst_mult_8_56  = SUM(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q ) ) + ( Xd_0__inst_mult_8_55  ) + ( Xd_0__inst_mult_8_54  ))
// Xd_0__inst_mult_8_57  = CARRY(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q ) ) + ( Xd_0__inst_mult_8_55  ) + ( Xd_0__inst_mult_8_54  ))
// Xd_0__inst_mult_8_58  = SHARE((Xd_0__inst_mult_8_8_q  & Xd_0__inst_mult_8_9_q ))

	.dataa(!Xd_0__inst_mult_8_8_q ),
	.datab(!Xd_0__inst_mult_8_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_54 ),
	.sharein(Xd_0__inst_mult_8_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_56 ),
	.cout(Xd_0__inst_mult_8_57 ),
	.shareout(Xd_0__inst_mult_8_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_21 (
// Equation(s):
// Xd_0__inst_mult_9_56  = SUM(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q ) ) + ( Xd_0__inst_mult_9_55  ) + ( Xd_0__inst_mult_9_54  ))
// Xd_0__inst_mult_9_57  = CARRY(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q ) ) + ( Xd_0__inst_mult_9_55  ) + ( Xd_0__inst_mult_9_54  ))
// Xd_0__inst_mult_9_58  = SHARE((Xd_0__inst_mult_9_8_q  & Xd_0__inst_mult_9_9_q ))

	.dataa(!Xd_0__inst_mult_9_8_q ),
	.datab(!Xd_0__inst_mult_9_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_54 ),
	.sharein(Xd_0__inst_mult_9_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_56 ),
	.cout(Xd_0__inst_mult_9_57 ),
	.shareout(Xd_0__inst_mult_9_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_21 (
// Equation(s):
// Xd_0__inst_mult_6_56  = SUM(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_55  ) + ( Xd_0__inst_mult_6_54  ))
// Xd_0__inst_mult_6_57  = CARRY(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_55  ) + ( Xd_0__inst_mult_6_54  ))
// Xd_0__inst_mult_6_58  = SHARE((Xd_0__inst_mult_6_8_q  & Xd_0__inst_mult_6_9_q ))

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_54 ),
	.sharein(Xd_0__inst_mult_6_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_56 ),
	.cout(Xd_0__inst_mult_6_57 ),
	.shareout(Xd_0__inst_mult_6_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_21 (
// Equation(s):
// Xd_0__inst_mult_7_56  = SUM(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_55  ) + ( Xd_0__inst_mult_7_54  ))
// Xd_0__inst_mult_7_57  = CARRY(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_55  ) + ( Xd_0__inst_mult_7_54  ))
// Xd_0__inst_mult_7_58  = SHARE((Xd_0__inst_mult_7_8_q  & Xd_0__inst_mult_7_9_q ))

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_54 ),
	.sharein(Xd_0__inst_mult_7_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_56 ),
	.cout(Xd_0__inst_mult_7_57 ),
	.shareout(Xd_0__inst_mult_7_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_21 (
// Equation(s):
// Xd_0__inst_mult_4_56  = SUM(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_55  ) + ( Xd_0__inst_mult_4_54  ))
// Xd_0__inst_mult_4_57  = CARRY(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_55  ) + ( Xd_0__inst_mult_4_54  ))
// Xd_0__inst_mult_4_58  = SHARE((Xd_0__inst_mult_4_8_q  & Xd_0__inst_mult_4_9_q ))

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_54 ),
	.sharein(Xd_0__inst_mult_4_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_56 ),
	.cout(Xd_0__inst_mult_4_57 ),
	.shareout(Xd_0__inst_mult_4_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_21 (
// Equation(s):
// Xd_0__inst_mult_5_56  = SUM(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_55  ) + ( Xd_0__inst_mult_5_54  ))
// Xd_0__inst_mult_5_57  = CARRY(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_55  ) + ( Xd_0__inst_mult_5_54  ))
// Xd_0__inst_mult_5_58  = SHARE((Xd_0__inst_mult_5_8_q  & Xd_0__inst_mult_5_9_q ))

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_54 ),
	.sharein(Xd_0__inst_mult_5_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_56 ),
	.cout(Xd_0__inst_mult_5_57 ),
	.shareout(Xd_0__inst_mult_5_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_21 (
// Equation(s):
// Xd_0__inst_mult_2_56  = SUM(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_55  ) + ( Xd_0__inst_mult_2_54  ))
// Xd_0__inst_mult_2_57  = CARRY(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_55  ) + ( Xd_0__inst_mult_2_54  ))
// Xd_0__inst_mult_2_58  = SHARE((Xd_0__inst_mult_2_8_q  & Xd_0__inst_mult_2_9_q ))

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_54 ),
	.sharein(Xd_0__inst_mult_2_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_56 ),
	.cout(Xd_0__inst_mult_2_57 ),
	.shareout(Xd_0__inst_mult_2_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_21 (
// Equation(s):
// Xd_0__inst_mult_3_56  = SUM(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_55  ) + ( Xd_0__inst_mult_3_54  ))
// Xd_0__inst_mult_3_57  = CARRY(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_55  ) + ( Xd_0__inst_mult_3_54  ))
// Xd_0__inst_mult_3_58  = SHARE((Xd_0__inst_mult_3_8_q  & Xd_0__inst_mult_3_9_q ))

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_54 ),
	.sharein(Xd_0__inst_mult_3_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_56 ),
	.cout(Xd_0__inst_mult_3_57 ),
	.shareout(Xd_0__inst_mult_3_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_21 (
// Equation(s):
// Xd_0__inst_mult_0_56  = SUM(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_55  ) + ( Xd_0__inst_mult_0_54  ))
// Xd_0__inst_mult_0_57  = CARRY(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_55  ) + ( Xd_0__inst_mult_0_54  ))
// Xd_0__inst_mult_0_58  = SHARE((Xd_0__inst_mult_0_8_q  & Xd_0__inst_mult_0_9_q ))

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_54 ),
	.sharein(Xd_0__inst_mult_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_56 ),
	.cout(Xd_0__inst_mult_0_57 ),
	.shareout(Xd_0__inst_mult_0_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_21 (
// Equation(s):
// Xd_0__inst_mult_1_56  = SUM(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_55  ) + ( Xd_0__inst_mult_1_54  ))
// Xd_0__inst_mult_1_57  = CARRY(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_55  ) + ( Xd_0__inst_mult_1_54  ))
// Xd_0__inst_mult_1_58  = SHARE((Xd_0__inst_mult_1_8_q  & Xd_0__inst_mult_1_9_q ))

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_54 ),
	.sharein(Xd_0__inst_mult_1_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_56 ),
	.cout(Xd_0__inst_mult_1_57 ),
	.shareout(Xd_0__inst_mult_1_58 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_28_22 (
// Equation(s):
// Xd_0__inst_mult_28_60  = SUM(( !Xd_0__inst_mult_28_10_q  $ (!Xd_0__inst_mult_28_11_q  $ (((Xd_0__inst_mult_28_2_q  & Xd_0__inst_mult_28_1_q )))) ) + ( Xd_0__inst_mult_28_58  ) + ( Xd_0__inst_mult_28_57  ))
// Xd_0__inst_mult_28_61  = CARRY(( !Xd_0__inst_mult_28_10_q  $ (!Xd_0__inst_mult_28_11_q  $ (((Xd_0__inst_mult_28_2_q  & Xd_0__inst_mult_28_1_q )))) ) + ( Xd_0__inst_mult_28_58  ) + ( Xd_0__inst_mult_28_57  ))
// Xd_0__inst_mult_28_62  = SHARE((!Xd_0__inst_mult_28_10_q  & (Xd_0__inst_mult_28_11_q  & (Xd_0__inst_mult_28_2_q  & Xd_0__inst_mult_28_1_q ))) # (Xd_0__inst_mult_28_10_q  & (((Xd_0__inst_mult_28_2_q  & Xd_0__inst_mult_28_1_q )) # (Xd_0__inst_mult_28_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_28_10_q ),
	.datab(!Xd_0__inst_mult_28_11_q ),
	.datac(!Xd_0__inst_mult_28_2_q ),
	.datad(!Xd_0__inst_mult_28_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_57 ),
	.sharein(Xd_0__inst_mult_28_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_60 ),
	.cout(Xd_0__inst_mult_28_61 ),
	.shareout(Xd_0__inst_mult_28_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_29_22 (
// Equation(s):
// Xd_0__inst_mult_29_60  = SUM(( !Xd_0__inst_mult_29_10_q  $ (!Xd_0__inst_mult_29_11_q  $ (((Xd_0__inst_mult_29_2_q  & Xd_0__inst_mult_29_1_q )))) ) + ( Xd_0__inst_mult_29_58  ) + ( Xd_0__inst_mult_29_57  ))
// Xd_0__inst_mult_29_61  = CARRY(( !Xd_0__inst_mult_29_10_q  $ (!Xd_0__inst_mult_29_11_q  $ (((Xd_0__inst_mult_29_2_q  & Xd_0__inst_mult_29_1_q )))) ) + ( Xd_0__inst_mult_29_58  ) + ( Xd_0__inst_mult_29_57  ))
// Xd_0__inst_mult_29_62  = SHARE((!Xd_0__inst_mult_29_10_q  & (Xd_0__inst_mult_29_11_q  & (Xd_0__inst_mult_29_2_q  & Xd_0__inst_mult_29_1_q ))) # (Xd_0__inst_mult_29_10_q  & (((Xd_0__inst_mult_29_2_q  & Xd_0__inst_mult_29_1_q )) # (Xd_0__inst_mult_29_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_29_10_q ),
	.datab(!Xd_0__inst_mult_29_11_q ),
	.datac(!Xd_0__inst_mult_29_2_q ),
	.datad(!Xd_0__inst_mult_29_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_57 ),
	.sharein(Xd_0__inst_mult_29_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_60 ),
	.cout(Xd_0__inst_mult_29_61 ),
	.shareout(Xd_0__inst_mult_29_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_26_22 (
// Equation(s):
// Xd_0__inst_mult_26_60  = SUM(( !Xd_0__inst_mult_26_10_q  $ (!Xd_0__inst_mult_26_11_q  $ (((Xd_0__inst_mult_26_2_q  & Xd_0__inst_mult_26_1_q )))) ) + ( Xd_0__inst_mult_26_58  ) + ( Xd_0__inst_mult_26_57  ))
// Xd_0__inst_mult_26_61  = CARRY(( !Xd_0__inst_mult_26_10_q  $ (!Xd_0__inst_mult_26_11_q  $ (((Xd_0__inst_mult_26_2_q  & Xd_0__inst_mult_26_1_q )))) ) + ( Xd_0__inst_mult_26_58  ) + ( Xd_0__inst_mult_26_57  ))
// Xd_0__inst_mult_26_62  = SHARE((!Xd_0__inst_mult_26_10_q  & (Xd_0__inst_mult_26_11_q  & (Xd_0__inst_mult_26_2_q  & Xd_0__inst_mult_26_1_q ))) # (Xd_0__inst_mult_26_10_q  & (((Xd_0__inst_mult_26_2_q  & Xd_0__inst_mult_26_1_q )) # (Xd_0__inst_mult_26_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_26_10_q ),
	.datab(!Xd_0__inst_mult_26_11_q ),
	.datac(!Xd_0__inst_mult_26_2_q ),
	.datad(!Xd_0__inst_mult_26_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_57 ),
	.sharein(Xd_0__inst_mult_26_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_60 ),
	.cout(Xd_0__inst_mult_26_61 ),
	.shareout(Xd_0__inst_mult_26_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_27_22 (
// Equation(s):
// Xd_0__inst_mult_27_60  = SUM(( !Xd_0__inst_mult_27_10_q  $ (!Xd_0__inst_mult_27_11_q  $ (((Xd_0__inst_mult_27_2_q  & Xd_0__inst_mult_27_1_q )))) ) + ( Xd_0__inst_mult_27_58  ) + ( Xd_0__inst_mult_27_57  ))
// Xd_0__inst_mult_27_61  = CARRY(( !Xd_0__inst_mult_27_10_q  $ (!Xd_0__inst_mult_27_11_q  $ (((Xd_0__inst_mult_27_2_q  & Xd_0__inst_mult_27_1_q )))) ) + ( Xd_0__inst_mult_27_58  ) + ( Xd_0__inst_mult_27_57  ))
// Xd_0__inst_mult_27_62  = SHARE((!Xd_0__inst_mult_27_10_q  & (Xd_0__inst_mult_27_11_q  & (Xd_0__inst_mult_27_2_q  & Xd_0__inst_mult_27_1_q ))) # (Xd_0__inst_mult_27_10_q  & (((Xd_0__inst_mult_27_2_q  & Xd_0__inst_mult_27_1_q )) # (Xd_0__inst_mult_27_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_27_10_q ),
	.datab(!Xd_0__inst_mult_27_11_q ),
	.datac(!Xd_0__inst_mult_27_2_q ),
	.datad(!Xd_0__inst_mult_27_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_57 ),
	.sharein(Xd_0__inst_mult_27_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_60 ),
	.cout(Xd_0__inst_mult_27_61 ),
	.shareout(Xd_0__inst_mult_27_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_24_22 (
// Equation(s):
// Xd_0__inst_mult_24_60  = SUM(( !Xd_0__inst_mult_24_10_q  $ (!Xd_0__inst_mult_24_11_q  $ (((Xd_0__inst_mult_24_2_q  & Xd_0__inst_mult_24_1_q )))) ) + ( Xd_0__inst_mult_24_58  ) + ( Xd_0__inst_mult_24_57  ))
// Xd_0__inst_mult_24_61  = CARRY(( !Xd_0__inst_mult_24_10_q  $ (!Xd_0__inst_mult_24_11_q  $ (((Xd_0__inst_mult_24_2_q  & Xd_0__inst_mult_24_1_q )))) ) + ( Xd_0__inst_mult_24_58  ) + ( Xd_0__inst_mult_24_57  ))
// Xd_0__inst_mult_24_62  = SHARE((!Xd_0__inst_mult_24_10_q  & (Xd_0__inst_mult_24_11_q  & (Xd_0__inst_mult_24_2_q  & Xd_0__inst_mult_24_1_q ))) # (Xd_0__inst_mult_24_10_q  & (((Xd_0__inst_mult_24_2_q  & Xd_0__inst_mult_24_1_q )) # (Xd_0__inst_mult_24_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_24_10_q ),
	.datab(!Xd_0__inst_mult_24_11_q ),
	.datac(!Xd_0__inst_mult_24_2_q ),
	.datad(!Xd_0__inst_mult_24_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_57 ),
	.sharein(Xd_0__inst_mult_24_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_60 ),
	.cout(Xd_0__inst_mult_24_61 ),
	.shareout(Xd_0__inst_mult_24_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_25_22 (
// Equation(s):
// Xd_0__inst_mult_25_60  = SUM(( !Xd_0__inst_mult_25_10_q  $ (!Xd_0__inst_mult_25_11_q  $ (((Xd_0__inst_mult_25_2_q  & Xd_0__inst_mult_25_1_q )))) ) + ( Xd_0__inst_mult_25_58  ) + ( Xd_0__inst_mult_25_57  ))
// Xd_0__inst_mult_25_61  = CARRY(( !Xd_0__inst_mult_25_10_q  $ (!Xd_0__inst_mult_25_11_q  $ (((Xd_0__inst_mult_25_2_q  & Xd_0__inst_mult_25_1_q )))) ) + ( Xd_0__inst_mult_25_58  ) + ( Xd_0__inst_mult_25_57  ))
// Xd_0__inst_mult_25_62  = SHARE((!Xd_0__inst_mult_25_10_q  & (Xd_0__inst_mult_25_11_q  & (Xd_0__inst_mult_25_2_q  & Xd_0__inst_mult_25_1_q ))) # (Xd_0__inst_mult_25_10_q  & (((Xd_0__inst_mult_25_2_q  & Xd_0__inst_mult_25_1_q )) # (Xd_0__inst_mult_25_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_25_10_q ),
	.datab(!Xd_0__inst_mult_25_11_q ),
	.datac(!Xd_0__inst_mult_25_2_q ),
	.datad(!Xd_0__inst_mult_25_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_57 ),
	.sharein(Xd_0__inst_mult_25_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_60 ),
	.cout(Xd_0__inst_mult_25_61 ),
	.shareout(Xd_0__inst_mult_25_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_22_22 (
// Equation(s):
// Xd_0__inst_mult_22_60  = SUM(( !Xd_0__inst_mult_22_10_q  $ (!Xd_0__inst_mult_22_11_q  $ (((Xd_0__inst_mult_22_2_q  & Xd_0__inst_mult_22_1_q )))) ) + ( Xd_0__inst_mult_22_58  ) + ( Xd_0__inst_mult_22_57  ))
// Xd_0__inst_mult_22_61  = CARRY(( !Xd_0__inst_mult_22_10_q  $ (!Xd_0__inst_mult_22_11_q  $ (((Xd_0__inst_mult_22_2_q  & Xd_0__inst_mult_22_1_q )))) ) + ( Xd_0__inst_mult_22_58  ) + ( Xd_0__inst_mult_22_57  ))
// Xd_0__inst_mult_22_62  = SHARE((!Xd_0__inst_mult_22_10_q  & (Xd_0__inst_mult_22_11_q  & (Xd_0__inst_mult_22_2_q  & Xd_0__inst_mult_22_1_q ))) # (Xd_0__inst_mult_22_10_q  & (((Xd_0__inst_mult_22_2_q  & Xd_0__inst_mult_22_1_q )) # (Xd_0__inst_mult_22_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_22_10_q ),
	.datab(!Xd_0__inst_mult_22_11_q ),
	.datac(!Xd_0__inst_mult_22_2_q ),
	.datad(!Xd_0__inst_mult_22_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_57 ),
	.sharein(Xd_0__inst_mult_22_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_60 ),
	.cout(Xd_0__inst_mult_22_61 ),
	.shareout(Xd_0__inst_mult_22_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_23_22 (
// Equation(s):
// Xd_0__inst_mult_23_60  = SUM(( !Xd_0__inst_mult_23_10_q  $ (!Xd_0__inst_mult_23_11_q  $ (((Xd_0__inst_mult_23_2_q  & Xd_0__inst_mult_23_1_q )))) ) + ( Xd_0__inst_mult_23_58  ) + ( Xd_0__inst_mult_23_57  ))
// Xd_0__inst_mult_23_61  = CARRY(( !Xd_0__inst_mult_23_10_q  $ (!Xd_0__inst_mult_23_11_q  $ (((Xd_0__inst_mult_23_2_q  & Xd_0__inst_mult_23_1_q )))) ) + ( Xd_0__inst_mult_23_58  ) + ( Xd_0__inst_mult_23_57  ))
// Xd_0__inst_mult_23_62  = SHARE((!Xd_0__inst_mult_23_10_q  & (Xd_0__inst_mult_23_11_q  & (Xd_0__inst_mult_23_2_q  & Xd_0__inst_mult_23_1_q ))) # (Xd_0__inst_mult_23_10_q  & (((Xd_0__inst_mult_23_2_q  & Xd_0__inst_mult_23_1_q )) # (Xd_0__inst_mult_23_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_23_10_q ),
	.datab(!Xd_0__inst_mult_23_11_q ),
	.datac(!Xd_0__inst_mult_23_2_q ),
	.datad(!Xd_0__inst_mult_23_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_57 ),
	.sharein(Xd_0__inst_mult_23_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_60 ),
	.cout(Xd_0__inst_mult_23_61 ),
	.shareout(Xd_0__inst_mult_23_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_20_22 (
// Equation(s):
// Xd_0__inst_mult_20_60  = SUM(( !Xd_0__inst_mult_20_10_q  $ (!Xd_0__inst_mult_20_11_q  $ (((Xd_0__inst_mult_20_2_q  & Xd_0__inst_mult_20_1_q )))) ) + ( Xd_0__inst_mult_20_58  ) + ( Xd_0__inst_mult_20_57  ))
// Xd_0__inst_mult_20_61  = CARRY(( !Xd_0__inst_mult_20_10_q  $ (!Xd_0__inst_mult_20_11_q  $ (((Xd_0__inst_mult_20_2_q  & Xd_0__inst_mult_20_1_q )))) ) + ( Xd_0__inst_mult_20_58  ) + ( Xd_0__inst_mult_20_57  ))
// Xd_0__inst_mult_20_62  = SHARE((!Xd_0__inst_mult_20_10_q  & (Xd_0__inst_mult_20_11_q  & (Xd_0__inst_mult_20_2_q  & Xd_0__inst_mult_20_1_q ))) # (Xd_0__inst_mult_20_10_q  & (((Xd_0__inst_mult_20_2_q  & Xd_0__inst_mult_20_1_q )) # (Xd_0__inst_mult_20_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_20_10_q ),
	.datab(!Xd_0__inst_mult_20_11_q ),
	.datac(!Xd_0__inst_mult_20_2_q ),
	.datad(!Xd_0__inst_mult_20_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_57 ),
	.sharein(Xd_0__inst_mult_20_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_60 ),
	.cout(Xd_0__inst_mult_20_61 ),
	.shareout(Xd_0__inst_mult_20_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_21_22 (
// Equation(s):
// Xd_0__inst_mult_21_60  = SUM(( !Xd_0__inst_mult_21_10_q  $ (!Xd_0__inst_mult_21_11_q  $ (((Xd_0__inst_mult_21_2_q  & Xd_0__inst_mult_21_1_q )))) ) + ( Xd_0__inst_mult_21_58  ) + ( Xd_0__inst_mult_21_57  ))
// Xd_0__inst_mult_21_61  = CARRY(( !Xd_0__inst_mult_21_10_q  $ (!Xd_0__inst_mult_21_11_q  $ (((Xd_0__inst_mult_21_2_q  & Xd_0__inst_mult_21_1_q )))) ) + ( Xd_0__inst_mult_21_58  ) + ( Xd_0__inst_mult_21_57  ))
// Xd_0__inst_mult_21_62  = SHARE((!Xd_0__inst_mult_21_10_q  & (Xd_0__inst_mult_21_11_q  & (Xd_0__inst_mult_21_2_q  & Xd_0__inst_mult_21_1_q ))) # (Xd_0__inst_mult_21_10_q  & (((Xd_0__inst_mult_21_2_q  & Xd_0__inst_mult_21_1_q )) # (Xd_0__inst_mult_21_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_21_10_q ),
	.datab(!Xd_0__inst_mult_21_11_q ),
	.datac(!Xd_0__inst_mult_21_2_q ),
	.datad(!Xd_0__inst_mult_21_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_57 ),
	.sharein(Xd_0__inst_mult_21_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_60 ),
	.cout(Xd_0__inst_mult_21_61 ),
	.shareout(Xd_0__inst_mult_21_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_18_22 (
// Equation(s):
// Xd_0__inst_mult_18_60  = SUM(( !Xd_0__inst_mult_18_10_q  $ (!Xd_0__inst_mult_18_11_q  $ (((Xd_0__inst_mult_18_2_q  & Xd_0__inst_mult_18_1_q )))) ) + ( Xd_0__inst_mult_18_58  ) + ( Xd_0__inst_mult_18_57  ))
// Xd_0__inst_mult_18_61  = CARRY(( !Xd_0__inst_mult_18_10_q  $ (!Xd_0__inst_mult_18_11_q  $ (((Xd_0__inst_mult_18_2_q  & Xd_0__inst_mult_18_1_q )))) ) + ( Xd_0__inst_mult_18_58  ) + ( Xd_0__inst_mult_18_57  ))
// Xd_0__inst_mult_18_62  = SHARE((!Xd_0__inst_mult_18_10_q  & (Xd_0__inst_mult_18_11_q  & (Xd_0__inst_mult_18_2_q  & Xd_0__inst_mult_18_1_q ))) # (Xd_0__inst_mult_18_10_q  & (((Xd_0__inst_mult_18_2_q  & Xd_0__inst_mult_18_1_q )) # (Xd_0__inst_mult_18_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_18_10_q ),
	.datab(!Xd_0__inst_mult_18_11_q ),
	.datac(!Xd_0__inst_mult_18_2_q ),
	.datad(!Xd_0__inst_mult_18_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_57 ),
	.sharein(Xd_0__inst_mult_18_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_60 ),
	.cout(Xd_0__inst_mult_18_61 ),
	.shareout(Xd_0__inst_mult_18_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_19_22 (
// Equation(s):
// Xd_0__inst_mult_19_60  = SUM(( !Xd_0__inst_mult_19_10_q  $ (!Xd_0__inst_mult_19_11_q  $ (((Xd_0__inst_mult_19_2_q  & Xd_0__inst_mult_19_1_q )))) ) + ( Xd_0__inst_mult_19_58  ) + ( Xd_0__inst_mult_19_57  ))
// Xd_0__inst_mult_19_61  = CARRY(( !Xd_0__inst_mult_19_10_q  $ (!Xd_0__inst_mult_19_11_q  $ (((Xd_0__inst_mult_19_2_q  & Xd_0__inst_mult_19_1_q )))) ) + ( Xd_0__inst_mult_19_58  ) + ( Xd_0__inst_mult_19_57  ))
// Xd_0__inst_mult_19_62  = SHARE((!Xd_0__inst_mult_19_10_q  & (Xd_0__inst_mult_19_11_q  & (Xd_0__inst_mult_19_2_q  & Xd_0__inst_mult_19_1_q ))) # (Xd_0__inst_mult_19_10_q  & (((Xd_0__inst_mult_19_2_q  & Xd_0__inst_mult_19_1_q )) # (Xd_0__inst_mult_19_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_19_10_q ),
	.datab(!Xd_0__inst_mult_19_11_q ),
	.datac(!Xd_0__inst_mult_19_2_q ),
	.datad(!Xd_0__inst_mult_19_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_57 ),
	.sharein(Xd_0__inst_mult_19_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_60 ),
	.cout(Xd_0__inst_mult_19_61 ),
	.shareout(Xd_0__inst_mult_19_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_16_22 (
// Equation(s):
// Xd_0__inst_mult_16_60  = SUM(( !Xd_0__inst_mult_16_10_q  $ (!Xd_0__inst_mult_16_11_q  $ (((Xd_0__inst_mult_16_2_q  & Xd_0__inst_mult_16_1_q )))) ) + ( Xd_0__inst_mult_16_58  ) + ( Xd_0__inst_mult_16_57  ))
// Xd_0__inst_mult_16_61  = CARRY(( !Xd_0__inst_mult_16_10_q  $ (!Xd_0__inst_mult_16_11_q  $ (((Xd_0__inst_mult_16_2_q  & Xd_0__inst_mult_16_1_q )))) ) + ( Xd_0__inst_mult_16_58  ) + ( Xd_0__inst_mult_16_57  ))
// Xd_0__inst_mult_16_62  = SHARE((!Xd_0__inst_mult_16_10_q  & (Xd_0__inst_mult_16_11_q  & (Xd_0__inst_mult_16_2_q  & Xd_0__inst_mult_16_1_q ))) # (Xd_0__inst_mult_16_10_q  & (((Xd_0__inst_mult_16_2_q  & Xd_0__inst_mult_16_1_q )) # (Xd_0__inst_mult_16_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_16_10_q ),
	.datab(!Xd_0__inst_mult_16_11_q ),
	.datac(!Xd_0__inst_mult_16_2_q ),
	.datad(!Xd_0__inst_mult_16_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_57 ),
	.sharein(Xd_0__inst_mult_16_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_60 ),
	.cout(Xd_0__inst_mult_16_61 ),
	.shareout(Xd_0__inst_mult_16_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_17_22 (
// Equation(s):
// Xd_0__inst_mult_17_60  = SUM(( !Xd_0__inst_mult_17_10_q  $ (!Xd_0__inst_mult_17_11_q  $ (((Xd_0__inst_mult_17_2_q  & Xd_0__inst_mult_17_1_q )))) ) + ( Xd_0__inst_mult_17_58  ) + ( Xd_0__inst_mult_17_57  ))
// Xd_0__inst_mult_17_61  = CARRY(( !Xd_0__inst_mult_17_10_q  $ (!Xd_0__inst_mult_17_11_q  $ (((Xd_0__inst_mult_17_2_q  & Xd_0__inst_mult_17_1_q )))) ) + ( Xd_0__inst_mult_17_58  ) + ( Xd_0__inst_mult_17_57  ))
// Xd_0__inst_mult_17_62  = SHARE((!Xd_0__inst_mult_17_10_q  & (Xd_0__inst_mult_17_11_q  & (Xd_0__inst_mult_17_2_q  & Xd_0__inst_mult_17_1_q ))) # (Xd_0__inst_mult_17_10_q  & (((Xd_0__inst_mult_17_2_q  & Xd_0__inst_mult_17_1_q )) # (Xd_0__inst_mult_17_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_17_10_q ),
	.datab(!Xd_0__inst_mult_17_11_q ),
	.datac(!Xd_0__inst_mult_17_2_q ),
	.datad(!Xd_0__inst_mult_17_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_57 ),
	.sharein(Xd_0__inst_mult_17_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_60 ),
	.cout(Xd_0__inst_mult_17_61 ),
	.shareout(Xd_0__inst_mult_17_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_22 (
// Equation(s):
// Xd_0__inst_mult_14_60  = SUM(( !Xd_0__inst_mult_14_10_q  $ (!Xd_0__inst_mult_14_11_q  $ (((Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_1_q )))) ) + ( Xd_0__inst_mult_14_58  ) + ( Xd_0__inst_mult_14_57  ))
// Xd_0__inst_mult_14_61  = CARRY(( !Xd_0__inst_mult_14_10_q  $ (!Xd_0__inst_mult_14_11_q  $ (((Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_1_q )))) ) + ( Xd_0__inst_mult_14_58  ) + ( Xd_0__inst_mult_14_57  ))
// Xd_0__inst_mult_14_62  = SHARE((!Xd_0__inst_mult_14_10_q  & (Xd_0__inst_mult_14_11_q  & (Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_1_q ))) # (Xd_0__inst_mult_14_10_q  & (((Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_1_q )) # (Xd_0__inst_mult_14_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_14_10_q ),
	.datab(!Xd_0__inst_mult_14_11_q ),
	.datac(!Xd_0__inst_mult_14_2_q ),
	.datad(!Xd_0__inst_mult_14_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_57 ),
	.sharein(Xd_0__inst_mult_14_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_60 ),
	.cout(Xd_0__inst_mult_14_61 ),
	.shareout(Xd_0__inst_mult_14_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_22 (
// Equation(s):
// Xd_0__inst_mult_15_60  = SUM(( !Xd_0__inst_mult_15_10_q  $ (!Xd_0__inst_mult_15_11_q  $ (((Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_1_q )))) ) + ( Xd_0__inst_mult_15_58  ) + ( Xd_0__inst_mult_15_57  ))
// Xd_0__inst_mult_15_61  = CARRY(( !Xd_0__inst_mult_15_10_q  $ (!Xd_0__inst_mult_15_11_q  $ (((Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_1_q )))) ) + ( Xd_0__inst_mult_15_58  ) + ( Xd_0__inst_mult_15_57  ))
// Xd_0__inst_mult_15_62  = SHARE((!Xd_0__inst_mult_15_10_q  & (Xd_0__inst_mult_15_11_q  & (Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_1_q ))) # (Xd_0__inst_mult_15_10_q  & (((Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_1_q )) # (Xd_0__inst_mult_15_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_15_10_q ),
	.datab(!Xd_0__inst_mult_15_11_q ),
	.datac(!Xd_0__inst_mult_15_2_q ),
	.datad(!Xd_0__inst_mult_15_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_57 ),
	.sharein(Xd_0__inst_mult_15_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_60 ),
	.cout(Xd_0__inst_mult_15_61 ),
	.shareout(Xd_0__inst_mult_15_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_22 (
// Equation(s):
// Xd_0__inst_mult_12_60  = SUM(( !Xd_0__inst_mult_12_10_q  $ (!Xd_0__inst_mult_12_11_q  $ (((Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_1_q )))) ) + ( Xd_0__inst_mult_12_58  ) + ( Xd_0__inst_mult_12_57  ))
// Xd_0__inst_mult_12_61  = CARRY(( !Xd_0__inst_mult_12_10_q  $ (!Xd_0__inst_mult_12_11_q  $ (((Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_1_q )))) ) + ( Xd_0__inst_mult_12_58  ) + ( Xd_0__inst_mult_12_57  ))
// Xd_0__inst_mult_12_62  = SHARE((!Xd_0__inst_mult_12_10_q  & (Xd_0__inst_mult_12_11_q  & (Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_1_q ))) # (Xd_0__inst_mult_12_10_q  & (((Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_1_q )) # (Xd_0__inst_mult_12_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_12_10_q ),
	.datab(!Xd_0__inst_mult_12_11_q ),
	.datac(!Xd_0__inst_mult_12_2_q ),
	.datad(!Xd_0__inst_mult_12_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_57 ),
	.sharein(Xd_0__inst_mult_12_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_60 ),
	.cout(Xd_0__inst_mult_12_61 ),
	.shareout(Xd_0__inst_mult_12_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_22 (
// Equation(s):
// Xd_0__inst_mult_13_60  = SUM(( !Xd_0__inst_mult_13_10_q  $ (!Xd_0__inst_mult_13_11_q  $ (((Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_1_q )))) ) + ( Xd_0__inst_mult_13_58  ) + ( Xd_0__inst_mult_13_57  ))
// Xd_0__inst_mult_13_61  = CARRY(( !Xd_0__inst_mult_13_10_q  $ (!Xd_0__inst_mult_13_11_q  $ (((Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_1_q )))) ) + ( Xd_0__inst_mult_13_58  ) + ( Xd_0__inst_mult_13_57  ))
// Xd_0__inst_mult_13_62  = SHARE((!Xd_0__inst_mult_13_10_q  & (Xd_0__inst_mult_13_11_q  & (Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_1_q ))) # (Xd_0__inst_mult_13_10_q  & (((Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_1_q )) # (Xd_0__inst_mult_13_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_13_10_q ),
	.datab(!Xd_0__inst_mult_13_11_q ),
	.datac(!Xd_0__inst_mult_13_2_q ),
	.datad(!Xd_0__inst_mult_13_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_57 ),
	.sharein(Xd_0__inst_mult_13_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_60 ),
	.cout(Xd_0__inst_mult_13_61 ),
	.shareout(Xd_0__inst_mult_13_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_22 (
// Equation(s):
// Xd_0__inst_mult_10_60  = SUM(( !Xd_0__inst_mult_10_10_q  $ (!Xd_0__inst_mult_10_11_q  $ (((Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_1_q )))) ) + ( Xd_0__inst_mult_10_58  ) + ( Xd_0__inst_mult_10_57  ))
// Xd_0__inst_mult_10_61  = CARRY(( !Xd_0__inst_mult_10_10_q  $ (!Xd_0__inst_mult_10_11_q  $ (((Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_1_q )))) ) + ( Xd_0__inst_mult_10_58  ) + ( Xd_0__inst_mult_10_57  ))
// Xd_0__inst_mult_10_62  = SHARE((!Xd_0__inst_mult_10_10_q  & (Xd_0__inst_mult_10_11_q  & (Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_1_q ))) # (Xd_0__inst_mult_10_10_q  & (((Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_1_q )) # (Xd_0__inst_mult_10_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_10_10_q ),
	.datab(!Xd_0__inst_mult_10_11_q ),
	.datac(!Xd_0__inst_mult_10_2_q ),
	.datad(!Xd_0__inst_mult_10_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_57 ),
	.sharein(Xd_0__inst_mult_10_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_60 ),
	.cout(Xd_0__inst_mult_10_61 ),
	.shareout(Xd_0__inst_mult_10_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_22 (
// Equation(s):
// Xd_0__inst_mult_11_60  = SUM(( !Xd_0__inst_mult_11_10_q  $ (!Xd_0__inst_mult_11_11_q  $ (((Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_1_q )))) ) + ( Xd_0__inst_mult_11_58  ) + ( Xd_0__inst_mult_11_57  ))
// Xd_0__inst_mult_11_61  = CARRY(( !Xd_0__inst_mult_11_10_q  $ (!Xd_0__inst_mult_11_11_q  $ (((Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_1_q )))) ) + ( Xd_0__inst_mult_11_58  ) + ( Xd_0__inst_mult_11_57  ))
// Xd_0__inst_mult_11_62  = SHARE((!Xd_0__inst_mult_11_10_q  & (Xd_0__inst_mult_11_11_q  & (Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_1_q ))) # (Xd_0__inst_mult_11_10_q  & (((Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_1_q )) # (Xd_0__inst_mult_11_11_q 
// ))))

	.dataa(!Xd_0__inst_mult_11_10_q ),
	.datab(!Xd_0__inst_mult_11_11_q ),
	.datac(!Xd_0__inst_mult_11_2_q ),
	.datad(!Xd_0__inst_mult_11_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_57 ),
	.sharein(Xd_0__inst_mult_11_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_60 ),
	.cout(Xd_0__inst_mult_11_61 ),
	.shareout(Xd_0__inst_mult_11_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_22 (
// Equation(s):
// Xd_0__inst_mult_8_60  = SUM(( !Xd_0__inst_mult_8_10_q  $ (!Xd_0__inst_mult_8_11_q  $ (((Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_1_q )))) ) + ( Xd_0__inst_mult_8_58  ) + ( Xd_0__inst_mult_8_57  ))
// Xd_0__inst_mult_8_61  = CARRY(( !Xd_0__inst_mult_8_10_q  $ (!Xd_0__inst_mult_8_11_q  $ (((Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_1_q )))) ) + ( Xd_0__inst_mult_8_58  ) + ( Xd_0__inst_mult_8_57  ))
// Xd_0__inst_mult_8_62  = SHARE((!Xd_0__inst_mult_8_10_q  & (Xd_0__inst_mult_8_11_q  & (Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_1_q ))) # (Xd_0__inst_mult_8_10_q  & (((Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_1_q )) # (Xd_0__inst_mult_8_11_q ))))

	.dataa(!Xd_0__inst_mult_8_10_q ),
	.datab(!Xd_0__inst_mult_8_11_q ),
	.datac(!Xd_0__inst_mult_8_2_q ),
	.datad(!Xd_0__inst_mult_8_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_57 ),
	.sharein(Xd_0__inst_mult_8_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_60 ),
	.cout(Xd_0__inst_mult_8_61 ),
	.shareout(Xd_0__inst_mult_8_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_22 (
// Equation(s):
// Xd_0__inst_mult_9_60  = SUM(( !Xd_0__inst_mult_9_10_q  $ (!Xd_0__inst_mult_9_11_q  $ (((Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_1_q )))) ) + ( Xd_0__inst_mult_9_58  ) + ( Xd_0__inst_mult_9_57  ))
// Xd_0__inst_mult_9_61  = CARRY(( !Xd_0__inst_mult_9_10_q  $ (!Xd_0__inst_mult_9_11_q  $ (((Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_1_q )))) ) + ( Xd_0__inst_mult_9_58  ) + ( Xd_0__inst_mult_9_57  ))
// Xd_0__inst_mult_9_62  = SHARE((!Xd_0__inst_mult_9_10_q  & (Xd_0__inst_mult_9_11_q  & (Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_1_q ))) # (Xd_0__inst_mult_9_10_q  & (((Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_1_q )) # (Xd_0__inst_mult_9_11_q ))))

	.dataa(!Xd_0__inst_mult_9_10_q ),
	.datab(!Xd_0__inst_mult_9_11_q ),
	.datac(!Xd_0__inst_mult_9_2_q ),
	.datad(!Xd_0__inst_mult_9_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_57 ),
	.sharein(Xd_0__inst_mult_9_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_60 ),
	.cout(Xd_0__inst_mult_9_61 ),
	.shareout(Xd_0__inst_mult_9_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_22 (
// Equation(s):
// Xd_0__inst_mult_6_60  = SUM(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q  $ (((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_1_q )))) ) + ( Xd_0__inst_mult_6_58  ) + ( Xd_0__inst_mult_6_57  ))
// Xd_0__inst_mult_6_61  = CARRY(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q  $ (((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_1_q )))) ) + ( Xd_0__inst_mult_6_58  ) + ( Xd_0__inst_mult_6_57  ))
// Xd_0__inst_mult_6_62  = SHARE((!Xd_0__inst_mult_6_10_q  & (Xd_0__inst_mult_6_11_q  & (Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_1_q ))) # (Xd_0__inst_mult_6_10_q  & (((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_1_q )) # (Xd_0__inst_mult_6_11_q ))))

	.dataa(!Xd_0__inst_mult_6_10_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(!Xd_0__inst_mult_6_2_q ),
	.datad(!Xd_0__inst_mult_6_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_57 ),
	.sharein(Xd_0__inst_mult_6_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_60 ),
	.cout(Xd_0__inst_mult_6_61 ),
	.shareout(Xd_0__inst_mult_6_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_22 (
// Equation(s):
// Xd_0__inst_mult_7_60  = SUM(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q  $ (((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_1_q )))) ) + ( Xd_0__inst_mult_7_58  ) + ( Xd_0__inst_mult_7_57  ))
// Xd_0__inst_mult_7_61  = CARRY(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q  $ (((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_1_q )))) ) + ( Xd_0__inst_mult_7_58  ) + ( Xd_0__inst_mult_7_57  ))
// Xd_0__inst_mult_7_62  = SHARE((!Xd_0__inst_mult_7_10_q  & (Xd_0__inst_mult_7_11_q  & (Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_1_q ))) # (Xd_0__inst_mult_7_10_q  & (((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_1_q )) # (Xd_0__inst_mult_7_11_q ))))

	.dataa(!Xd_0__inst_mult_7_10_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(!Xd_0__inst_mult_7_2_q ),
	.datad(!Xd_0__inst_mult_7_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_57 ),
	.sharein(Xd_0__inst_mult_7_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_60 ),
	.cout(Xd_0__inst_mult_7_61 ),
	.shareout(Xd_0__inst_mult_7_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_22 (
// Equation(s):
// Xd_0__inst_mult_4_60  = SUM(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q  $ (((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_1_q )))) ) + ( Xd_0__inst_mult_4_58  ) + ( Xd_0__inst_mult_4_57  ))
// Xd_0__inst_mult_4_61  = CARRY(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q  $ (((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_1_q )))) ) + ( Xd_0__inst_mult_4_58  ) + ( Xd_0__inst_mult_4_57  ))
// Xd_0__inst_mult_4_62  = SHARE((!Xd_0__inst_mult_4_10_q  & (Xd_0__inst_mult_4_11_q  & (Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_1_q ))) # (Xd_0__inst_mult_4_10_q  & (((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_1_q )) # (Xd_0__inst_mult_4_11_q ))))

	.dataa(!Xd_0__inst_mult_4_10_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(!Xd_0__inst_mult_4_2_q ),
	.datad(!Xd_0__inst_mult_4_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_57 ),
	.sharein(Xd_0__inst_mult_4_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_60 ),
	.cout(Xd_0__inst_mult_4_61 ),
	.shareout(Xd_0__inst_mult_4_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_22 (
// Equation(s):
// Xd_0__inst_mult_5_60  = SUM(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q  $ (((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_1_q )))) ) + ( Xd_0__inst_mult_5_58  ) + ( Xd_0__inst_mult_5_57  ))
// Xd_0__inst_mult_5_61  = CARRY(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q  $ (((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_1_q )))) ) + ( Xd_0__inst_mult_5_58  ) + ( Xd_0__inst_mult_5_57  ))
// Xd_0__inst_mult_5_62  = SHARE((!Xd_0__inst_mult_5_10_q  & (Xd_0__inst_mult_5_11_q  & (Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_1_q ))) # (Xd_0__inst_mult_5_10_q  & (((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_1_q )) # (Xd_0__inst_mult_5_11_q ))))

	.dataa(!Xd_0__inst_mult_5_10_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(!Xd_0__inst_mult_5_2_q ),
	.datad(!Xd_0__inst_mult_5_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_57 ),
	.sharein(Xd_0__inst_mult_5_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_60 ),
	.cout(Xd_0__inst_mult_5_61 ),
	.shareout(Xd_0__inst_mult_5_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_22 (
// Equation(s):
// Xd_0__inst_mult_2_60  = SUM(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q  $ (((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_1_q )))) ) + ( Xd_0__inst_mult_2_58  ) + ( Xd_0__inst_mult_2_57  ))
// Xd_0__inst_mult_2_61  = CARRY(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q  $ (((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_1_q )))) ) + ( Xd_0__inst_mult_2_58  ) + ( Xd_0__inst_mult_2_57  ))
// Xd_0__inst_mult_2_62  = SHARE((!Xd_0__inst_mult_2_10_q  & (Xd_0__inst_mult_2_11_q  & (Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_1_q ))) # (Xd_0__inst_mult_2_10_q  & (((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_1_q )) # (Xd_0__inst_mult_2_11_q ))))

	.dataa(!Xd_0__inst_mult_2_10_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(!Xd_0__inst_mult_2_2_q ),
	.datad(!Xd_0__inst_mult_2_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_57 ),
	.sharein(Xd_0__inst_mult_2_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_60 ),
	.cout(Xd_0__inst_mult_2_61 ),
	.shareout(Xd_0__inst_mult_2_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_22 (
// Equation(s):
// Xd_0__inst_mult_3_60  = SUM(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q  $ (((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_1_q )))) ) + ( Xd_0__inst_mult_3_58  ) + ( Xd_0__inst_mult_3_57  ))
// Xd_0__inst_mult_3_61  = CARRY(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q  $ (((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_1_q )))) ) + ( Xd_0__inst_mult_3_58  ) + ( Xd_0__inst_mult_3_57  ))
// Xd_0__inst_mult_3_62  = SHARE((!Xd_0__inst_mult_3_10_q  & (Xd_0__inst_mult_3_11_q  & (Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_1_q ))) # (Xd_0__inst_mult_3_10_q  & (((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_1_q )) # (Xd_0__inst_mult_3_11_q ))))

	.dataa(!Xd_0__inst_mult_3_10_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(!Xd_0__inst_mult_3_2_q ),
	.datad(!Xd_0__inst_mult_3_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_57 ),
	.sharein(Xd_0__inst_mult_3_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_60 ),
	.cout(Xd_0__inst_mult_3_61 ),
	.shareout(Xd_0__inst_mult_3_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_22 (
// Equation(s):
// Xd_0__inst_mult_0_60  = SUM(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q  $ (((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_1_q )))) ) + ( Xd_0__inst_mult_0_58  ) + ( Xd_0__inst_mult_0_57  ))
// Xd_0__inst_mult_0_61  = CARRY(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q  $ (((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_1_q )))) ) + ( Xd_0__inst_mult_0_58  ) + ( Xd_0__inst_mult_0_57  ))
// Xd_0__inst_mult_0_62  = SHARE((!Xd_0__inst_mult_0_10_q  & (Xd_0__inst_mult_0_11_q  & (Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_1_q ))) # (Xd_0__inst_mult_0_10_q  & (((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_1_q )) # (Xd_0__inst_mult_0_11_q ))))

	.dataa(!Xd_0__inst_mult_0_10_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(!Xd_0__inst_mult_0_2_q ),
	.datad(!Xd_0__inst_mult_0_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_57 ),
	.sharein(Xd_0__inst_mult_0_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_60 ),
	.cout(Xd_0__inst_mult_0_61 ),
	.shareout(Xd_0__inst_mult_0_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_22 (
// Equation(s):
// Xd_0__inst_mult_1_60  = SUM(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q  $ (((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_1_q )))) ) + ( Xd_0__inst_mult_1_58  ) + ( Xd_0__inst_mult_1_57  ))
// Xd_0__inst_mult_1_61  = CARRY(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q  $ (((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_1_q )))) ) + ( Xd_0__inst_mult_1_58  ) + ( Xd_0__inst_mult_1_57  ))
// Xd_0__inst_mult_1_62  = SHARE((!Xd_0__inst_mult_1_10_q  & (Xd_0__inst_mult_1_11_q  & (Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_1_q ))) # (Xd_0__inst_mult_1_10_q  & (((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_1_q )) # (Xd_0__inst_mult_1_11_q ))))

	.dataa(!Xd_0__inst_mult_1_10_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(!Xd_0__inst_mult_1_2_q ),
	.datad(!Xd_0__inst_mult_1_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_57 ),
	.sharein(Xd_0__inst_mult_1_58 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_60 ),
	.cout(Xd_0__inst_mult_1_61 ),
	.shareout(Xd_0__inst_mult_1_62 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_28_23 (
// Equation(s):
// Xd_0__inst_mult_28_64  = SUM(( !Xd_0__inst_mult_28_12_q  $ (!Xd_0__inst_mult_28_13_q ) ) + ( Xd_0__inst_mult_28_62  ) + ( Xd_0__inst_mult_28_61  ))
// Xd_0__inst_mult_28_65  = CARRY(( !Xd_0__inst_mult_28_12_q  $ (!Xd_0__inst_mult_28_13_q ) ) + ( Xd_0__inst_mult_28_62  ) + ( Xd_0__inst_mult_28_61  ))
// Xd_0__inst_mult_28_66  = SHARE((Xd_0__inst_mult_28_12_q  & Xd_0__inst_mult_28_13_q ))

	.dataa(!Xd_0__inst_mult_28_12_q ),
	.datab(!Xd_0__inst_mult_28_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_61 ),
	.sharein(Xd_0__inst_mult_28_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_64 ),
	.cout(Xd_0__inst_mult_28_65 ),
	.shareout(Xd_0__inst_mult_28_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_29_23 (
// Equation(s):
// Xd_0__inst_mult_29_64  = SUM(( !Xd_0__inst_mult_29_12_q  $ (!Xd_0__inst_mult_29_13_q ) ) + ( Xd_0__inst_mult_29_62  ) + ( Xd_0__inst_mult_29_61  ))
// Xd_0__inst_mult_29_65  = CARRY(( !Xd_0__inst_mult_29_12_q  $ (!Xd_0__inst_mult_29_13_q ) ) + ( Xd_0__inst_mult_29_62  ) + ( Xd_0__inst_mult_29_61  ))
// Xd_0__inst_mult_29_66  = SHARE((Xd_0__inst_mult_29_12_q  & Xd_0__inst_mult_29_13_q ))

	.dataa(!Xd_0__inst_mult_29_12_q ),
	.datab(!Xd_0__inst_mult_29_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_61 ),
	.sharein(Xd_0__inst_mult_29_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_64 ),
	.cout(Xd_0__inst_mult_29_65 ),
	.shareout(Xd_0__inst_mult_29_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_26_23 (
// Equation(s):
// Xd_0__inst_mult_26_64  = SUM(( !Xd_0__inst_mult_26_12_q  $ (!Xd_0__inst_mult_26_13_q ) ) + ( Xd_0__inst_mult_26_62  ) + ( Xd_0__inst_mult_26_61  ))
// Xd_0__inst_mult_26_65  = CARRY(( !Xd_0__inst_mult_26_12_q  $ (!Xd_0__inst_mult_26_13_q ) ) + ( Xd_0__inst_mult_26_62  ) + ( Xd_0__inst_mult_26_61  ))
// Xd_0__inst_mult_26_66  = SHARE((Xd_0__inst_mult_26_12_q  & Xd_0__inst_mult_26_13_q ))

	.dataa(!Xd_0__inst_mult_26_12_q ),
	.datab(!Xd_0__inst_mult_26_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_61 ),
	.sharein(Xd_0__inst_mult_26_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_64 ),
	.cout(Xd_0__inst_mult_26_65 ),
	.shareout(Xd_0__inst_mult_26_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_27_23 (
// Equation(s):
// Xd_0__inst_mult_27_64  = SUM(( !Xd_0__inst_mult_27_12_q  $ (!Xd_0__inst_mult_27_13_q ) ) + ( Xd_0__inst_mult_27_62  ) + ( Xd_0__inst_mult_27_61  ))
// Xd_0__inst_mult_27_65  = CARRY(( !Xd_0__inst_mult_27_12_q  $ (!Xd_0__inst_mult_27_13_q ) ) + ( Xd_0__inst_mult_27_62  ) + ( Xd_0__inst_mult_27_61  ))
// Xd_0__inst_mult_27_66  = SHARE((Xd_0__inst_mult_27_12_q  & Xd_0__inst_mult_27_13_q ))

	.dataa(!Xd_0__inst_mult_27_12_q ),
	.datab(!Xd_0__inst_mult_27_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_61 ),
	.sharein(Xd_0__inst_mult_27_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_64 ),
	.cout(Xd_0__inst_mult_27_65 ),
	.shareout(Xd_0__inst_mult_27_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_24_23 (
// Equation(s):
// Xd_0__inst_mult_24_64  = SUM(( !Xd_0__inst_mult_24_12_q  $ (!Xd_0__inst_mult_24_13_q ) ) + ( Xd_0__inst_mult_24_62  ) + ( Xd_0__inst_mult_24_61  ))
// Xd_0__inst_mult_24_65  = CARRY(( !Xd_0__inst_mult_24_12_q  $ (!Xd_0__inst_mult_24_13_q ) ) + ( Xd_0__inst_mult_24_62  ) + ( Xd_0__inst_mult_24_61  ))
// Xd_0__inst_mult_24_66  = SHARE((Xd_0__inst_mult_24_12_q  & Xd_0__inst_mult_24_13_q ))

	.dataa(!Xd_0__inst_mult_24_12_q ),
	.datab(!Xd_0__inst_mult_24_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_61 ),
	.sharein(Xd_0__inst_mult_24_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_64 ),
	.cout(Xd_0__inst_mult_24_65 ),
	.shareout(Xd_0__inst_mult_24_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_25_23 (
// Equation(s):
// Xd_0__inst_mult_25_64  = SUM(( !Xd_0__inst_mult_25_12_q  $ (!Xd_0__inst_mult_25_13_q ) ) + ( Xd_0__inst_mult_25_62  ) + ( Xd_0__inst_mult_25_61  ))
// Xd_0__inst_mult_25_65  = CARRY(( !Xd_0__inst_mult_25_12_q  $ (!Xd_0__inst_mult_25_13_q ) ) + ( Xd_0__inst_mult_25_62  ) + ( Xd_0__inst_mult_25_61  ))
// Xd_0__inst_mult_25_66  = SHARE((Xd_0__inst_mult_25_12_q  & Xd_0__inst_mult_25_13_q ))

	.dataa(!Xd_0__inst_mult_25_12_q ),
	.datab(!Xd_0__inst_mult_25_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_61 ),
	.sharein(Xd_0__inst_mult_25_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_64 ),
	.cout(Xd_0__inst_mult_25_65 ),
	.shareout(Xd_0__inst_mult_25_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_22_23 (
// Equation(s):
// Xd_0__inst_mult_22_64  = SUM(( !Xd_0__inst_mult_22_12_q  $ (!Xd_0__inst_mult_22_13_q ) ) + ( Xd_0__inst_mult_22_62  ) + ( Xd_0__inst_mult_22_61  ))
// Xd_0__inst_mult_22_65  = CARRY(( !Xd_0__inst_mult_22_12_q  $ (!Xd_0__inst_mult_22_13_q ) ) + ( Xd_0__inst_mult_22_62  ) + ( Xd_0__inst_mult_22_61  ))
// Xd_0__inst_mult_22_66  = SHARE((Xd_0__inst_mult_22_12_q  & Xd_0__inst_mult_22_13_q ))

	.dataa(!Xd_0__inst_mult_22_12_q ),
	.datab(!Xd_0__inst_mult_22_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_61 ),
	.sharein(Xd_0__inst_mult_22_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_64 ),
	.cout(Xd_0__inst_mult_22_65 ),
	.shareout(Xd_0__inst_mult_22_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_23_23 (
// Equation(s):
// Xd_0__inst_mult_23_64  = SUM(( !Xd_0__inst_mult_23_12_q  $ (!Xd_0__inst_mult_23_13_q ) ) + ( Xd_0__inst_mult_23_62  ) + ( Xd_0__inst_mult_23_61  ))
// Xd_0__inst_mult_23_65  = CARRY(( !Xd_0__inst_mult_23_12_q  $ (!Xd_0__inst_mult_23_13_q ) ) + ( Xd_0__inst_mult_23_62  ) + ( Xd_0__inst_mult_23_61  ))
// Xd_0__inst_mult_23_66  = SHARE((Xd_0__inst_mult_23_12_q  & Xd_0__inst_mult_23_13_q ))

	.dataa(!Xd_0__inst_mult_23_12_q ),
	.datab(!Xd_0__inst_mult_23_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_61 ),
	.sharein(Xd_0__inst_mult_23_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_64 ),
	.cout(Xd_0__inst_mult_23_65 ),
	.shareout(Xd_0__inst_mult_23_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_20_23 (
// Equation(s):
// Xd_0__inst_mult_20_64  = SUM(( !Xd_0__inst_mult_20_12_q  $ (!Xd_0__inst_mult_20_13_q ) ) + ( Xd_0__inst_mult_20_62  ) + ( Xd_0__inst_mult_20_61  ))
// Xd_0__inst_mult_20_65  = CARRY(( !Xd_0__inst_mult_20_12_q  $ (!Xd_0__inst_mult_20_13_q ) ) + ( Xd_0__inst_mult_20_62  ) + ( Xd_0__inst_mult_20_61  ))
// Xd_0__inst_mult_20_66  = SHARE((Xd_0__inst_mult_20_12_q  & Xd_0__inst_mult_20_13_q ))

	.dataa(!Xd_0__inst_mult_20_12_q ),
	.datab(!Xd_0__inst_mult_20_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_61 ),
	.sharein(Xd_0__inst_mult_20_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_64 ),
	.cout(Xd_0__inst_mult_20_65 ),
	.shareout(Xd_0__inst_mult_20_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_21_23 (
// Equation(s):
// Xd_0__inst_mult_21_64  = SUM(( !Xd_0__inst_mult_21_12_q  $ (!Xd_0__inst_mult_21_13_q ) ) + ( Xd_0__inst_mult_21_62  ) + ( Xd_0__inst_mult_21_61  ))
// Xd_0__inst_mult_21_65  = CARRY(( !Xd_0__inst_mult_21_12_q  $ (!Xd_0__inst_mult_21_13_q ) ) + ( Xd_0__inst_mult_21_62  ) + ( Xd_0__inst_mult_21_61  ))
// Xd_0__inst_mult_21_66  = SHARE((Xd_0__inst_mult_21_12_q  & Xd_0__inst_mult_21_13_q ))

	.dataa(!Xd_0__inst_mult_21_12_q ),
	.datab(!Xd_0__inst_mult_21_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_61 ),
	.sharein(Xd_0__inst_mult_21_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_64 ),
	.cout(Xd_0__inst_mult_21_65 ),
	.shareout(Xd_0__inst_mult_21_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_18_23 (
// Equation(s):
// Xd_0__inst_mult_18_64  = SUM(( !Xd_0__inst_mult_18_12_q  $ (!Xd_0__inst_mult_18_13_q ) ) + ( Xd_0__inst_mult_18_62  ) + ( Xd_0__inst_mult_18_61  ))
// Xd_0__inst_mult_18_65  = CARRY(( !Xd_0__inst_mult_18_12_q  $ (!Xd_0__inst_mult_18_13_q ) ) + ( Xd_0__inst_mult_18_62  ) + ( Xd_0__inst_mult_18_61  ))
// Xd_0__inst_mult_18_66  = SHARE((Xd_0__inst_mult_18_12_q  & Xd_0__inst_mult_18_13_q ))

	.dataa(!Xd_0__inst_mult_18_12_q ),
	.datab(!Xd_0__inst_mult_18_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_61 ),
	.sharein(Xd_0__inst_mult_18_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_64 ),
	.cout(Xd_0__inst_mult_18_65 ),
	.shareout(Xd_0__inst_mult_18_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_19_23 (
// Equation(s):
// Xd_0__inst_mult_19_64  = SUM(( !Xd_0__inst_mult_19_12_q  $ (!Xd_0__inst_mult_19_13_q ) ) + ( Xd_0__inst_mult_19_62  ) + ( Xd_0__inst_mult_19_61  ))
// Xd_0__inst_mult_19_65  = CARRY(( !Xd_0__inst_mult_19_12_q  $ (!Xd_0__inst_mult_19_13_q ) ) + ( Xd_0__inst_mult_19_62  ) + ( Xd_0__inst_mult_19_61  ))
// Xd_0__inst_mult_19_66  = SHARE((Xd_0__inst_mult_19_12_q  & Xd_0__inst_mult_19_13_q ))

	.dataa(!Xd_0__inst_mult_19_12_q ),
	.datab(!Xd_0__inst_mult_19_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_61 ),
	.sharein(Xd_0__inst_mult_19_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_64 ),
	.cout(Xd_0__inst_mult_19_65 ),
	.shareout(Xd_0__inst_mult_19_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_16_23 (
// Equation(s):
// Xd_0__inst_mult_16_64  = SUM(( !Xd_0__inst_mult_16_12_q  $ (!Xd_0__inst_mult_16_13_q ) ) + ( Xd_0__inst_mult_16_62  ) + ( Xd_0__inst_mult_16_61  ))
// Xd_0__inst_mult_16_65  = CARRY(( !Xd_0__inst_mult_16_12_q  $ (!Xd_0__inst_mult_16_13_q ) ) + ( Xd_0__inst_mult_16_62  ) + ( Xd_0__inst_mult_16_61  ))
// Xd_0__inst_mult_16_66  = SHARE((Xd_0__inst_mult_16_12_q  & Xd_0__inst_mult_16_13_q ))

	.dataa(!Xd_0__inst_mult_16_12_q ),
	.datab(!Xd_0__inst_mult_16_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_61 ),
	.sharein(Xd_0__inst_mult_16_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_64 ),
	.cout(Xd_0__inst_mult_16_65 ),
	.shareout(Xd_0__inst_mult_16_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_17_23 (
// Equation(s):
// Xd_0__inst_mult_17_64  = SUM(( !Xd_0__inst_mult_17_12_q  $ (!Xd_0__inst_mult_17_13_q ) ) + ( Xd_0__inst_mult_17_62  ) + ( Xd_0__inst_mult_17_61  ))
// Xd_0__inst_mult_17_65  = CARRY(( !Xd_0__inst_mult_17_12_q  $ (!Xd_0__inst_mult_17_13_q ) ) + ( Xd_0__inst_mult_17_62  ) + ( Xd_0__inst_mult_17_61  ))
// Xd_0__inst_mult_17_66  = SHARE((Xd_0__inst_mult_17_12_q  & Xd_0__inst_mult_17_13_q ))

	.dataa(!Xd_0__inst_mult_17_12_q ),
	.datab(!Xd_0__inst_mult_17_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_61 ),
	.sharein(Xd_0__inst_mult_17_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_64 ),
	.cout(Xd_0__inst_mult_17_65 ),
	.shareout(Xd_0__inst_mult_17_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_23 (
// Equation(s):
// Xd_0__inst_mult_14_64  = SUM(( !Xd_0__inst_mult_14_12_q  $ (!Xd_0__inst_mult_14_13_q ) ) + ( Xd_0__inst_mult_14_62  ) + ( Xd_0__inst_mult_14_61  ))
// Xd_0__inst_mult_14_65  = CARRY(( !Xd_0__inst_mult_14_12_q  $ (!Xd_0__inst_mult_14_13_q ) ) + ( Xd_0__inst_mult_14_62  ) + ( Xd_0__inst_mult_14_61  ))
// Xd_0__inst_mult_14_66  = SHARE((Xd_0__inst_mult_14_12_q  & Xd_0__inst_mult_14_13_q ))

	.dataa(!Xd_0__inst_mult_14_12_q ),
	.datab(!Xd_0__inst_mult_14_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_61 ),
	.sharein(Xd_0__inst_mult_14_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_64 ),
	.cout(Xd_0__inst_mult_14_65 ),
	.shareout(Xd_0__inst_mult_14_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_23 (
// Equation(s):
// Xd_0__inst_mult_15_64  = SUM(( !Xd_0__inst_mult_15_12_q  $ (!Xd_0__inst_mult_15_13_q ) ) + ( Xd_0__inst_mult_15_62  ) + ( Xd_0__inst_mult_15_61  ))
// Xd_0__inst_mult_15_65  = CARRY(( !Xd_0__inst_mult_15_12_q  $ (!Xd_0__inst_mult_15_13_q ) ) + ( Xd_0__inst_mult_15_62  ) + ( Xd_0__inst_mult_15_61  ))
// Xd_0__inst_mult_15_66  = SHARE((Xd_0__inst_mult_15_12_q  & Xd_0__inst_mult_15_13_q ))

	.dataa(!Xd_0__inst_mult_15_12_q ),
	.datab(!Xd_0__inst_mult_15_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_61 ),
	.sharein(Xd_0__inst_mult_15_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_64 ),
	.cout(Xd_0__inst_mult_15_65 ),
	.shareout(Xd_0__inst_mult_15_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_23 (
// Equation(s):
// Xd_0__inst_mult_12_64  = SUM(( !Xd_0__inst_mult_12_12_q  $ (!Xd_0__inst_mult_12_13_q ) ) + ( Xd_0__inst_mult_12_62  ) + ( Xd_0__inst_mult_12_61  ))
// Xd_0__inst_mult_12_65  = CARRY(( !Xd_0__inst_mult_12_12_q  $ (!Xd_0__inst_mult_12_13_q ) ) + ( Xd_0__inst_mult_12_62  ) + ( Xd_0__inst_mult_12_61  ))
// Xd_0__inst_mult_12_66  = SHARE((Xd_0__inst_mult_12_12_q  & Xd_0__inst_mult_12_13_q ))

	.dataa(!Xd_0__inst_mult_12_12_q ),
	.datab(!Xd_0__inst_mult_12_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_61 ),
	.sharein(Xd_0__inst_mult_12_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_64 ),
	.cout(Xd_0__inst_mult_12_65 ),
	.shareout(Xd_0__inst_mult_12_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_23 (
// Equation(s):
// Xd_0__inst_mult_13_64  = SUM(( !Xd_0__inst_mult_13_12_q  $ (!Xd_0__inst_mult_13_13_q ) ) + ( Xd_0__inst_mult_13_62  ) + ( Xd_0__inst_mult_13_61  ))
// Xd_0__inst_mult_13_65  = CARRY(( !Xd_0__inst_mult_13_12_q  $ (!Xd_0__inst_mult_13_13_q ) ) + ( Xd_0__inst_mult_13_62  ) + ( Xd_0__inst_mult_13_61  ))
// Xd_0__inst_mult_13_66  = SHARE((Xd_0__inst_mult_13_12_q  & Xd_0__inst_mult_13_13_q ))

	.dataa(!Xd_0__inst_mult_13_12_q ),
	.datab(!Xd_0__inst_mult_13_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_61 ),
	.sharein(Xd_0__inst_mult_13_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_64 ),
	.cout(Xd_0__inst_mult_13_65 ),
	.shareout(Xd_0__inst_mult_13_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_23 (
// Equation(s):
// Xd_0__inst_mult_10_64  = SUM(( !Xd_0__inst_mult_10_12_q  $ (!Xd_0__inst_mult_10_13_q ) ) + ( Xd_0__inst_mult_10_62  ) + ( Xd_0__inst_mult_10_61  ))
// Xd_0__inst_mult_10_65  = CARRY(( !Xd_0__inst_mult_10_12_q  $ (!Xd_0__inst_mult_10_13_q ) ) + ( Xd_0__inst_mult_10_62  ) + ( Xd_0__inst_mult_10_61  ))
// Xd_0__inst_mult_10_66  = SHARE((Xd_0__inst_mult_10_12_q  & Xd_0__inst_mult_10_13_q ))

	.dataa(!Xd_0__inst_mult_10_12_q ),
	.datab(!Xd_0__inst_mult_10_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_61 ),
	.sharein(Xd_0__inst_mult_10_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_64 ),
	.cout(Xd_0__inst_mult_10_65 ),
	.shareout(Xd_0__inst_mult_10_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_23 (
// Equation(s):
// Xd_0__inst_mult_11_64  = SUM(( !Xd_0__inst_mult_11_12_q  $ (!Xd_0__inst_mult_11_13_q ) ) + ( Xd_0__inst_mult_11_62  ) + ( Xd_0__inst_mult_11_61  ))
// Xd_0__inst_mult_11_65  = CARRY(( !Xd_0__inst_mult_11_12_q  $ (!Xd_0__inst_mult_11_13_q ) ) + ( Xd_0__inst_mult_11_62  ) + ( Xd_0__inst_mult_11_61  ))
// Xd_0__inst_mult_11_66  = SHARE((Xd_0__inst_mult_11_12_q  & Xd_0__inst_mult_11_13_q ))

	.dataa(!Xd_0__inst_mult_11_12_q ),
	.datab(!Xd_0__inst_mult_11_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_61 ),
	.sharein(Xd_0__inst_mult_11_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_64 ),
	.cout(Xd_0__inst_mult_11_65 ),
	.shareout(Xd_0__inst_mult_11_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_23 (
// Equation(s):
// Xd_0__inst_mult_8_64  = SUM(( !Xd_0__inst_mult_8_12_q  $ (!Xd_0__inst_mult_8_13_q ) ) + ( Xd_0__inst_mult_8_62  ) + ( Xd_0__inst_mult_8_61  ))
// Xd_0__inst_mult_8_65  = CARRY(( !Xd_0__inst_mult_8_12_q  $ (!Xd_0__inst_mult_8_13_q ) ) + ( Xd_0__inst_mult_8_62  ) + ( Xd_0__inst_mult_8_61  ))
// Xd_0__inst_mult_8_66  = SHARE((Xd_0__inst_mult_8_12_q  & Xd_0__inst_mult_8_13_q ))

	.dataa(!Xd_0__inst_mult_8_12_q ),
	.datab(!Xd_0__inst_mult_8_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_61 ),
	.sharein(Xd_0__inst_mult_8_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_64 ),
	.cout(Xd_0__inst_mult_8_65 ),
	.shareout(Xd_0__inst_mult_8_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_23 (
// Equation(s):
// Xd_0__inst_mult_9_64  = SUM(( !Xd_0__inst_mult_9_12_q  $ (!Xd_0__inst_mult_9_13_q ) ) + ( Xd_0__inst_mult_9_62  ) + ( Xd_0__inst_mult_9_61  ))
// Xd_0__inst_mult_9_65  = CARRY(( !Xd_0__inst_mult_9_12_q  $ (!Xd_0__inst_mult_9_13_q ) ) + ( Xd_0__inst_mult_9_62  ) + ( Xd_0__inst_mult_9_61  ))
// Xd_0__inst_mult_9_66  = SHARE((Xd_0__inst_mult_9_12_q  & Xd_0__inst_mult_9_13_q ))

	.dataa(!Xd_0__inst_mult_9_12_q ),
	.datab(!Xd_0__inst_mult_9_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_61 ),
	.sharein(Xd_0__inst_mult_9_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_64 ),
	.cout(Xd_0__inst_mult_9_65 ),
	.shareout(Xd_0__inst_mult_9_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_23 (
// Equation(s):
// Xd_0__inst_mult_6_64  = SUM(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_62  ) + ( Xd_0__inst_mult_6_61  ))
// Xd_0__inst_mult_6_65  = CARRY(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_62  ) + ( Xd_0__inst_mult_6_61  ))
// Xd_0__inst_mult_6_66  = SHARE((Xd_0__inst_mult_6_12_q  & Xd_0__inst_mult_6_13_q ))

	.dataa(!Xd_0__inst_mult_6_12_q ),
	.datab(!Xd_0__inst_mult_6_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_61 ),
	.sharein(Xd_0__inst_mult_6_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_64 ),
	.cout(Xd_0__inst_mult_6_65 ),
	.shareout(Xd_0__inst_mult_6_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_23 (
// Equation(s):
// Xd_0__inst_mult_7_64  = SUM(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_62  ) + ( Xd_0__inst_mult_7_61  ))
// Xd_0__inst_mult_7_65  = CARRY(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_62  ) + ( Xd_0__inst_mult_7_61  ))
// Xd_0__inst_mult_7_66  = SHARE((Xd_0__inst_mult_7_12_q  & Xd_0__inst_mult_7_13_q ))

	.dataa(!Xd_0__inst_mult_7_12_q ),
	.datab(!Xd_0__inst_mult_7_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_61 ),
	.sharein(Xd_0__inst_mult_7_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_64 ),
	.cout(Xd_0__inst_mult_7_65 ),
	.shareout(Xd_0__inst_mult_7_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_23 (
// Equation(s):
// Xd_0__inst_mult_4_64  = SUM(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_62  ) + ( Xd_0__inst_mult_4_61  ))
// Xd_0__inst_mult_4_65  = CARRY(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_62  ) + ( Xd_0__inst_mult_4_61  ))
// Xd_0__inst_mult_4_66  = SHARE((Xd_0__inst_mult_4_12_q  & Xd_0__inst_mult_4_13_q ))

	.dataa(!Xd_0__inst_mult_4_12_q ),
	.datab(!Xd_0__inst_mult_4_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_61 ),
	.sharein(Xd_0__inst_mult_4_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_64 ),
	.cout(Xd_0__inst_mult_4_65 ),
	.shareout(Xd_0__inst_mult_4_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_23 (
// Equation(s):
// Xd_0__inst_mult_5_64  = SUM(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_62  ) + ( Xd_0__inst_mult_5_61  ))
// Xd_0__inst_mult_5_65  = CARRY(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_62  ) + ( Xd_0__inst_mult_5_61  ))
// Xd_0__inst_mult_5_66  = SHARE((Xd_0__inst_mult_5_12_q  & Xd_0__inst_mult_5_13_q ))

	.dataa(!Xd_0__inst_mult_5_12_q ),
	.datab(!Xd_0__inst_mult_5_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_61 ),
	.sharein(Xd_0__inst_mult_5_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_64 ),
	.cout(Xd_0__inst_mult_5_65 ),
	.shareout(Xd_0__inst_mult_5_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_23 (
// Equation(s):
// Xd_0__inst_mult_2_64  = SUM(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_62  ) + ( Xd_0__inst_mult_2_61  ))
// Xd_0__inst_mult_2_65  = CARRY(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_62  ) + ( Xd_0__inst_mult_2_61  ))
// Xd_0__inst_mult_2_66  = SHARE((Xd_0__inst_mult_2_12_q  & Xd_0__inst_mult_2_13_q ))

	.dataa(!Xd_0__inst_mult_2_12_q ),
	.datab(!Xd_0__inst_mult_2_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_61 ),
	.sharein(Xd_0__inst_mult_2_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_64 ),
	.cout(Xd_0__inst_mult_2_65 ),
	.shareout(Xd_0__inst_mult_2_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_23 (
// Equation(s):
// Xd_0__inst_mult_3_64  = SUM(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_62  ) + ( Xd_0__inst_mult_3_61  ))
// Xd_0__inst_mult_3_65  = CARRY(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_62  ) + ( Xd_0__inst_mult_3_61  ))
// Xd_0__inst_mult_3_66  = SHARE((Xd_0__inst_mult_3_12_q  & Xd_0__inst_mult_3_13_q ))

	.dataa(!Xd_0__inst_mult_3_12_q ),
	.datab(!Xd_0__inst_mult_3_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_61 ),
	.sharein(Xd_0__inst_mult_3_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_64 ),
	.cout(Xd_0__inst_mult_3_65 ),
	.shareout(Xd_0__inst_mult_3_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_23 (
// Equation(s):
// Xd_0__inst_mult_0_64  = SUM(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_62  ) + ( Xd_0__inst_mult_0_61  ))
// Xd_0__inst_mult_0_65  = CARRY(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_62  ) + ( Xd_0__inst_mult_0_61  ))
// Xd_0__inst_mult_0_66  = SHARE((Xd_0__inst_mult_0_12_q  & Xd_0__inst_mult_0_13_q ))

	.dataa(!Xd_0__inst_mult_0_12_q ),
	.datab(!Xd_0__inst_mult_0_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_61 ),
	.sharein(Xd_0__inst_mult_0_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_64 ),
	.cout(Xd_0__inst_mult_0_65 ),
	.shareout(Xd_0__inst_mult_0_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_23 (
// Equation(s):
// Xd_0__inst_mult_1_64  = SUM(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_62  ) + ( Xd_0__inst_mult_1_61  ))
// Xd_0__inst_mult_1_65  = CARRY(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_62  ) + ( Xd_0__inst_mult_1_61  ))
// Xd_0__inst_mult_1_66  = SHARE((Xd_0__inst_mult_1_12_q  & Xd_0__inst_mult_1_13_q ))

	.dataa(!Xd_0__inst_mult_1_12_q ),
	.datab(!Xd_0__inst_mult_1_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_61 ),
	.sharein(Xd_0__inst_mult_1_62 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_64 ),
	.cout(Xd_0__inst_mult_1_65 ),
	.shareout(Xd_0__inst_mult_1_66 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_28_24 (
// Equation(s):
// Xd_0__inst_mult_28_68  = SUM(( !Xd_0__inst_mult_28_14_q  $ (!Xd_0__inst_mult_28_15_q ) ) + ( Xd_0__inst_mult_28_66  ) + ( Xd_0__inst_mult_28_65  ))
// Xd_0__inst_mult_28_69  = CARRY(( !Xd_0__inst_mult_28_14_q  $ (!Xd_0__inst_mult_28_15_q ) ) + ( Xd_0__inst_mult_28_66  ) + ( Xd_0__inst_mult_28_65  ))
// Xd_0__inst_mult_28_70  = SHARE((Xd_0__inst_mult_28_14_q  & Xd_0__inst_mult_28_15_q ))

	.dataa(!Xd_0__inst_mult_28_14_q ),
	.datab(!Xd_0__inst_mult_28_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_65 ),
	.sharein(Xd_0__inst_mult_28_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_68 ),
	.cout(Xd_0__inst_mult_28_69 ),
	.shareout(Xd_0__inst_mult_28_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_29_24 (
// Equation(s):
// Xd_0__inst_mult_29_68  = SUM(( !Xd_0__inst_mult_29_14_q  $ (!Xd_0__inst_mult_29_15_q ) ) + ( Xd_0__inst_mult_29_66  ) + ( Xd_0__inst_mult_29_65  ))
// Xd_0__inst_mult_29_69  = CARRY(( !Xd_0__inst_mult_29_14_q  $ (!Xd_0__inst_mult_29_15_q ) ) + ( Xd_0__inst_mult_29_66  ) + ( Xd_0__inst_mult_29_65  ))
// Xd_0__inst_mult_29_70  = SHARE((Xd_0__inst_mult_29_14_q  & Xd_0__inst_mult_29_15_q ))

	.dataa(!Xd_0__inst_mult_29_14_q ),
	.datab(!Xd_0__inst_mult_29_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_65 ),
	.sharein(Xd_0__inst_mult_29_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_68 ),
	.cout(Xd_0__inst_mult_29_69 ),
	.shareout(Xd_0__inst_mult_29_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_26_24 (
// Equation(s):
// Xd_0__inst_mult_26_68  = SUM(( !Xd_0__inst_mult_26_14_q  $ (!Xd_0__inst_mult_26_15_q ) ) + ( Xd_0__inst_mult_26_66  ) + ( Xd_0__inst_mult_26_65  ))
// Xd_0__inst_mult_26_69  = CARRY(( !Xd_0__inst_mult_26_14_q  $ (!Xd_0__inst_mult_26_15_q ) ) + ( Xd_0__inst_mult_26_66  ) + ( Xd_0__inst_mult_26_65  ))
// Xd_0__inst_mult_26_70  = SHARE((Xd_0__inst_mult_26_14_q  & Xd_0__inst_mult_26_15_q ))

	.dataa(!Xd_0__inst_mult_26_14_q ),
	.datab(!Xd_0__inst_mult_26_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_65 ),
	.sharein(Xd_0__inst_mult_26_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_68 ),
	.cout(Xd_0__inst_mult_26_69 ),
	.shareout(Xd_0__inst_mult_26_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_27_24 (
// Equation(s):
// Xd_0__inst_mult_27_68  = SUM(( !Xd_0__inst_mult_27_14_q  $ (!Xd_0__inst_mult_27_15_q ) ) + ( Xd_0__inst_mult_27_66  ) + ( Xd_0__inst_mult_27_65  ))
// Xd_0__inst_mult_27_69  = CARRY(( !Xd_0__inst_mult_27_14_q  $ (!Xd_0__inst_mult_27_15_q ) ) + ( Xd_0__inst_mult_27_66  ) + ( Xd_0__inst_mult_27_65  ))
// Xd_0__inst_mult_27_70  = SHARE((Xd_0__inst_mult_27_14_q  & Xd_0__inst_mult_27_15_q ))

	.dataa(!Xd_0__inst_mult_27_14_q ),
	.datab(!Xd_0__inst_mult_27_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_65 ),
	.sharein(Xd_0__inst_mult_27_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_68 ),
	.cout(Xd_0__inst_mult_27_69 ),
	.shareout(Xd_0__inst_mult_27_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_24_24 (
// Equation(s):
// Xd_0__inst_mult_24_68  = SUM(( !Xd_0__inst_mult_24_14_q  $ (!Xd_0__inst_mult_24_15_q ) ) + ( Xd_0__inst_mult_24_66  ) + ( Xd_0__inst_mult_24_65  ))
// Xd_0__inst_mult_24_69  = CARRY(( !Xd_0__inst_mult_24_14_q  $ (!Xd_0__inst_mult_24_15_q ) ) + ( Xd_0__inst_mult_24_66  ) + ( Xd_0__inst_mult_24_65  ))
// Xd_0__inst_mult_24_70  = SHARE((Xd_0__inst_mult_24_14_q  & Xd_0__inst_mult_24_15_q ))

	.dataa(!Xd_0__inst_mult_24_14_q ),
	.datab(!Xd_0__inst_mult_24_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_65 ),
	.sharein(Xd_0__inst_mult_24_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_68 ),
	.cout(Xd_0__inst_mult_24_69 ),
	.shareout(Xd_0__inst_mult_24_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_25_24 (
// Equation(s):
// Xd_0__inst_mult_25_68  = SUM(( !Xd_0__inst_mult_25_14_q  $ (!Xd_0__inst_mult_25_15_q ) ) + ( Xd_0__inst_mult_25_66  ) + ( Xd_0__inst_mult_25_65  ))
// Xd_0__inst_mult_25_69  = CARRY(( !Xd_0__inst_mult_25_14_q  $ (!Xd_0__inst_mult_25_15_q ) ) + ( Xd_0__inst_mult_25_66  ) + ( Xd_0__inst_mult_25_65  ))
// Xd_0__inst_mult_25_70  = SHARE((Xd_0__inst_mult_25_14_q  & Xd_0__inst_mult_25_15_q ))

	.dataa(!Xd_0__inst_mult_25_14_q ),
	.datab(!Xd_0__inst_mult_25_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_65 ),
	.sharein(Xd_0__inst_mult_25_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_68 ),
	.cout(Xd_0__inst_mult_25_69 ),
	.shareout(Xd_0__inst_mult_25_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_22_24 (
// Equation(s):
// Xd_0__inst_mult_22_68  = SUM(( !Xd_0__inst_mult_22_14_q  $ (!Xd_0__inst_mult_22_15_q ) ) + ( Xd_0__inst_mult_22_66  ) + ( Xd_0__inst_mult_22_65  ))
// Xd_0__inst_mult_22_69  = CARRY(( !Xd_0__inst_mult_22_14_q  $ (!Xd_0__inst_mult_22_15_q ) ) + ( Xd_0__inst_mult_22_66  ) + ( Xd_0__inst_mult_22_65  ))
// Xd_0__inst_mult_22_70  = SHARE((Xd_0__inst_mult_22_14_q  & Xd_0__inst_mult_22_15_q ))

	.dataa(!Xd_0__inst_mult_22_14_q ),
	.datab(!Xd_0__inst_mult_22_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_65 ),
	.sharein(Xd_0__inst_mult_22_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_68 ),
	.cout(Xd_0__inst_mult_22_69 ),
	.shareout(Xd_0__inst_mult_22_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_23_24 (
// Equation(s):
// Xd_0__inst_mult_23_68  = SUM(( !Xd_0__inst_mult_23_14_q  $ (!Xd_0__inst_mult_23_15_q ) ) + ( Xd_0__inst_mult_23_66  ) + ( Xd_0__inst_mult_23_65  ))
// Xd_0__inst_mult_23_69  = CARRY(( !Xd_0__inst_mult_23_14_q  $ (!Xd_0__inst_mult_23_15_q ) ) + ( Xd_0__inst_mult_23_66  ) + ( Xd_0__inst_mult_23_65  ))
// Xd_0__inst_mult_23_70  = SHARE((Xd_0__inst_mult_23_14_q  & Xd_0__inst_mult_23_15_q ))

	.dataa(!Xd_0__inst_mult_23_14_q ),
	.datab(!Xd_0__inst_mult_23_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_65 ),
	.sharein(Xd_0__inst_mult_23_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_68 ),
	.cout(Xd_0__inst_mult_23_69 ),
	.shareout(Xd_0__inst_mult_23_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_20_24 (
// Equation(s):
// Xd_0__inst_mult_20_68  = SUM(( !Xd_0__inst_mult_20_14_q  $ (!Xd_0__inst_mult_20_15_q ) ) + ( Xd_0__inst_mult_20_66  ) + ( Xd_0__inst_mult_20_65  ))
// Xd_0__inst_mult_20_69  = CARRY(( !Xd_0__inst_mult_20_14_q  $ (!Xd_0__inst_mult_20_15_q ) ) + ( Xd_0__inst_mult_20_66  ) + ( Xd_0__inst_mult_20_65  ))
// Xd_0__inst_mult_20_70  = SHARE((Xd_0__inst_mult_20_14_q  & Xd_0__inst_mult_20_15_q ))

	.dataa(!Xd_0__inst_mult_20_14_q ),
	.datab(!Xd_0__inst_mult_20_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_65 ),
	.sharein(Xd_0__inst_mult_20_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_68 ),
	.cout(Xd_0__inst_mult_20_69 ),
	.shareout(Xd_0__inst_mult_20_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_21_24 (
// Equation(s):
// Xd_0__inst_mult_21_68  = SUM(( !Xd_0__inst_mult_21_14_q  $ (!Xd_0__inst_mult_21_15_q ) ) + ( Xd_0__inst_mult_21_66  ) + ( Xd_0__inst_mult_21_65  ))
// Xd_0__inst_mult_21_69  = CARRY(( !Xd_0__inst_mult_21_14_q  $ (!Xd_0__inst_mult_21_15_q ) ) + ( Xd_0__inst_mult_21_66  ) + ( Xd_0__inst_mult_21_65  ))
// Xd_0__inst_mult_21_70  = SHARE((Xd_0__inst_mult_21_14_q  & Xd_0__inst_mult_21_15_q ))

	.dataa(!Xd_0__inst_mult_21_14_q ),
	.datab(!Xd_0__inst_mult_21_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_65 ),
	.sharein(Xd_0__inst_mult_21_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_68 ),
	.cout(Xd_0__inst_mult_21_69 ),
	.shareout(Xd_0__inst_mult_21_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_18_24 (
// Equation(s):
// Xd_0__inst_mult_18_68  = SUM(( !Xd_0__inst_mult_18_14_q  $ (!Xd_0__inst_mult_18_15_q ) ) + ( Xd_0__inst_mult_18_66  ) + ( Xd_0__inst_mult_18_65  ))
// Xd_0__inst_mult_18_69  = CARRY(( !Xd_0__inst_mult_18_14_q  $ (!Xd_0__inst_mult_18_15_q ) ) + ( Xd_0__inst_mult_18_66  ) + ( Xd_0__inst_mult_18_65  ))
// Xd_0__inst_mult_18_70  = SHARE((Xd_0__inst_mult_18_14_q  & Xd_0__inst_mult_18_15_q ))

	.dataa(!Xd_0__inst_mult_18_14_q ),
	.datab(!Xd_0__inst_mult_18_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_65 ),
	.sharein(Xd_0__inst_mult_18_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_68 ),
	.cout(Xd_0__inst_mult_18_69 ),
	.shareout(Xd_0__inst_mult_18_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_19_24 (
// Equation(s):
// Xd_0__inst_mult_19_68  = SUM(( !Xd_0__inst_mult_19_14_q  $ (!Xd_0__inst_mult_19_15_q ) ) + ( Xd_0__inst_mult_19_66  ) + ( Xd_0__inst_mult_19_65  ))
// Xd_0__inst_mult_19_69  = CARRY(( !Xd_0__inst_mult_19_14_q  $ (!Xd_0__inst_mult_19_15_q ) ) + ( Xd_0__inst_mult_19_66  ) + ( Xd_0__inst_mult_19_65  ))
// Xd_0__inst_mult_19_70  = SHARE((Xd_0__inst_mult_19_14_q  & Xd_0__inst_mult_19_15_q ))

	.dataa(!Xd_0__inst_mult_19_14_q ),
	.datab(!Xd_0__inst_mult_19_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_65 ),
	.sharein(Xd_0__inst_mult_19_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_68 ),
	.cout(Xd_0__inst_mult_19_69 ),
	.shareout(Xd_0__inst_mult_19_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_16_24 (
// Equation(s):
// Xd_0__inst_mult_16_68  = SUM(( !Xd_0__inst_mult_16_14_q  $ (!Xd_0__inst_mult_16_15_q ) ) + ( Xd_0__inst_mult_16_66  ) + ( Xd_0__inst_mult_16_65  ))
// Xd_0__inst_mult_16_69  = CARRY(( !Xd_0__inst_mult_16_14_q  $ (!Xd_0__inst_mult_16_15_q ) ) + ( Xd_0__inst_mult_16_66  ) + ( Xd_0__inst_mult_16_65  ))
// Xd_0__inst_mult_16_70  = SHARE((Xd_0__inst_mult_16_14_q  & Xd_0__inst_mult_16_15_q ))

	.dataa(!Xd_0__inst_mult_16_14_q ),
	.datab(!Xd_0__inst_mult_16_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_65 ),
	.sharein(Xd_0__inst_mult_16_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_68 ),
	.cout(Xd_0__inst_mult_16_69 ),
	.shareout(Xd_0__inst_mult_16_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_17_24 (
// Equation(s):
// Xd_0__inst_mult_17_68  = SUM(( !Xd_0__inst_mult_17_14_q  $ (!Xd_0__inst_mult_17_15_q ) ) + ( Xd_0__inst_mult_17_66  ) + ( Xd_0__inst_mult_17_65  ))
// Xd_0__inst_mult_17_69  = CARRY(( !Xd_0__inst_mult_17_14_q  $ (!Xd_0__inst_mult_17_15_q ) ) + ( Xd_0__inst_mult_17_66  ) + ( Xd_0__inst_mult_17_65  ))
// Xd_0__inst_mult_17_70  = SHARE((Xd_0__inst_mult_17_14_q  & Xd_0__inst_mult_17_15_q ))

	.dataa(!Xd_0__inst_mult_17_14_q ),
	.datab(!Xd_0__inst_mult_17_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_65 ),
	.sharein(Xd_0__inst_mult_17_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_68 ),
	.cout(Xd_0__inst_mult_17_69 ),
	.shareout(Xd_0__inst_mult_17_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14_24 (
// Equation(s):
// Xd_0__inst_mult_14_68  = SUM(( !Xd_0__inst_mult_14_14_q  $ (!Xd_0__inst_mult_14_15_q ) ) + ( Xd_0__inst_mult_14_66  ) + ( Xd_0__inst_mult_14_65  ))
// Xd_0__inst_mult_14_69  = CARRY(( !Xd_0__inst_mult_14_14_q  $ (!Xd_0__inst_mult_14_15_q ) ) + ( Xd_0__inst_mult_14_66  ) + ( Xd_0__inst_mult_14_65  ))
// Xd_0__inst_mult_14_70  = SHARE((Xd_0__inst_mult_14_14_q  & Xd_0__inst_mult_14_15_q ))

	.dataa(!Xd_0__inst_mult_14_14_q ),
	.datab(!Xd_0__inst_mult_14_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_65 ),
	.sharein(Xd_0__inst_mult_14_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_68 ),
	.cout(Xd_0__inst_mult_14_69 ),
	.shareout(Xd_0__inst_mult_14_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15_24 (
// Equation(s):
// Xd_0__inst_mult_15_68  = SUM(( !Xd_0__inst_mult_15_14_q  $ (!Xd_0__inst_mult_15_15_q ) ) + ( Xd_0__inst_mult_15_66  ) + ( Xd_0__inst_mult_15_65  ))
// Xd_0__inst_mult_15_69  = CARRY(( !Xd_0__inst_mult_15_14_q  $ (!Xd_0__inst_mult_15_15_q ) ) + ( Xd_0__inst_mult_15_66  ) + ( Xd_0__inst_mult_15_65  ))
// Xd_0__inst_mult_15_70  = SHARE((Xd_0__inst_mult_15_14_q  & Xd_0__inst_mult_15_15_q ))

	.dataa(!Xd_0__inst_mult_15_14_q ),
	.datab(!Xd_0__inst_mult_15_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_65 ),
	.sharein(Xd_0__inst_mult_15_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_68 ),
	.cout(Xd_0__inst_mult_15_69 ),
	.shareout(Xd_0__inst_mult_15_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12_24 (
// Equation(s):
// Xd_0__inst_mult_12_68  = SUM(( !Xd_0__inst_mult_12_14_q  $ (!Xd_0__inst_mult_12_15_q ) ) + ( Xd_0__inst_mult_12_66  ) + ( Xd_0__inst_mult_12_65  ))
// Xd_0__inst_mult_12_69  = CARRY(( !Xd_0__inst_mult_12_14_q  $ (!Xd_0__inst_mult_12_15_q ) ) + ( Xd_0__inst_mult_12_66  ) + ( Xd_0__inst_mult_12_65  ))
// Xd_0__inst_mult_12_70  = SHARE((Xd_0__inst_mult_12_14_q  & Xd_0__inst_mult_12_15_q ))

	.dataa(!Xd_0__inst_mult_12_14_q ),
	.datab(!Xd_0__inst_mult_12_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_65 ),
	.sharein(Xd_0__inst_mult_12_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_68 ),
	.cout(Xd_0__inst_mult_12_69 ),
	.shareout(Xd_0__inst_mult_12_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13_24 (
// Equation(s):
// Xd_0__inst_mult_13_68  = SUM(( !Xd_0__inst_mult_13_14_q  $ (!Xd_0__inst_mult_13_15_q ) ) + ( Xd_0__inst_mult_13_66  ) + ( Xd_0__inst_mult_13_65  ))
// Xd_0__inst_mult_13_69  = CARRY(( !Xd_0__inst_mult_13_14_q  $ (!Xd_0__inst_mult_13_15_q ) ) + ( Xd_0__inst_mult_13_66  ) + ( Xd_0__inst_mult_13_65  ))
// Xd_0__inst_mult_13_70  = SHARE((Xd_0__inst_mult_13_14_q  & Xd_0__inst_mult_13_15_q ))

	.dataa(!Xd_0__inst_mult_13_14_q ),
	.datab(!Xd_0__inst_mult_13_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_65 ),
	.sharein(Xd_0__inst_mult_13_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_68 ),
	.cout(Xd_0__inst_mult_13_69 ),
	.shareout(Xd_0__inst_mult_13_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10_24 (
// Equation(s):
// Xd_0__inst_mult_10_68  = SUM(( !Xd_0__inst_mult_10_14_q  $ (!Xd_0__inst_mult_10_15_q ) ) + ( Xd_0__inst_mult_10_66  ) + ( Xd_0__inst_mult_10_65  ))
// Xd_0__inst_mult_10_69  = CARRY(( !Xd_0__inst_mult_10_14_q  $ (!Xd_0__inst_mult_10_15_q ) ) + ( Xd_0__inst_mult_10_66  ) + ( Xd_0__inst_mult_10_65  ))
// Xd_0__inst_mult_10_70  = SHARE((Xd_0__inst_mult_10_14_q  & Xd_0__inst_mult_10_15_q ))

	.dataa(!Xd_0__inst_mult_10_14_q ),
	.datab(!Xd_0__inst_mult_10_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_65 ),
	.sharein(Xd_0__inst_mult_10_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_68 ),
	.cout(Xd_0__inst_mult_10_69 ),
	.shareout(Xd_0__inst_mult_10_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_24 (
// Equation(s):
// Xd_0__inst_mult_11_68  = SUM(( !Xd_0__inst_mult_11_14_q  $ (!Xd_0__inst_mult_11_15_q ) ) + ( Xd_0__inst_mult_11_66  ) + ( Xd_0__inst_mult_11_65  ))
// Xd_0__inst_mult_11_69  = CARRY(( !Xd_0__inst_mult_11_14_q  $ (!Xd_0__inst_mult_11_15_q ) ) + ( Xd_0__inst_mult_11_66  ) + ( Xd_0__inst_mult_11_65  ))
// Xd_0__inst_mult_11_70  = SHARE((Xd_0__inst_mult_11_14_q  & Xd_0__inst_mult_11_15_q ))

	.dataa(!Xd_0__inst_mult_11_14_q ),
	.datab(!Xd_0__inst_mult_11_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_65 ),
	.sharein(Xd_0__inst_mult_11_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_68 ),
	.cout(Xd_0__inst_mult_11_69 ),
	.shareout(Xd_0__inst_mult_11_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8_24 (
// Equation(s):
// Xd_0__inst_mult_8_68  = SUM(( !Xd_0__inst_mult_8_14_q  $ (!Xd_0__inst_mult_8_15_q ) ) + ( Xd_0__inst_mult_8_66  ) + ( Xd_0__inst_mult_8_65  ))
// Xd_0__inst_mult_8_69  = CARRY(( !Xd_0__inst_mult_8_14_q  $ (!Xd_0__inst_mult_8_15_q ) ) + ( Xd_0__inst_mult_8_66  ) + ( Xd_0__inst_mult_8_65  ))
// Xd_0__inst_mult_8_70  = SHARE((Xd_0__inst_mult_8_14_q  & Xd_0__inst_mult_8_15_q ))

	.dataa(!Xd_0__inst_mult_8_14_q ),
	.datab(!Xd_0__inst_mult_8_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_65 ),
	.sharein(Xd_0__inst_mult_8_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_68 ),
	.cout(Xd_0__inst_mult_8_69 ),
	.shareout(Xd_0__inst_mult_8_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9_24 (
// Equation(s):
// Xd_0__inst_mult_9_68  = SUM(( !Xd_0__inst_mult_9_14_q  $ (!Xd_0__inst_mult_9_15_q ) ) + ( Xd_0__inst_mult_9_66  ) + ( Xd_0__inst_mult_9_65  ))
// Xd_0__inst_mult_9_69  = CARRY(( !Xd_0__inst_mult_9_14_q  $ (!Xd_0__inst_mult_9_15_q ) ) + ( Xd_0__inst_mult_9_66  ) + ( Xd_0__inst_mult_9_65  ))
// Xd_0__inst_mult_9_70  = SHARE((Xd_0__inst_mult_9_14_q  & Xd_0__inst_mult_9_15_q ))

	.dataa(!Xd_0__inst_mult_9_14_q ),
	.datab(!Xd_0__inst_mult_9_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_65 ),
	.sharein(Xd_0__inst_mult_9_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_68 ),
	.cout(Xd_0__inst_mult_9_69 ),
	.shareout(Xd_0__inst_mult_9_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_24 (
// Equation(s):
// Xd_0__inst_mult_6_68  = SUM(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_66  ) + ( Xd_0__inst_mult_6_65  ))
// Xd_0__inst_mult_6_69  = CARRY(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_66  ) + ( Xd_0__inst_mult_6_65  ))
// Xd_0__inst_mult_6_70  = SHARE((Xd_0__inst_mult_6_14_q  & Xd_0__inst_mult_6_15_q ))

	.dataa(!Xd_0__inst_mult_6_14_q ),
	.datab(!Xd_0__inst_mult_6_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_65 ),
	.sharein(Xd_0__inst_mult_6_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_68 ),
	.cout(Xd_0__inst_mult_6_69 ),
	.shareout(Xd_0__inst_mult_6_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_24 (
// Equation(s):
// Xd_0__inst_mult_7_68  = SUM(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_66  ) + ( Xd_0__inst_mult_7_65  ))
// Xd_0__inst_mult_7_69  = CARRY(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_66  ) + ( Xd_0__inst_mult_7_65  ))
// Xd_0__inst_mult_7_70  = SHARE((Xd_0__inst_mult_7_14_q  & Xd_0__inst_mult_7_15_q ))

	.dataa(!Xd_0__inst_mult_7_14_q ),
	.datab(!Xd_0__inst_mult_7_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_65 ),
	.sharein(Xd_0__inst_mult_7_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_68 ),
	.cout(Xd_0__inst_mult_7_69 ),
	.shareout(Xd_0__inst_mult_7_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_24 (
// Equation(s):
// Xd_0__inst_mult_4_68  = SUM(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_66  ) + ( Xd_0__inst_mult_4_65  ))
// Xd_0__inst_mult_4_69  = CARRY(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_66  ) + ( Xd_0__inst_mult_4_65  ))
// Xd_0__inst_mult_4_70  = SHARE((Xd_0__inst_mult_4_14_q  & Xd_0__inst_mult_4_15_q ))

	.dataa(!Xd_0__inst_mult_4_14_q ),
	.datab(!Xd_0__inst_mult_4_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_65 ),
	.sharein(Xd_0__inst_mult_4_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_68 ),
	.cout(Xd_0__inst_mult_4_69 ),
	.shareout(Xd_0__inst_mult_4_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_24 (
// Equation(s):
// Xd_0__inst_mult_5_68  = SUM(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_66  ) + ( Xd_0__inst_mult_5_65  ))
// Xd_0__inst_mult_5_69  = CARRY(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_66  ) + ( Xd_0__inst_mult_5_65  ))
// Xd_0__inst_mult_5_70  = SHARE((Xd_0__inst_mult_5_14_q  & Xd_0__inst_mult_5_15_q ))

	.dataa(!Xd_0__inst_mult_5_14_q ),
	.datab(!Xd_0__inst_mult_5_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_65 ),
	.sharein(Xd_0__inst_mult_5_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_68 ),
	.cout(Xd_0__inst_mult_5_69 ),
	.shareout(Xd_0__inst_mult_5_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_24 (
// Equation(s):
// Xd_0__inst_mult_2_68  = SUM(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_66  ) + ( Xd_0__inst_mult_2_65  ))
// Xd_0__inst_mult_2_69  = CARRY(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_66  ) + ( Xd_0__inst_mult_2_65  ))
// Xd_0__inst_mult_2_70  = SHARE((Xd_0__inst_mult_2_14_q  & Xd_0__inst_mult_2_15_q ))

	.dataa(!Xd_0__inst_mult_2_14_q ),
	.datab(!Xd_0__inst_mult_2_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_65 ),
	.sharein(Xd_0__inst_mult_2_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_68 ),
	.cout(Xd_0__inst_mult_2_69 ),
	.shareout(Xd_0__inst_mult_2_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_24 (
// Equation(s):
// Xd_0__inst_mult_3_68  = SUM(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_66  ) + ( Xd_0__inst_mult_3_65  ))
// Xd_0__inst_mult_3_69  = CARRY(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_66  ) + ( Xd_0__inst_mult_3_65  ))
// Xd_0__inst_mult_3_70  = SHARE((Xd_0__inst_mult_3_14_q  & Xd_0__inst_mult_3_15_q ))

	.dataa(!Xd_0__inst_mult_3_14_q ),
	.datab(!Xd_0__inst_mult_3_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_65 ),
	.sharein(Xd_0__inst_mult_3_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_68 ),
	.cout(Xd_0__inst_mult_3_69 ),
	.shareout(Xd_0__inst_mult_3_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_24 (
// Equation(s):
// Xd_0__inst_mult_0_68  = SUM(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_66  ) + ( Xd_0__inst_mult_0_65  ))
// Xd_0__inst_mult_0_69  = CARRY(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_66  ) + ( Xd_0__inst_mult_0_65  ))
// Xd_0__inst_mult_0_70  = SHARE((Xd_0__inst_mult_0_14_q  & Xd_0__inst_mult_0_15_q ))

	.dataa(!Xd_0__inst_mult_0_14_q ),
	.datab(!Xd_0__inst_mult_0_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_65 ),
	.sharein(Xd_0__inst_mult_0_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_68 ),
	.cout(Xd_0__inst_mult_0_69 ),
	.shareout(Xd_0__inst_mult_0_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_24 (
// Equation(s):
// Xd_0__inst_mult_1_68  = SUM(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_66  ) + ( Xd_0__inst_mult_1_65  ))
// Xd_0__inst_mult_1_69  = CARRY(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_66  ) + ( Xd_0__inst_mult_1_65  ))
// Xd_0__inst_mult_1_70  = SHARE((Xd_0__inst_mult_1_14_q  & Xd_0__inst_mult_1_15_q ))

	.dataa(!Xd_0__inst_mult_1_14_q ),
	.datab(!Xd_0__inst_mult_1_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_65 ),
	.sharein(Xd_0__inst_mult_1_66 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_68 ),
	.cout(Xd_0__inst_mult_1_69 ),
	.shareout(Xd_0__inst_mult_1_70 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_28_25 (
// Equation(s):
// Xd_0__inst_mult_28_72  = SUM(( !Xd_0__inst_mult_28_16_q  $ (!Xd_0__inst_mult_28_17_q  $ (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_18_q )))) ) + ( Xd_0__inst_mult_28_70  ) + ( Xd_0__inst_mult_28_69  ))
// Xd_0__inst_mult_28_73  = CARRY(( !Xd_0__inst_mult_28_16_q  $ (!Xd_0__inst_mult_28_17_q  $ (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_18_q )))) ) + ( Xd_0__inst_mult_28_70  ) + ( Xd_0__inst_mult_28_69  ))
// Xd_0__inst_mult_28_74  = SHARE((!Xd_0__inst_mult_28_16_q  & (Xd_0__inst_mult_28_17_q  & (Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_18_q ))) # (Xd_0__inst_mult_28_16_q  & (((Xd_0__inst_mult_28_7_q  & Xd_0__inst_mult_28_18_q )) # (Xd_0__inst_mult_28_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_28_16_q ),
	.datab(!Xd_0__inst_mult_28_17_q ),
	.datac(!Xd_0__inst_mult_28_7_q ),
	.datad(!Xd_0__inst_mult_28_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_69 ),
	.sharein(Xd_0__inst_mult_28_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_72 ),
	.cout(Xd_0__inst_mult_28_73 ),
	.shareout(Xd_0__inst_mult_28_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_29_25 (
// Equation(s):
// Xd_0__inst_mult_29_72  = SUM(( !Xd_0__inst_mult_29_16_q  $ (!Xd_0__inst_mult_29_17_q  $ (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_18_q )))) ) + ( Xd_0__inst_mult_29_70  ) + ( Xd_0__inst_mult_29_69  ))
// Xd_0__inst_mult_29_73  = CARRY(( !Xd_0__inst_mult_29_16_q  $ (!Xd_0__inst_mult_29_17_q  $ (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_18_q )))) ) + ( Xd_0__inst_mult_29_70  ) + ( Xd_0__inst_mult_29_69  ))
// Xd_0__inst_mult_29_74  = SHARE((!Xd_0__inst_mult_29_16_q  & (Xd_0__inst_mult_29_17_q  & (Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_18_q ))) # (Xd_0__inst_mult_29_16_q  & (((Xd_0__inst_mult_29_7_q  & Xd_0__inst_mult_29_18_q )) # (Xd_0__inst_mult_29_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_29_16_q ),
	.datab(!Xd_0__inst_mult_29_17_q ),
	.datac(!Xd_0__inst_mult_29_7_q ),
	.datad(!Xd_0__inst_mult_29_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_69 ),
	.sharein(Xd_0__inst_mult_29_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_72 ),
	.cout(Xd_0__inst_mult_29_73 ),
	.shareout(Xd_0__inst_mult_29_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_26_25 (
// Equation(s):
// Xd_0__inst_mult_26_72  = SUM(( !Xd_0__inst_mult_26_16_q  $ (!Xd_0__inst_mult_26_17_q  $ (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_18_q )))) ) + ( Xd_0__inst_mult_26_70  ) + ( Xd_0__inst_mult_26_69  ))
// Xd_0__inst_mult_26_73  = CARRY(( !Xd_0__inst_mult_26_16_q  $ (!Xd_0__inst_mult_26_17_q  $ (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_18_q )))) ) + ( Xd_0__inst_mult_26_70  ) + ( Xd_0__inst_mult_26_69  ))
// Xd_0__inst_mult_26_74  = SHARE((!Xd_0__inst_mult_26_16_q  & (Xd_0__inst_mult_26_17_q  & (Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_18_q ))) # (Xd_0__inst_mult_26_16_q  & (((Xd_0__inst_mult_26_7_q  & Xd_0__inst_mult_26_18_q )) # (Xd_0__inst_mult_26_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_26_16_q ),
	.datab(!Xd_0__inst_mult_26_17_q ),
	.datac(!Xd_0__inst_mult_26_7_q ),
	.datad(!Xd_0__inst_mult_26_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_69 ),
	.sharein(Xd_0__inst_mult_26_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_72 ),
	.cout(Xd_0__inst_mult_26_73 ),
	.shareout(Xd_0__inst_mult_26_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_27_25 (
// Equation(s):
// Xd_0__inst_mult_27_72  = SUM(( !Xd_0__inst_mult_27_16_q  $ (!Xd_0__inst_mult_27_17_q  $ (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_18_q )))) ) + ( Xd_0__inst_mult_27_70  ) + ( Xd_0__inst_mult_27_69  ))
// Xd_0__inst_mult_27_73  = CARRY(( !Xd_0__inst_mult_27_16_q  $ (!Xd_0__inst_mult_27_17_q  $ (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_18_q )))) ) + ( Xd_0__inst_mult_27_70  ) + ( Xd_0__inst_mult_27_69  ))
// Xd_0__inst_mult_27_74  = SHARE((!Xd_0__inst_mult_27_16_q  & (Xd_0__inst_mult_27_17_q  & (Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_18_q ))) # (Xd_0__inst_mult_27_16_q  & (((Xd_0__inst_mult_27_7_q  & Xd_0__inst_mult_27_18_q )) # (Xd_0__inst_mult_27_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_27_16_q ),
	.datab(!Xd_0__inst_mult_27_17_q ),
	.datac(!Xd_0__inst_mult_27_7_q ),
	.datad(!Xd_0__inst_mult_27_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_69 ),
	.sharein(Xd_0__inst_mult_27_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_72 ),
	.cout(Xd_0__inst_mult_27_73 ),
	.shareout(Xd_0__inst_mult_27_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_24_25 (
// Equation(s):
// Xd_0__inst_mult_24_72  = SUM(( !Xd_0__inst_mult_24_16_q  $ (!Xd_0__inst_mult_24_17_q  $ (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_18_q )))) ) + ( Xd_0__inst_mult_24_70  ) + ( Xd_0__inst_mult_24_69  ))
// Xd_0__inst_mult_24_73  = CARRY(( !Xd_0__inst_mult_24_16_q  $ (!Xd_0__inst_mult_24_17_q  $ (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_18_q )))) ) + ( Xd_0__inst_mult_24_70  ) + ( Xd_0__inst_mult_24_69  ))
// Xd_0__inst_mult_24_74  = SHARE((!Xd_0__inst_mult_24_16_q  & (Xd_0__inst_mult_24_17_q  & (Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_18_q ))) # (Xd_0__inst_mult_24_16_q  & (((Xd_0__inst_mult_24_7_q  & Xd_0__inst_mult_24_18_q )) # (Xd_0__inst_mult_24_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_24_16_q ),
	.datab(!Xd_0__inst_mult_24_17_q ),
	.datac(!Xd_0__inst_mult_24_7_q ),
	.datad(!Xd_0__inst_mult_24_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_69 ),
	.sharein(Xd_0__inst_mult_24_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_72 ),
	.cout(Xd_0__inst_mult_24_73 ),
	.shareout(Xd_0__inst_mult_24_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_25_25 (
// Equation(s):
// Xd_0__inst_mult_25_72  = SUM(( !Xd_0__inst_mult_25_16_q  $ (!Xd_0__inst_mult_25_17_q  $ (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_18_q )))) ) + ( Xd_0__inst_mult_25_70  ) + ( Xd_0__inst_mult_25_69  ))
// Xd_0__inst_mult_25_73  = CARRY(( !Xd_0__inst_mult_25_16_q  $ (!Xd_0__inst_mult_25_17_q  $ (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_18_q )))) ) + ( Xd_0__inst_mult_25_70  ) + ( Xd_0__inst_mult_25_69  ))
// Xd_0__inst_mult_25_74  = SHARE((!Xd_0__inst_mult_25_16_q  & (Xd_0__inst_mult_25_17_q  & (Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_18_q ))) # (Xd_0__inst_mult_25_16_q  & (((Xd_0__inst_mult_25_7_q  & Xd_0__inst_mult_25_18_q )) # (Xd_0__inst_mult_25_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_25_16_q ),
	.datab(!Xd_0__inst_mult_25_17_q ),
	.datac(!Xd_0__inst_mult_25_7_q ),
	.datad(!Xd_0__inst_mult_25_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_69 ),
	.sharein(Xd_0__inst_mult_25_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_72 ),
	.cout(Xd_0__inst_mult_25_73 ),
	.shareout(Xd_0__inst_mult_25_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_22_25 (
// Equation(s):
// Xd_0__inst_mult_22_72  = SUM(( !Xd_0__inst_mult_22_16_q  $ (!Xd_0__inst_mult_22_17_q  $ (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_18_q )))) ) + ( Xd_0__inst_mult_22_70  ) + ( Xd_0__inst_mult_22_69  ))
// Xd_0__inst_mult_22_73  = CARRY(( !Xd_0__inst_mult_22_16_q  $ (!Xd_0__inst_mult_22_17_q  $ (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_18_q )))) ) + ( Xd_0__inst_mult_22_70  ) + ( Xd_0__inst_mult_22_69  ))
// Xd_0__inst_mult_22_74  = SHARE((!Xd_0__inst_mult_22_16_q  & (Xd_0__inst_mult_22_17_q  & (Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_18_q ))) # (Xd_0__inst_mult_22_16_q  & (((Xd_0__inst_mult_22_7_q  & Xd_0__inst_mult_22_18_q )) # (Xd_0__inst_mult_22_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_22_16_q ),
	.datab(!Xd_0__inst_mult_22_17_q ),
	.datac(!Xd_0__inst_mult_22_7_q ),
	.datad(!Xd_0__inst_mult_22_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_69 ),
	.sharein(Xd_0__inst_mult_22_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_72 ),
	.cout(Xd_0__inst_mult_22_73 ),
	.shareout(Xd_0__inst_mult_22_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_23_25 (
// Equation(s):
// Xd_0__inst_mult_23_72  = SUM(( !Xd_0__inst_mult_23_16_q  $ (!Xd_0__inst_mult_23_17_q  $ (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_18_q )))) ) + ( Xd_0__inst_mult_23_70  ) + ( Xd_0__inst_mult_23_69  ))
// Xd_0__inst_mult_23_73  = CARRY(( !Xd_0__inst_mult_23_16_q  $ (!Xd_0__inst_mult_23_17_q  $ (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_18_q )))) ) + ( Xd_0__inst_mult_23_70  ) + ( Xd_0__inst_mult_23_69  ))
// Xd_0__inst_mult_23_74  = SHARE((!Xd_0__inst_mult_23_16_q  & (Xd_0__inst_mult_23_17_q  & (Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_18_q ))) # (Xd_0__inst_mult_23_16_q  & (((Xd_0__inst_mult_23_7_q  & Xd_0__inst_mult_23_18_q )) # (Xd_0__inst_mult_23_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_23_16_q ),
	.datab(!Xd_0__inst_mult_23_17_q ),
	.datac(!Xd_0__inst_mult_23_7_q ),
	.datad(!Xd_0__inst_mult_23_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_69 ),
	.sharein(Xd_0__inst_mult_23_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_72 ),
	.cout(Xd_0__inst_mult_23_73 ),
	.shareout(Xd_0__inst_mult_23_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_20_25 (
// Equation(s):
// Xd_0__inst_mult_20_72  = SUM(( !Xd_0__inst_mult_20_16_q  $ (!Xd_0__inst_mult_20_17_q  $ (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_18_q )))) ) + ( Xd_0__inst_mult_20_70  ) + ( Xd_0__inst_mult_20_69  ))
// Xd_0__inst_mult_20_73  = CARRY(( !Xd_0__inst_mult_20_16_q  $ (!Xd_0__inst_mult_20_17_q  $ (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_18_q )))) ) + ( Xd_0__inst_mult_20_70  ) + ( Xd_0__inst_mult_20_69  ))
// Xd_0__inst_mult_20_74  = SHARE((!Xd_0__inst_mult_20_16_q  & (Xd_0__inst_mult_20_17_q  & (Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_18_q ))) # (Xd_0__inst_mult_20_16_q  & (((Xd_0__inst_mult_20_7_q  & Xd_0__inst_mult_20_18_q )) # (Xd_0__inst_mult_20_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_20_16_q ),
	.datab(!Xd_0__inst_mult_20_17_q ),
	.datac(!Xd_0__inst_mult_20_7_q ),
	.datad(!Xd_0__inst_mult_20_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_69 ),
	.sharein(Xd_0__inst_mult_20_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_72 ),
	.cout(Xd_0__inst_mult_20_73 ),
	.shareout(Xd_0__inst_mult_20_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_21_25 (
// Equation(s):
// Xd_0__inst_mult_21_72  = SUM(( !Xd_0__inst_mult_21_16_q  $ (!Xd_0__inst_mult_21_17_q  $ (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_18_q )))) ) + ( Xd_0__inst_mult_21_70  ) + ( Xd_0__inst_mult_21_69  ))
// Xd_0__inst_mult_21_73  = CARRY(( !Xd_0__inst_mult_21_16_q  $ (!Xd_0__inst_mult_21_17_q  $ (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_18_q )))) ) + ( Xd_0__inst_mult_21_70  ) + ( Xd_0__inst_mult_21_69  ))
// Xd_0__inst_mult_21_74  = SHARE((!Xd_0__inst_mult_21_16_q  & (Xd_0__inst_mult_21_17_q  & (Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_18_q ))) # (Xd_0__inst_mult_21_16_q  & (((Xd_0__inst_mult_21_7_q  & Xd_0__inst_mult_21_18_q )) # (Xd_0__inst_mult_21_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_21_16_q ),
	.datab(!Xd_0__inst_mult_21_17_q ),
	.datac(!Xd_0__inst_mult_21_7_q ),
	.datad(!Xd_0__inst_mult_21_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_69 ),
	.sharein(Xd_0__inst_mult_21_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_72 ),
	.cout(Xd_0__inst_mult_21_73 ),
	.shareout(Xd_0__inst_mult_21_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_18_25 (
// Equation(s):
// Xd_0__inst_mult_18_72  = SUM(( !Xd_0__inst_mult_18_16_q  $ (!Xd_0__inst_mult_18_17_q  $ (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_18_q )))) ) + ( Xd_0__inst_mult_18_70  ) + ( Xd_0__inst_mult_18_69  ))
// Xd_0__inst_mult_18_73  = CARRY(( !Xd_0__inst_mult_18_16_q  $ (!Xd_0__inst_mult_18_17_q  $ (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_18_q )))) ) + ( Xd_0__inst_mult_18_70  ) + ( Xd_0__inst_mult_18_69  ))
// Xd_0__inst_mult_18_74  = SHARE((!Xd_0__inst_mult_18_16_q  & (Xd_0__inst_mult_18_17_q  & (Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_18_q ))) # (Xd_0__inst_mult_18_16_q  & (((Xd_0__inst_mult_18_7_q  & Xd_0__inst_mult_18_18_q )) # (Xd_0__inst_mult_18_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_18_16_q ),
	.datab(!Xd_0__inst_mult_18_17_q ),
	.datac(!Xd_0__inst_mult_18_7_q ),
	.datad(!Xd_0__inst_mult_18_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_69 ),
	.sharein(Xd_0__inst_mult_18_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_72 ),
	.cout(Xd_0__inst_mult_18_73 ),
	.shareout(Xd_0__inst_mult_18_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_19_25 (
// Equation(s):
// Xd_0__inst_mult_19_72  = SUM(( !Xd_0__inst_mult_19_16_q  $ (!Xd_0__inst_mult_19_17_q  $ (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_18_q )))) ) + ( Xd_0__inst_mult_19_70  ) + ( Xd_0__inst_mult_19_69  ))
// Xd_0__inst_mult_19_73  = CARRY(( !Xd_0__inst_mult_19_16_q  $ (!Xd_0__inst_mult_19_17_q  $ (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_18_q )))) ) + ( Xd_0__inst_mult_19_70  ) + ( Xd_0__inst_mult_19_69  ))
// Xd_0__inst_mult_19_74  = SHARE((!Xd_0__inst_mult_19_16_q  & (Xd_0__inst_mult_19_17_q  & (Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_18_q ))) # (Xd_0__inst_mult_19_16_q  & (((Xd_0__inst_mult_19_7_q  & Xd_0__inst_mult_19_18_q )) # (Xd_0__inst_mult_19_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_19_16_q ),
	.datab(!Xd_0__inst_mult_19_17_q ),
	.datac(!Xd_0__inst_mult_19_7_q ),
	.datad(!Xd_0__inst_mult_19_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_69 ),
	.sharein(Xd_0__inst_mult_19_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_72 ),
	.cout(Xd_0__inst_mult_19_73 ),
	.shareout(Xd_0__inst_mult_19_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_16_25 (
// Equation(s):
// Xd_0__inst_mult_16_72  = SUM(( !Xd_0__inst_mult_16_16_q  $ (!Xd_0__inst_mult_16_17_q  $ (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_18_q )))) ) + ( Xd_0__inst_mult_16_70  ) + ( Xd_0__inst_mult_16_69  ))
// Xd_0__inst_mult_16_73  = CARRY(( !Xd_0__inst_mult_16_16_q  $ (!Xd_0__inst_mult_16_17_q  $ (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_18_q )))) ) + ( Xd_0__inst_mult_16_70  ) + ( Xd_0__inst_mult_16_69  ))
// Xd_0__inst_mult_16_74  = SHARE((!Xd_0__inst_mult_16_16_q  & (Xd_0__inst_mult_16_17_q  & (Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_18_q ))) # (Xd_0__inst_mult_16_16_q  & (((Xd_0__inst_mult_16_7_q  & Xd_0__inst_mult_16_18_q )) # (Xd_0__inst_mult_16_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_16_16_q ),
	.datab(!Xd_0__inst_mult_16_17_q ),
	.datac(!Xd_0__inst_mult_16_7_q ),
	.datad(!Xd_0__inst_mult_16_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_69 ),
	.sharein(Xd_0__inst_mult_16_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_72 ),
	.cout(Xd_0__inst_mult_16_73 ),
	.shareout(Xd_0__inst_mult_16_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_17_25 (
// Equation(s):
// Xd_0__inst_mult_17_72  = SUM(( !Xd_0__inst_mult_17_16_q  $ (!Xd_0__inst_mult_17_17_q  $ (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_18_q )))) ) + ( Xd_0__inst_mult_17_70  ) + ( Xd_0__inst_mult_17_69  ))
// Xd_0__inst_mult_17_73  = CARRY(( !Xd_0__inst_mult_17_16_q  $ (!Xd_0__inst_mult_17_17_q  $ (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_18_q )))) ) + ( Xd_0__inst_mult_17_70  ) + ( Xd_0__inst_mult_17_69  ))
// Xd_0__inst_mult_17_74  = SHARE((!Xd_0__inst_mult_17_16_q  & (Xd_0__inst_mult_17_17_q  & (Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_18_q ))) # (Xd_0__inst_mult_17_16_q  & (((Xd_0__inst_mult_17_7_q  & Xd_0__inst_mult_17_18_q )) # (Xd_0__inst_mult_17_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_17_16_q ),
	.datab(!Xd_0__inst_mult_17_17_q ),
	.datac(!Xd_0__inst_mult_17_7_q ),
	.datad(!Xd_0__inst_mult_17_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_69 ),
	.sharein(Xd_0__inst_mult_17_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_72 ),
	.cout(Xd_0__inst_mult_17_73 ),
	.shareout(Xd_0__inst_mult_17_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_25 (
// Equation(s):
// Xd_0__inst_mult_14_72  = SUM(( !Xd_0__inst_mult_14_16_q  $ (!Xd_0__inst_mult_14_17_q  $ (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_18_q )))) ) + ( Xd_0__inst_mult_14_70  ) + ( Xd_0__inst_mult_14_69  ))
// Xd_0__inst_mult_14_73  = CARRY(( !Xd_0__inst_mult_14_16_q  $ (!Xd_0__inst_mult_14_17_q  $ (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_18_q )))) ) + ( Xd_0__inst_mult_14_70  ) + ( Xd_0__inst_mult_14_69  ))
// Xd_0__inst_mult_14_74  = SHARE((!Xd_0__inst_mult_14_16_q  & (Xd_0__inst_mult_14_17_q  & (Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_18_q ))) # (Xd_0__inst_mult_14_16_q  & (((Xd_0__inst_mult_14_7_q  & Xd_0__inst_mult_14_18_q )) # (Xd_0__inst_mult_14_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_14_16_q ),
	.datab(!Xd_0__inst_mult_14_17_q ),
	.datac(!Xd_0__inst_mult_14_7_q ),
	.datad(!Xd_0__inst_mult_14_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_69 ),
	.sharein(Xd_0__inst_mult_14_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_72 ),
	.cout(Xd_0__inst_mult_14_73 ),
	.shareout(Xd_0__inst_mult_14_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_25 (
// Equation(s):
// Xd_0__inst_mult_15_72  = SUM(( !Xd_0__inst_mult_15_16_q  $ (!Xd_0__inst_mult_15_17_q  $ (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_18_q )))) ) + ( Xd_0__inst_mult_15_70  ) + ( Xd_0__inst_mult_15_69  ))
// Xd_0__inst_mult_15_73  = CARRY(( !Xd_0__inst_mult_15_16_q  $ (!Xd_0__inst_mult_15_17_q  $ (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_18_q )))) ) + ( Xd_0__inst_mult_15_70  ) + ( Xd_0__inst_mult_15_69  ))
// Xd_0__inst_mult_15_74  = SHARE((!Xd_0__inst_mult_15_16_q  & (Xd_0__inst_mult_15_17_q  & (Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_18_q ))) # (Xd_0__inst_mult_15_16_q  & (((Xd_0__inst_mult_15_7_q  & Xd_0__inst_mult_15_18_q )) # (Xd_0__inst_mult_15_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_15_16_q ),
	.datab(!Xd_0__inst_mult_15_17_q ),
	.datac(!Xd_0__inst_mult_15_7_q ),
	.datad(!Xd_0__inst_mult_15_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_69 ),
	.sharein(Xd_0__inst_mult_15_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_72 ),
	.cout(Xd_0__inst_mult_15_73 ),
	.shareout(Xd_0__inst_mult_15_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_25 (
// Equation(s):
// Xd_0__inst_mult_12_72  = SUM(( !Xd_0__inst_mult_12_16_q  $ (!Xd_0__inst_mult_12_17_q  $ (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_18_q )))) ) + ( Xd_0__inst_mult_12_70  ) + ( Xd_0__inst_mult_12_69  ))
// Xd_0__inst_mult_12_73  = CARRY(( !Xd_0__inst_mult_12_16_q  $ (!Xd_0__inst_mult_12_17_q  $ (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_18_q )))) ) + ( Xd_0__inst_mult_12_70  ) + ( Xd_0__inst_mult_12_69  ))
// Xd_0__inst_mult_12_74  = SHARE((!Xd_0__inst_mult_12_16_q  & (Xd_0__inst_mult_12_17_q  & (Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_18_q ))) # (Xd_0__inst_mult_12_16_q  & (((Xd_0__inst_mult_12_7_q  & Xd_0__inst_mult_12_18_q )) # (Xd_0__inst_mult_12_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_12_16_q ),
	.datab(!Xd_0__inst_mult_12_17_q ),
	.datac(!Xd_0__inst_mult_12_7_q ),
	.datad(!Xd_0__inst_mult_12_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_69 ),
	.sharein(Xd_0__inst_mult_12_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_72 ),
	.cout(Xd_0__inst_mult_12_73 ),
	.shareout(Xd_0__inst_mult_12_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_25 (
// Equation(s):
// Xd_0__inst_mult_13_72  = SUM(( !Xd_0__inst_mult_13_16_q  $ (!Xd_0__inst_mult_13_17_q  $ (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_18_q )))) ) + ( Xd_0__inst_mult_13_70  ) + ( Xd_0__inst_mult_13_69  ))
// Xd_0__inst_mult_13_73  = CARRY(( !Xd_0__inst_mult_13_16_q  $ (!Xd_0__inst_mult_13_17_q  $ (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_18_q )))) ) + ( Xd_0__inst_mult_13_70  ) + ( Xd_0__inst_mult_13_69  ))
// Xd_0__inst_mult_13_74  = SHARE((!Xd_0__inst_mult_13_16_q  & (Xd_0__inst_mult_13_17_q  & (Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_18_q ))) # (Xd_0__inst_mult_13_16_q  & (((Xd_0__inst_mult_13_7_q  & Xd_0__inst_mult_13_18_q )) # (Xd_0__inst_mult_13_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_13_16_q ),
	.datab(!Xd_0__inst_mult_13_17_q ),
	.datac(!Xd_0__inst_mult_13_7_q ),
	.datad(!Xd_0__inst_mult_13_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_69 ),
	.sharein(Xd_0__inst_mult_13_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_72 ),
	.cout(Xd_0__inst_mult_13_73 ),
	.shareout(Xd_0__inst_mult_13_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_25 (
// Equation(s):
// Xd_0__inst_mult_10_72  = SUM(( !Xd_0__inst_mult_10_16_q  $ (!Xd_0__inst_mult_10_17_q  $ (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_18_q )))) ) + ( Xd_0__inst_mult_10_70  ) + ( Xd_0__inst_mult_10_69  ))
// Xd_0__inst_mult_10_73  = CARRY(( !Xd_0__inst_mult_10_16_q  $ (!Xd_0__inst_mult_10_17_q  $ (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_18_q )))) ) + ( Xd_0__inst_mult_10_70  ) + ( Xd_0__inst_mult_10_69  ))
// Xd_0__inst_mult_10_74  = SHARE((!Xd_0__inst_mult_10_16_q  & (Xd_0__inst_mult_10_17_q  & (Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_18_q ))) # (Xd_0__inst_mult_10_16_q  & (((Xd_0__inst_mult_10_7_q  & Xd_0__inst_mult_10_18_q )) # (Xd_0__inst_mult_10_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_10_16_q ),
	.datab(!Xd_0__inst_mult_10_17_q ),
	.datac(!Xd_0__inst_mult_10_7_q ),
	.datad(!Xd_0__inst_mult_10_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_69 ),
	.sharein(Xd_0__inst_mult_10_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_72 ),
	.cout(Xd_0__inst_mult_10_73 ),
	.shareout(Xd_0__inst_mult_10_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_25 (
// Equation(s):
// Xd_0__inst_mult_11_72  = SUM(( !Xd_0__inst_mult_11_16_q  $ (!Xd_0__inst_mult_11_17_q  $ (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_18_q )))) ) + ( Xd_0__inst_mult_11_70  ) + ( Xd_0__inst_mult_11_69  ))
// Xd_0__inst_mult_11_73  = CARRY(( !Xd_0__inst_mult_11_16_q  $ (!Xd_0__inst_mult_11_17_q  $ (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_18_q )))) ) + ( Xd_0__inst_mult_11_70  ) + ( Xd_0__inst_mult_11_69  ))
// Xd_0__inst_mult_11_74  = SHARE((!Xd_0__inst_mult_11_16_q  & (Xd_0__inst_mult_11_17_q  & (Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_18_q ))) # (Xd_0__inst_mult_11_16_q  & (((Xd_0__inst_mult_11_7_q  & Xd_0__inst_mult_11_18_q )) # (Xd_0__inst_mult_11_17_q 
// ))))

	.dataa(!Xd_0__inst_mult_11_16_q ),
	.datab(!Xd_0__inst_mult_11_17_q ),
	.datac(!Xd_0__inst_mult_11_7_q ),
	.datad(!Xd_0__inst_mult_11_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_69 ),
	.sharein(Xd_0__inst_mult_11_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_72 ),
	.cout(Xd_0__inst_mult_11_73 ),
	.shareout(Xd_0__inst_mult_11_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_25 (
// Equation(s):
// Xd_0__inst_mult_8_72  = SUM(( !Xd_0__inst_mult_8_16_q  $ (!Xd_0__inst_mult_8_17_q  $ (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_18_q )))) ) + ( Xd_0__inst_mult_8_70  ) + ( Xd_0__inst_mult_8_69  ))
// Xd_0__inst_mult_8_73  = CARRY(( !Xd_0__inst_mult_8_16_q  $ (!Xd_0__inst_mult_8_17_q  $ (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_18_q )))) ) + ( Xd_0__inst_mult_8_70  ) + ( Xd_0__inst_mult_8_69  ))
// Xd_0__inst_mult_8_74  = SHARE((!Xd_0__inst_mult_8_16_q  & (Xd_0__inst_mult_8_17_q  & (Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_18_q ))) # (Xd_0__inst_mult_8_16_q  & (((Xd_0__inst_mult_8_7_q  & Xd_0__inst_mult_8_18_q )) # (Xd_0__inst_mult_8_17_q ))))

	.dataa(!Xd_0__inst_mult_8_16_q ),
	.datab(!Xd_0__inst_mult_8_17_q ),
	.datac(!Xd_0__inst_mult_8_7_q ),
	.datad(!Xd_0__inst_mult_8_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_69 ),
	.sharein(Xd_0__inst_mult_8_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_72 ),
	.cout(Xd_0__inst_mult_8_73 ),
	.shareout(Xd_0__inst_mult_8_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_25 (
// Equation(s):
// Xd_0__inst_mult_9_72  = SUM(( !Xd_0__inst_mult_9_16_q  $ (!Xd_0__inst_mult_9_17_q  $ (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_18_q )))) ) + ( Xd_0__inst_mult_9_70  ) + ( Xd_0__inst_mult_9_69  ))
// Xd_0__inst_mult_9_73  = CARRY(( !Xd_0__inst_mult_9_16_q  $ (!Xd_0__inst_mult_9_17_q  $ (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_18_q )))) ) + ( Xd_0__inst_mult_9_70  ) + ( Xd_0__inst_mult_9_69  ))
// Xd_0__inst_mult_9_74  = SHARE((!Xd_0__inst_mult_9_16_q  & (Xd_0__inst_mult_9_17_q  & (Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_18_q ))) # (Xd_0__inst_mult_9_16_q  & (((Xd_0__inst_mult_9_7_q  & Xd_0__inst_mult_9_18_q )) # (Xd_0__inst_mult_9_17_q ))))

	.dataa(!Xd_0__inst_mult_9_16_q ),
	.datab(!Xd_0__inst_mult_9_17_q ),
	.datac(!Xd_0__inst_mult_9_7_q ),
	.datad(!Xd_0__inst_mult_9_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_69 ),
	.sharein(Xd_0__inst_mult_9_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_72 ),
	.cout(Xd_0__inst_mult_9_73 ),
	.shareout(Xd_0__inst_mult_9_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_25 (
// Equation(s):
// Xd_0__inst_mult_6_72  = SUM(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q  $ (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_18_q )))) ) + ( Xd_0__inst_mult_6_70  ) + ( Xd_0__inst_mult_6_69  ))
// Xd_0__inst_mult_6_73  = CARRY(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q  $ (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_18_q )))) ) + ( Xd_0__inst_mult_6_70  ) + ( Xd_0__inst_mult_6_69  ))
// Xd_0__inst_mult_6_74  = SHARE((!Xd_0__inst_mult_6_16_q  & (Xd_0__inst_mult_6_17_q  & (Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_18_q ))) # (Xd_0__inst_mult_6_16_q  & (((Xd_0__inst_mult_6_7_q  & Xd_0__inst_mult_6_18_q )) # (Xd_0__inst_mult_6_17_q ))))

	.dataa(!Xd_0__inst_mult_6_16_q ),
	.datab(!Xd_0__inst_mult_6_17_q ),
	.datac(!Xd_0__inst_mult_6_7_q ),
	.datad(!Xd_0__inst_mult_6_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_69 ),
	.sharein(Xd_0__inst_mult_6_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_72 ),
	.cout(Xd_0__inst_mult_6_73 ),
	.shareout(Xd_0__inst_mult_6_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_25 (
// Equation(s):
// Xd_0__inst_mult_7_72  = SUM(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q  $ (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_18_q )))) ) + ( Xd_0__inst_mult_7_70  ) + ( Xd_0__inst_mult_7_69  ))
// Xd_0__inst_mult_7_73  = CARRY(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q  $ (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_18_q )))) ) + ( Xd_0__inst_mult_7_70  ) + ( Xd_0__inst_mult_7_69  ))
// Xd_0__inst_mult_7_74  = SHARE((!Xd_0__inst_mult_7_16_q  & (Xd_0__inst_mult_7_17_q  & (Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_18_q ))) # (Xd_0__inst_mult_7_16_q  & (((Xd_0__inst_mult_7_7_q  & Xd_0__inst_mult_7_18_q )) # (Xd_0__inst_mult_7_17_q ))))

	.dataa(!Xd_0__inst_mult_7_16_q ),
	.datab(!Xd_0__inst_mult_7_17_q ),
	.datac(!Xd_0__inst_mult_7_7_q ),
	.datad(!Xd_0__inst_mult_7_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_69 ),
	.sharein(Xd_0__inst_mult_7_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_72 ),
	.cout(Xd_0__inst_mult_7_73 ),
	.shareout(Xd_0__inst_mult_7_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_25 (
// Equation(s):
// Xd_0__inst_mult_4_72  = SUM(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q  $ (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_18_q )))) ) + ( Xd_0__inst_mult_4_70  ) + ( Xd_0__inst_mult_4_69  ))
// Xd_0__inst_mult_4_73  = CARRY(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q  $ (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_18_q )))) ) + ( Xd_0__inst_mult_4_70  ) + ( Xd_0__inst_mult_4_69  ))
// Xd_0__inst_mult_4_74  = SHARE((!Xd_0__inst_mult_4_16_q  & (Xd_0__inst_mult_4_17_q  & (Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_18_q ))) # (Xd_0__inst_mult_4_16_q  & (((Xd_0__inst_mult_4_7_q  & Xd_0__inst_mult_4_18_q )) # (Xd_0__inst_mult_4_17_q ))))

	.dataa(!Xd_0__inst_mult_4_16_q ),
	.datab(!Xd_0__inst_mult_4_17_q ),
	.datac(!Xd_0__inst_mult_4_7_q ),
	.datad(!Xd_0__inst_mult_4_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_69 ),
	.sharein(Xd_0__inst_mult_4_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_72 ),
	.cout(Xd_0__inst_mult_4_73 ),
	.shareout(Xd_0__inst_mult_4_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_25 (
// Equation(s):
// Xd_0__inst_mult_5_72  = SUM(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q  $ (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_18_q )))) ) + ( Xd_0__inst_mult_5_70  ) + ( Xd_0__inst_mult_5_69  ))
// Xd_0__inst_mult_5_73  = CARRY(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q  $ (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_18_q )))) ) + ( Xd_0__inst_mult_5_70  ) + ( Xd_0__inst_mult_5_69  ))
// Xd_0__inst_mult_5_74  = SHARE((!Xd_0__inst_mult_5_16_q  & (Xd_0__inst_mult_5_17_q  & (Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_18_q ))) # (Xd_0__inst_mult_5_16_q  & (((Xd_0__inst_mult_5_7_q  & Xd_0__inst_mult_5_18_q )) # (Xd_0__inst_mult_5_17_q ))))

	.dataa(!Xd_0__inst_mult_5_16_q ),
	.datab(!Xd_0__inst_mult_5_17_q ),
	.datac(!Xd_0__inst_mult_5_7_q ),
	.datad(!Xd_0__inst_mult_5_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_69 ),
	.sharein(Xd_0__inst_mult_5_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_72 ),
	.cout(Xd_0__inst_mult_5_73 ),
	.shareout(Xd_0__inst_mult_5_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_25 (
// Equation(s):
// Xd_0__inst_mult_2_72  = SUM(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q  $ (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_18_q )))) ) + ( Xd_0__inst_mult_2_70  ) + ( Xd_0__inst_mult_2_69  ))
// Xd_0__inst_mult_2_73  = CARRY(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q  $ (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_18_q )))) ) + ( Xd_0__inst_mult_2_70  ) + ( Xd_0__inst_mult_2_69  ))
// Xd_0__inst_mult_2_74  = SHARE((!Xd_0__inst_mult_2_16_q  & (Xd_0__inst_mult_2_17_q  & (Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_18_q ))) # (Xd_0__inst_mult_2_16_q  & (((Xd_0__inst_mult_2_7_q  & Xd_0__inst_mult_2_18_q )) # (Xd_0__inst_mult_2_17_q ))))

	.dataa(!Xd_0__inst_mult_2_16_q ),
	.datab(!Xd_0__inst_mult_2_17_q ),
	.datac(!Xd_0__inst_mult_2_7_q ),
	.datad(!Xd_0__inst_mult_2_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_69 ),
	.sharein(Xd_0__inst_mult_2_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_72 ),
	.cout(Xd_0__inst_mult_2_73 ),
	.shareout(Xd_0__inst_mult_2_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_25 (
// Equation(s):
// Xd_0__inst_mult_3_72  = SUM(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q  $ (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_18_q )))) ) + ( Xd_0__inst_mult_3_70  ) + ( Xd_0__inst_mult_3_69  ))
// Xd_0__inst_mult_3_73  = CARRY(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q  $ (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_18_q )))) ) + ( Xd_0__inst_mult_3_70  ) + ( Xd_0__inst_mult_3_69  ))
// Xd_0__inst_mult_3_74  = SHARE((!Xd_0__inst_mult_3_16_q  & (Xd_0__inst_mult_3_17_q  & (Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_18_q ))) # (Xd_0__inst_mult_3_16_q  & (((Xd_0__inst_mult_3_7_q  & Xd_0__inst_mult_3_18_q )) # (Xd_0__inst_mult_3_17_q ))))

	.dataa(!Xd_0__inst_mult_3_16_q ),
	.datab(!Xd_0__inst_mult_3_17_q ),
	.datac(!Xd_0__inst_mult_3_7_q ),
	.datad(!Xd_0__inst_mult_3_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_69 ),
	.sharein(Xd_0__inst_mult_3_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_72 ),
	.cout(Xd_0__inst_mult_3_73 ),
	.shareout(Xd_0__inst_mult_3_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_25 (
// Equation(s):
// Xd_0__inst_mult_0_72  = SUM(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q  $ (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_18_q )))) ) + ( Xd_0__inst_mult_0_70  ) + ( Xd_0__inst_mult_0_69  ))
// Xd_0__inst_mult_0_73  = CARRY(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q  $ (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_18_q )))) ) + ( Xd_0__inst_mult_0_70  ) + ( Xd_0__inst_mult_0_69  ))
// Xd_0__inst_mult_0_74  = SHARE((!Xd_0__inst_mult_0_16_q  & (Xd_0__inst_mult_0_17_q  & (Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_18_q ))) # (Xd_0__inst_mult_0_16_q  & (((Xd_0__inst_mult_0_7_q  & Xd_0__inst_mult_0_18_q )) # (Xd_0__inst_mult_0_17_q ))))

	.dataa(!Xd_0__inst_mult_0_16_q ),
	.datab(!Xd_0__inst_mult_0_17_q ),
	.datac(!Xd_0__inst_mult_0_7_q ),
	.datad(!Xd_0__inst_mult_0_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_69 ),
	.sharein(Xd_0__inst_mult_0_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_72 ),
	.cout(Xd_0__inst_mult_0_73 ),
	.shareout(Xd_0__inst_mult_0_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_25 (
// Equation(s):
// Xd_0__inst_mult_1_72  = SUM(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q  $ (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_18_q )))) ) + ( Xd_0__inst_mult_1_70  ) + ( Xd_0__inst_mult_1_69  ))
// Xd_0__inst_mult_1_73  = CARRY(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q  $ (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_18_q )))) ) + ( Xd_0__inst_mult_1_70  ) + ( Xd_0__inst_mult_1_69  ))
// Xd_0__inst_mult_1_74  = SHARE((!Xd_0__inst_mult_1_16_q  & (Xd_0__inst_mult_1_17_q  & (Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_18_q ))) # (Xd_0__inst_mult_1_16_q  & (((Xd_0__inst_mult_1_7_q  & Xd_0__inst_mult_1_18_q )) # (Xd_0__inst_mult_1_17_q ))))

	.dataa(!Xd_0__inst_mult_1_16_q ),
	.datab(!Xd_0__inst_mult_1_17_q ),
	.datac(!Xd_0__inst_mult_1_7_q ),
	.datad(!Xd_0__inst_mult_1_18_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_69 ),
	.sharein(Xd_0__inst_mult_1_70 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_72 ),
	.cout(Xd_0__inst_mult_1_73 ),
	.shareout(Xd_0__inst_mult_1_74 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_28_26 (
// Equation(s):
// Xd_0__inst_mult_28_76  = SUM(( !Xd_0__inst_mult_28_20_q  $ (((!Xd_0__inst_mult_28_19_q ) # (!Xd_0__inst_mult_28_18_q ))) ) + ( Xd_0__inst_mult_28_74  ) + ( Xd_0__inst_mult_28_73  ))
// Xd_0__inst_mult_28_77  = CARRY(( !Xd_0__inst_mult_28_20_q  $ (((!Xd_0__inst_mult_28_19_q ) # (!Xd_0__inst_mult_28_18_q ))) ) + ( Xd_0__inst_mult_28_74  ) + ( Xd_0__inst_mult_28_73  ))
// Xd_0__inst_mult_28_78  = SHARE((Xd_0__inst_mult_28_19_q  & (Xd_0__inst_mult_28_18_q  & Xd_0__inst_mult_28_20_q )))

	.dataa(!Xd_0__inst_mult_28_19_q ),
	.datab(!Xd_0__inst_mult_28_18_q ),
	.datac(!Xd_0__inst_mult_28_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_73 ),
	.sharein(Xd_0__inst_mult_28_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_76 ),
	.cout(Xd_0__inst_mult_28_77 ),
	.shareout(Xd_0__inst_mult_28_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_29_26 (
// Equation(s):
// Xd_0__inst_mult_29_76  = SUM(( !Xd_0__inst_mult_29_20_q  $ (((!Xd_0__inst_mult_29_19_q ) # (!Xd_0__inst_mult_29_18_q ))) ) + ( Xd_0__inst_mult_29_74  ) + ( Xd_0__inst_mult_29_73  ))
// Xd_0__inst_mult_29_77  = CARRY(( !Xd_0__inst_mult_29_20_q  $ (((!Xd_0__inst_mult_29_19_q ) # (!Xd_0__inst_mult_29_18_q ))) ) + ( Xd_0__inst_mult_29_74  ) + ( Xd_0__inst_mult_29_73  ))
// Xd_0__inst_mult_29_78  = SHARE((Xd_0__inst_mult_29_19_q  & (Xd_0__inst_mult_29_18_q  & Xd_0__inst_mult_29_20_q )))

	.dataa(!Xd_0__inst_mult_29_19_q ),
	.datab(!Xd_0__inst_mult_29_18_q ),
	.datac(!Xd_0__inst_mult_29_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_73 ),
	.sharein(Xd_0__inst_mult_29_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_76 ),
	.cout(Xd_0__inst_mult_29_77 ),
	.shareout(Xd_0__inst_mult_29_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_26_26 (
// Equation(s):
// Xd_0__inst_mult_26_76  = SUM(( !Xd_0__inst_mult_26_20_q  $ (((!Xd_0__inst_mult_26_19_q ) # (!Xd_0__inst_mult_26_18_q ))) ) + ( Xd_0__inst_mult_26_74  ) + ( Xd_0__inst_mult_26_73  ))
// Xd_0__inst_mult_26_77  = CARRY(( !Xd_0__inst_mult_26_20_q  $ (((!Xd_0__inst_mult_26_19_q ) # (!Xd_0__inst_mult_26_18_q ))) ) + ( Xd_0__inst_mult_26_74  ) + ( Xd_0__inst_mult_26_73  ))
// Xd_0__inst_mult_26_78  = SHARE((Xd_0__inst_mult_26_19_q  & (Xd_0__inst_mult_26_18_q  & Xd_0__inst_mult_26_20_q )))

	.dataa(!Xd_0__inst_mult_26_19_q ),
	.datab(!Xd_0__inst_mult_26_18_q ),
	.datac(!Xd_0__inst_mult_26_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_73 ),
	.sharein(Xd_0__inst_mult_26_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_76 ),
	.cout(Xd_0__inst_mult_26_77 ),
	.shareout(Xd_0__inst_mult_26_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_27_26 (
// Equation(s):
// Xd_0__inst_mult_27_76  = SUM(( !Xd_0__inst_mult_27_20_q  $ (((!Xd_0__inst_mult_27_19_q ) # (!Xd_0__inst_mult_27_18_q ))) ) + ( Xd_0__inst_mult_27_74  ) + ( Xd_0__inst_mult_27_73  ))
// Xd_0__inst_mult_27_77  = CARRY(( !Xd_0__inst_mult_27_20_q  $ (((!Xd_0__inst_mult_27_19_q ) # (!Xd_0__inst_mult_27_18_q ))) ) + ( Xd_0__inst_mult_27_74  ) + ( Xd_0__inst_mult_27_73  ))
// Xd_0__inst_mult_27_78  = SHARE((Xd_0__inst_mult_27_19_q  & (Xd_0__inst_mult_27_18_q  & Xd_0__inst_mult_27_20_q )))

	.dataa(!Xd_0__inst_mult_27_19_q ),
	.datab(!Xd_0__inst_mult_27_18_q ),
	.datac(!Xd_0__inst_mult_27_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_73 ),
	.sharein(Xd_0__inst_mult_27_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_76 ),
	.cout(Xd_0__inst_mult_27_77 ),
	.shareout(Xd_0__inst_mult_27_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_24_26 (
// Equation(s):
// Xd_0__inst_mult_24_76  = SUM(( !Xd_0__inst_mult_24_20_q  $ (((!Xd_0__inst_mult_24_19_q ) # (!Xd_0__inst_mult_24_18_q ))) ) + ( Xd_0__inst_mult_24_74  ) + ( Xd_0__inst_mult_24_73  ))
// Xd_0__inst_mult_24_77  = CARRY(( !Xd_0__inst_mult_24_20_q  $ (((!Xd_0__inst_mult_24_19_q ) # (!Xd_0__inst_mult_24_18_q ))) ) + ( Xd_0__inst_mult_24_74  ) + ( Xd_0__inst_mult_24_73  ))
// Xd_0__inst_mult_24_78  = SHARE((Xd_0__inst_mult_24_19_q  & (Xd_0__inst_mult_24_18_q  & Xd_0__inst_mult_24_20_q )))

	.dataa(!Xd_0__inst_mult_24_19_q ),
	.datab(!Xd_0__inst_mult_24_18_q ),
	.datac(!Xd_0__inst_mult_24_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_73 ),
	.sharein(Xd_0__inst_mult_24_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_76 ),
	.cout(Xd_0__inst_mult_24_77 ),
	.shareout(Xd_0__inst_mult_24_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_25_26 (
// Equation(s):
// Xd_0__inst_mult_25_76  = SUM(( !Xd_0__inst_mult_25_20_q  $ (((!Xd_0__inst_mult_25_19_q ) # (!Xd_0__inst_mult_25_18_q ))) ) + ( Xd_0__inst_mult_25_74  ) + ( Xd_0__inst_mult_25_73  ))
// Xd_0__inst_mult_25_77  = CARRY(( !Xd_0__inst_mult_25_20_q  $ (((!Xd_0__inst_mult_25_19_q ) # (!Xd_0__inst_mult_25_18_q ))) ) + ( Xd_0__inst_mult_25_74  ) + ( Xd_0__inst_mult_25_73  ))
// Xd_0__inst_mult_25_78  = SHARE((Xd_0__inst_mult_25_19_q  & (Xd_0__inst_mult_25_18_q  & Xd_0__inst_mult_25_20_q )))

	.dataa(!Xd_0__inst_mult_25_19_q ),
	.datab(!Xd_0__inst_mult_25_18_q ),
	.datac(!Xd_0__inst_mult_25_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_73 ),
	.sharein(Xd_0__inst_mult_25_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_76 ),
	.cout(Xd_0__inst_mult_25_77 ),
	.shareout(Xd_0__inst_mult_25_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_22_26 (
// Equation(s):
// Xd_0__inst_mult_22_76  = SUM(( !Xd_0__inst_mult_22_20_q  $ (((!Xd_0__inst_mult_22_19_q ) # (!Xd_0__inst_mult_22_18_q ))) ) + ( Xd_0__inst_mult_22_74  ) + ( Xd_0__inst_mult_22_73  ))
// Xd_0__inst_mult_22_77  = CARRY(( !Xd_0__inst_mult_22_20_q  $ (((!Xd_0__inst_mult_22_19_q ) # (!Xd_0__inst_mult_22_18_q ))) ) + ( Xd_0__inst_mult_22_74  ) + ( Xd_0__inst_mult_22_73  ))
// Xd_0__inst_mult_22_78  = SHARE((Xd_0__inst_mult_22_19_q  & (Xd_0__inst_mult_22_18_q  & Xd_0__inst_mult_22_20_q )))

	.dataa(!Xd_0__inst_mult_22_19_q ),
	.datab(!Xd_0__inst_mult_22_18_q ),
	.datac(!Xd_0__inst_mult_22_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_73 ),
	.sharein(Xd_0__inst_mult_22_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_76 ),
	.cout(Xd_0__inst_mult_22_77 ),
	.shareout(Xd_0__inst_mult_22_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_23_26 (
// Equation(s):
// Xd_0__inst_mult_23_76  = SUM(( !Xd_0__inst_mult_23_20_q  $ (((!Xd_0__inst_mult_23_19_q ) # (!Xd_0__inst_mult_23_18_q ))) ) + ( Xd_0__inst_mult_23_74  ) + ( Xd_0__inst_mult_23_73  ))
// Xd_0__inst_mult_23_77  = CARRY(( !Xd_0__inst_mult_23_20_q  $ (((!Xd_0__inst_mult_23_19_q ) # (!Xd_0__inst_mult_23_18_q ))) ) + ( Xd_0__inst_mult_23_74  ) + ( Xd_0__inst_mult_23_73  ))
// Xd_0__inst_mult_23_78  = SHARE((Xd_0__inst_mult_23_19_q  & (Xd_0__inst_mult_23_18_q  & Xd_0__inst_mult_23_20_q )))

	.dataa(!Xd_0__inst_mult_23_19_q ),
	.datab(!Xd_0__inst_mult_23_18_q ),
	.datac(!Xd_0__inst_mult_23_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_73 ),
	.sharein(Xd_0__inst_mult_23_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_76 ),
	.cout(Xd_0__inst_mult_23_77 ),
	.shareout(Xd_0__inst_mult_23_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_20_26 (
// Equation(s):
// Xd_0__inst_mult_20_76  = SUM(( !Xd_0__inst_mult_20_20_q  $ (((!Xd_0__inst_mult_20_19_q ) # (!Xd_0__inst_mult_20_18_q ))) ) + ( Xd_0__inst_mult_20_74  ) + ( Xd_0__inst_mult_20_73  ))
// Xd_0__inst_mult_20_77  = CARRY(( !Xd_0__inst_mult_20_20_q  $ (((!Xd_0__inst_mult_20_19_q ) # (!Xd_0__inst_mult_20_18_q ))) ) + ( Xd_0__inst_mult_20_74  ) + ( Xd_0__inst_mult_20_73  ))
// Xd_0__inst_mult_20_78  = SHARE((Xd_0__inst_mult_20_19_q  & (Xd_0__inst_mult_20_18_q  & Xd_0__inst_mult_20_20_q )))

	.dataa(!Xd_0__inst_mult_20_19_q ),
	.datab(!Xd_0__inst_mult_20_18_q ),
	.datac(!Xd_0__inst_mult_20_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_73 ),
	.sharein(Xd_0__inst_mult_20_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_76 ),
	.cout(Xd_0__inst_mult_20_77 ),
	.shareout(Xd_0__inst_mult_20_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_21_26 (
// Equation(s):
// Xd_0__inst_mult_21_76  = SUM(( !Xd_0__inst_mult_21_20_q  $ (((!Xd_0__inst_mult_21_19_q ) # (!Xd_0__inst_mult_21_18_q ))) ) + ( Xd_0__inst_mult_21_74  ) + ( Xd_0__inst_mult_21_73  ))
// Xd_0__inst_mult_21_77  = CARRY(( !Xd_0__inst_mult_21_20_q  $ (((!Xd_0__inst_mult_21_19_q ) # (!Xd_0__inst_mult_21_18_q ))) ) + ( Xd_0__inst_mult_21_74  ) + ( Xd_0__inst_mult_21_73  ))
// Xd_0__inst_mult_21_78  = SHARE((Xd_0__inst_mult_21_19_q  & (Xd_0__inst_mult_21_18_q  & Xd_0__inst_mult_21_20_q )))

	.dataa(!Xd_0__inst_mult_21_19_q ),
	.datab(!Xd_0__inst_mult_21_18_q ),
	.datac(!Xd_0__inst_mult_21_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_73 ),
	.sharein(Xd_0__inst_mult_21_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_76 ),
	.cout(Xd_0__inst_mult_21_77 ),
	.shareout(Xd_0__inst_mult_21_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_18_26 (
// Equation(s):
// Xd_0__inst_mult_18_76  = SUM(( !Xd_0__inst_mult_18_20_q  $ (((!Xd_0__inst_mult_18_19_q ) # (!Xd_0__inst_mult_18_18_q ))) ) + ( Xd_0__inst_mult_18_74  ) + ( Xd_0__inst_mult_18_73  ))
// Xd_0__inst_mult_18_77  = CARRY(( !Xd_0__inst_mult_18_20_q  $ (((!Xd_0__inst_mult_18_19_q ) # (!Xd_0__inst_mult_18_18_q ))) ) + ( Xd_0__inst_mult_18_74  ) + ( Xd_0__inst_mult_18_73  ))
// Xd_0__inst_mult_18_78  = SHARE((Xd_0__inst_mult_18_19_q  & (Xd_0__inst_mult_18_18_q  & Xd_0__inst_mult_18_20_q )))

	.dataa(!Xd_0__inst_mult_18_19_q ),
	.datab(!Xd_0__inst_mult_18_18_q ),
	.datac(!Xd_0__inst_mult_18_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_73 ),
	.sharein(Xd_0__inst_mult_18_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_76 ),
	.cout(Xd_0__inst_mult_18_77 ),
	.shareout(Xd_0__inst_mult_18_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_19_26 (
// Equation(s):
// Xd_0__inst_mult_19_76  = SUM(( !Xd_0__inst_mult_19_20_q  $ (((!Xd_0__inst_mult_19_19_q ) # (!Xd_0__inst_mult_19_18_q ))) ) + ( Xd_0__inst_mult_19_74  ) + ( Xd_0__inst_mult_19_73  ))
// Xd_0__inst_mult_19_77  = CARRY(( !Xd_0__inst_mult_19_20_q  $ (((!Xd_0__inst_mult_19_19_q ) # (!Xd_0__inst_mult_19_18_q ))) ) + ( Xd_0__inst_mult_19_74  ) + ( Xd_0__inst_mult_19_73  ))
// Xd_0__inst_mult_19_78  = SHARE((Xd_0__inst_mult_19_19_q  & (Xd_0__inst_mult_19_18_q  & Xd_0__inst_mult_19_20_q )))

	.dataa(!Xd_0__inst_mult_19_19_q ),
	.datab(!Xd_0__inst_mult_19_18_q ),
	.datac(!Xd_0__inst_mult_19_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_73 ),
	.sharein(Xd_0__inst_mult_19_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_76 ),
	.cout(Xd_0__inst_mult_19_77 ),
	.shareout(Xd_0__inst_mult_19_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_16_26 (
// Equation(s):
// Xd_0__inst_mult_16_76  = SUM(( !Xd_0__inst_mult_16_20_q  $ (((!Xd_0__inst_mult_16_19_q ) # (!Xd_0__inst_mult_16_18_q ))) ) + ( Xd_0__inst_mult_16_74  ) + ( Xd_0__inst_mult_16_73  ))
// Xd_0__inst_mult_16_77  = CARRY(( !Xd_0__inst_mult_16_20_q  $ (((!Xd_0__inst_mult_16_19_q ) # (!Xd_0__inst_mult_16_18_q ))) ) + ( Xd_0__inst_mult_16_74  ) + ( Xd_0__inst_mult_16_73  ))
// Xd_0__inst_mult_16_78  = SHARE((Xd_0__inst_mult_16_19_q  & (Xd_0__inst_mult_16_18_q  & Xd_0__inst_mult_16_20_q )))

	.dataa(!Xd_0__inst_mult_16_19_q ),
	.datab(!Xd_0__inst_mult_16_18_q ),
	.datac(!Xd_0__inst_mult_16_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_73 ),
	.sharein(Xd_0__inst_mult_16_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_76 ),
	.cout(Xd_0__inst_mult_16_77 ),
	.shareout(Xd_0__inst_mult_16_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_17_26 (
// Equation(s):
// Xd_0__inst_mult_17_76  = SUM(( !Xd_0__inst_mult_17_20_q  $ (((!Xd_0__inst_mult_17_19_q ) # (!Xd_0__inst_mult_17_18_q ))) ) + ( Xd_0__inst_mult_17_74  ) + ( Xd_0__inst_mult_17_73  ))
// Xd_0__inst_mult_17_77  = CARRY(( !Xd_0__inst_mult_17_20_q  $ (((!Xd_0__inst_mult_17_19_q ) # (!Xd_0__inst_mult_17_18_q ))) ) + ( Xd_0__inst_mult_17_74  ) + ( Xd_0__inst_mult_17_73  ))
// Xd_0__inst_mult_17_78  = SHARE((Xd_0__inst_mult_17_19_q  & (Xd_0__inst_mult_17_18_q  & Xd_0__inst_mult_17_20_q )))

	.dataa(!Xd_0__inst_mult_17_19_q ),
	.datab(!Xd_0__inst_mult_17_18_q ),
	.datac(!Xd_0__inst_mult_17_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_73 ),
	.sharein(Xd_0__inst_mult_17_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_76 ),
	.cout(Xd_0__inst_mult_17_77 ),
	.shareout(Xd_0__inst_mult_17_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_26 (
// Equation(s):
// Xd_0__inst_mult_14_76  = SUM(( !Xd_0__inst_mult_14_20_q  $ (((!Xd_0__inst_mult_14_19_q ) # (!Xd_0__inst_mult_14_18_q ))) ) + ( Xd_0__inst_mult_14_74  ) + ( Xd_0__inst_mult_14_73  ))
// Xd_0__inst_mult_14_77  = CARRY(( !Xd_0__inst_mult_14_20_q  $ (((!Xd_0__inst_mult_14_19_q ) # (!Xd_0__inst_mult_14_18_q ))) ) + ( Xd_0__inst_mult_14_74  ) + ( Xd_0__inst_mult_14_73  ))
// Xd_0__inst_mult_14_78  = SHARE((Xd_0__inst_mult_14_19_q  & (Xd_0__inst_mult_14_18_q  & Xd_0__inst_mult_14_20_q )))

	.dataa(!Xd_0__inst_mult_14_19_q ),
	.datab(!Xd_0__inst_mult_14_18_q ),
	.datac(!Xd_0__inst_mult_14_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_73 ),
	.sharein(Xd_0__inst_mult_14_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_76 ),
	.cout(Xd_0__inst_mult_14_77 ),
	.shareout(Xd_0__inst_mult_14_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_26 (
// Equation(s):
// Xd_0__inst_mult_15_76  = SUM(( !Xd_0__inst_mult_15_20_q  $ (((!Xd_0__inst_mult_15_19_q ) # (!Xd_0__inst_mult_15_18_q ))) ) + ( Xd_0__inst_mult_15_74  ) + ( Xd_0__inst_mult_15_73  ))
// Xd_0__inst_mult_15_77  = CARRY(( !Xd_0__inst_mult_15_20_q  $ (((!Xd_0__inst_mult_15_19_q ) # (!Xd_0__inst_mult_15_18_q ))) ) + ( Xd_0__inst_mult_15_74  ) + ( Xd_0__inst_mult_15_73  ))
// Xd_0__inst_mult_15_78  = SHARE((Xd_0__inst_mult_15_19_q  & (Xd_0__inst_mult_15_18_q  & Xd_0__inst_mult_15_20_q )))

	.dataa(!Xd_0__inst_mult_15_19_q ),
	.datab(!Xd_0__inst_mult_15_18_q ),
	.datac(!Xd_0__inst_mult_15_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_73 ),
	.sharein(Xd_0__inst_mult_15_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_76 ),
	.cout(Xd_0__inst_mult_15_77 ),
	.shareout(Xd_0__inst_mult_15_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_26 (
// Equation(s):
// Xd_0__inst_mult_12_76  = SUM(( !Xd_0__inst_mult_12_20_q  $ (((!Xd_0__inst_mult_12_19_q ) # (!Xd_0__inst_mult_12_18_q ))) ) + ( Xd_0__inst_mult_12_74  ) + ( Xd_0__inst_mult_12_73  ))
// Xd_0__inst_mult_12_77  = CARRY(( !Xd_0__inst_mult_12_20_q  $ (((!Xd_0__inst_mult_12_19_q ) # (!Xd_0__inst_mult_12_18_q ))) ) + ( Xd_0__inst_mult_12_74  ) + ( Xd_0__inst_mult_12_73  ))
// Xd_0__inst_mult_12_78  = SHARE((Xd_0__inst_mult_12_19_q  & (Xd_0__inst_mult_12_18_q  & Xd_0__inst_mult_12_20_q )))

	.dataa(!Xd_0__inst_mult_12_19_q ),
	.datab(!Xd_0__inst_mult_12_18_q ),
	.datac(!Xd_0__inst_mult_12_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_73 ),
	.sharein(Xd_0__inst_mult_12_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_76 ),
	.cout(Xd_0__inst_mult_12_77 ),
	.shareout(Xd_0__inst_mult_12_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_26 (
// Equation(s):
// Xd_0__inst_mult_13_76  = SUM(( !Xd_0__inst_mult_13_20_q  $ (((!Xd_0__inst_mult_13_19_q ) # (!Xd_0__inst_mult_13_18_q ))) ) + ( Xd_0__inst_mult_13_74  ) + ( Xd_0__inst_mult_13_73  ))
// Xd_0__inst_mult_13_77  = CARRY(( !Xd_0__inst_mult_13_20_q  $ (((!Xd_0__inst_mult_13_19_q ) # (!Xd_0__inst_mult_13_18_q ))) ) + ( Xd_0__inst_mult_13_74  ) + ( Xd_0__inst_mult_13_73  ))
// Xd_0__inst_mult_13_78  = SHARE((Xd_0__inst_mult_13_19_q  & (Xd_0__inst_mult_13_18_q  & Xd_0__inst_mult_13_20_q )))

	.dataa(!Xd_0__inst_mult_13_19_q ),
	.datab(!Xd_0__inst_mult_13_18_q ),
	.datac(!Xd_0__inst_mult_13_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_73 ),
	.sharein(Xd_0__inst_mult_13_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_76 ),
	.cout(Xd_0__inst_mult_13_77 ),
	.shareout(Xd_0__inst_mult_13_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_26 (
// Equation(s):
// Xd_0__inst_mult_10_76  = SUM(( !Xd_0__inst_mult_10_20_q  $ (((!Xd_0__inst_mult_10_19_q ) # (!Xd_0__inst_mult_10_18_q ))) ) + ( Xd_0__inst_mult_10_74  ) + ( Xd_0__inst_mult_10_73  ))
// Xd_0__inst_mult_10_77  = CARRY(( !Xd_0__inst_mult_10_20_q  $ (((!Xd_0__inst_mult_10_19_q ) # (!Xd_0__inst_mult_10_18_q ))) ) + ( Xd_0__inst_mult_10_74  ) + ( Xd_0__inst_mult_10_73  ))
// Xd_0__inst_mult_10_78  = SHARE((Xd_0__inst_mult_10_19_q  & (Xd_0__inst_mult_10_18_q  & Xd_0__inst_mult_10_20_q )))

	.dataa(!Xd_0__inst_mult_10_19_q ),
	.datab(!Xd_0__inst_mult_10_18_q ),
	.datac(!Xd_0__inst_mult_10_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_73 ),
	.sharein(Xd_0__inst_mult_10_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_76 ),
	.cout(Xd_0__inst_mult_10_77 ),
	.shareout(Xd_0__inst_mult_10_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_26 (
// Equation(s):
// Xd_0__inst_mult_11_76  = SUM(( !Xd_0__inst_mult_11_20_q  $ (((!Xd_0__inst_mult_11_19_q ) # (!Xd_0__inst_mult_11_18_q ))) ) + ( Xd_0__inst_mult_11_74  ) + ( Xd_0__inst_mult_11_73  ))
// Xd_0__inst_mult_11_77  = CARRY(( !Xd_0__inst_mult_11_20_q  $ (((!Xd_0__inst_mult_11_19_q ) # (!Xd_0__inst_mult_11_18_q ))) ) + ( Xd_0__inst_mult_11_74  ) + ( Xd_0__inst_mult_11_73  ))
// Xd_0__inst_mult_11_78  = SHARE((Xd_0__inst_mult_11_19_q  & (Xd_0__inst_mult_11_18_q  & Xd_0__inst_mult_11_20_q )))

	.dataa(!Xd_0__inst_mult_11_19_q ),
	.datab(!Xd_0__inst_mult_11_18_q ),
	.datac(!Xd_0__inst_mult_11_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_73 ),
	.sharein(Xd_0__inst_mult_11_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_76 ),
	.cout(Xd_0__inst_mult_11_77 ),
	.shareout(Xd_0__inst_mult_11_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_26 (
// Equation(s):
// Xd_0__inst_mult_8_76  = SUM(( !Xd_0__inst_mult_8_20_q  $ (((!Xd_0__inst_mult_8_19_q ) # (!Xd_0__inst_mult_8_18_q ))) ) + ( Xd_0__inst_mult_8_74  ) + ( Xd_0__inst_mult_8_73  ))
// Xd_0__inst_mult_8_77  = CARRY(( !Xd_0__inst_mult_8_20_q  $ (((!Xd_0__inst_mult_8_19_q ) # (!Xd_0__inst_mult_8_18_q ))) ) + ( Xd_0__inst_mult_8_74  ) + ( Xd_0__inst_mult_8_73  ))
// Xd_0__inst_mult_8_78  = SHARE((Xd_0__inst_mult_8_19_q  & (Xd_0__inst_mult_8_18_q  & Xd_0__inst_mult_8_20_q )))

	.dataa(!Xd_0__inst_mult_8_19_q ),
	.datab(!Xd_0__inst_mult_8_18_q ),
	.datac(!Xd_0__inst_mult_8_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_73 ),
	.sharein(Xd_0__inst_mult_8_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_76 ),
	.cout(Xd_0__inst_mult_8_77 ),
	.shareout(Xd_0__inst_mult_8_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_26 (
// Equation(s):
// Xd_0__inst_mult_9_76  = SUM(( !Xd_0__inst_mult_9_20_q  $ (((!Xd_0__inst_mult_9_19_q ) # (!Xd_0__inst_mult_9_18_q ))) ) + ( Xd_0__inst_mult_9_74  ) + ( Xd_0__inst_mult_9_73  ))
// Xd_0__inst_mult_9_77  = CARRY(( !Xd_0__inst_mult_9_20_q  $ (((!Xd_0__inst_mult_9_19_q ) # (!Xd_0__inst_mult_9_18_q ))) ) + ( Xd_0__inst_mult_9_74  ) + ( Xd_0__inst_mult_9_73  ))
// Xd_0__inst_mult_9_78  = SHARE((Xd_0__inst_mult_9_19_q  & (Xd_0__inst_mult_9_18_q  & Xd_0__inst_mult_9_20_q )))

	.dataa(!Xd_0__inst_mult_9_19_q ),
	.datab(!Xd_0__inst_mult_9_18_q ),
	.datac(!Xd_0__inst_mult_9_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_73 ),
	.sharein(Xd_0__inst_mult_9_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_76 ),
	.cout(Xd_0__inst_mult_9_77 ),
	.shareout(Xd_0__inst_mult_9_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_26 (
// Equation(s):
// Xd_0__inst_mult_6_76  = SUM(( !Xd_0__inst_mult_6_20_q  $ (((!Xd_0__inst_mult_6_19_q ) # (!Xd_0__inst_mult_6_18_q ))) ) + ( Xd_0__inst_mult_6_74  ) + ( Xd_0__inst_mult_6_73  ))
// Xd_0__inst_mult_6_77  = CARRY(( !Xd_0__inst_mult_6_20_q  $ (((!Xd_0__inst_mult_6_19_q ) # (!Xd_0__inst_mult_6_18_q ))) ) + ( Xd_0__inst_mult_6_74  ) + ( Xd_0__inst_mult_6_73  ))
// Xd_0__inst_mult_6_78  = SHARE((Xd_0__inst_mult_6_19_q  & (Xd_0__inst_mult_6_18_q  & Xd_0__inst_mult_6_20_q )))

	.dataa(!Xd_0__inst_mult_6_19_q ),
	.datab(!Xd_0__inst_mult_6_18_q ),
	.datac(!Xd_0__inst_mult_6_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_73 ),
	.sharein(Xd_0__inst_mult_6_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_76 ),
	.cout(Xd_0__inst_mult_6_77 ),
	.shareout(Xd_0__inst_mult_6_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_26 (
// Equation(s):
// Xd_0__inst_mult_7_76  = SUM(( !Xd_0__inst_mult_7_20_q  $ (((!Xd_0__inst_mult_7_19_q ) # (!Xd_0__inst_mult_7_18_q ))) ) + ( Xd_0__inst_mult_7_74  ) + ( Xd_0__inst_mult_7_73  ))
// Xd_0__inst_mult_7_77  = CARRY(( !Xd_0__inst_mult_7_20_q  $ (((!Xd_0__inst_mult_7_19_q ) # (!Xd_0__inst_mult_7_18_q ))) ) + ( Xd_0__inst_mult_7_74  ) + ( Xd_0__inst_mult_7_73  ))
// Xd_0__inst_mult_7_78  = SHARE((Xd_0__inst_mult_7_19_q  & (Xd_0__inst_mult_7_18_q  & Xd_0__inst_mult_7_20_q )))

	.dataa(!Xd_0__inst_mult_7_19_q ),
	.datab(!Xd_0__inst_mult_7_18_q ),
	.datac(!Xd_0__inst_mult_7_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_73 ),
	.sharein(Xd_0__inst_mult_7_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_76 ),
	.cout(Xd_0__inst_mult_7_77 ),
	.shareout(Xd_0__inst_mult_7_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_26 (
// Equation(s):
// Xd_0__inst_mult_4_76  = SUM(( !Xd_0__inst_mult_4_20_q  $ (((!Xd_0__inst_mult_4_19_q ) # (!Xd_0__inst_mult_4_18_q ))) ) + ( Xd_0__inst_mult_4_74  ) + ( Xd_0__inst_mult_4_73  ))
// Xd_0__inst_mult_4_77  = CARRY(( !Xd_0__inst_mult_4_20_q  $ (((!Xd_0__inst_mult_4_19_q ) # (!Xd_0__inst_mult_4_18_q ))) ) + ( Xd_0__inst_mult_4_74  ) + ( Xd_0__inst_mult_4_73  ))
// Xd_0__inst_mult_4_78  = SHARE((Xd_0__inst_mult_4_19_q  & (Xd_0__inst_mult_4_18_q  & Xd_0__inst_mult_4_20_q )))

	.dataa(!Xd_0__inst_mult_4_19_q ),
	.datab(!Xd_0__inst_mult_4_18_q ),
	.datac(!Xd_0__inst_mult_4_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_73 ),
	.sharein(Xd_0__inst_mult_4_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_76 ),
	.cout(Xd_0__inst_mult_4_77 ),
	.shareout(Xd_0__inst_mult_4_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_26 (
// Equation(s):
// Xd_0__inst_mult_5_76  = SUM(( !Xd_0__inst_mult_5_20_q  $ (((!Xd_0__inst_mult_5_19_q ) # (!Xd_0__inst_mult_5_18_q ))) ) + ( Xd_0__inst_mult_5_74  ) + ( Xd_0__inst_mult_5_73  ))
// Xd_0__inst_mult_5_77  = CARRY(( !Xd_0__inst_mult_5_20_q  $ (((!Xd_0__inst_mult_5_19_q ) # (!Xd_0__inst_mult_5_18_q ))) ) + ( Xd_0__inst_mult_5_74  ) + ( Xd_0__inst_mult_5_73  ))
// Xd_0__inst_mult_5_78  = SHARE((Xd_0__inst_mult_5_19_q  & (Xd_0__inst_mult_5_18_q  & Xd_0__inst_mult_5_20_q )))

	.dataa(!Xd_0__inst_mult_5_19_q ),
	.datab(!Xd_0__inst_mult_5_18_q ),
	.datac(!Xd_0__inst_mult_5_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_73 ),
	.sharein(Xd_0__inst_mult_5_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_76 ),
	.cout(Xd_0__inst_mult_5_77 ),
	.shareout(Xd_0__inst_mult_5_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_26 (
// Equation(s):
// Xd_0__inst_mult_2_76  = SUM(( !Xd_0__inst_mult_2_20_q  $ (((!Xd_0__inst_mult_2_19_q ) # (!Xd_0__inst_mult_2_18_q ))) ) + ( Xd_0__inst_mult_2_74  ) + ( Xd_0__inst_mult_2_73  ))
// Xd_0__inst_mult_2_77  = CARRY(( !Xd_0__inst_mult_2_20_q  $ (((!Xd_0__inst_mult_2_19_q ) # (!Xd_0__inst_mult_2_18_q ))) ) + ( Xd_0__inst_mult_2_74  ) + ( Xd_0__inst_mult_2_73  ))
// Xd_0__inst_mult_2_78  = SHARE((Xd_0__inst_mult_2_19_q  & (Xd_0__inst_mult_2_18_q  & Xd_0__inst_mult_2_20_q )))

	.dataa(!Xd_0__inst_mult_2_19_q ),
	.datab(!Xd_0__inst_mult_2_18_q ),
	.datac(!Xd_0__inst_mult_2_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_73 ),
	.sharein(Xd_0__inst_mult_2_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_76 ),
	.cout(Xd_0__inst_mult_2_77 ),
	.shareout(Xd_0__inst_mult_2_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_26 (
// Equation(s):
// Xd_0__inst_mult_3_76  = SUM(( !Xd_0__inst_mult_3_20_q  $ (((!Xd_0__inst_mult_3_19_q ) # (!Xd_0__inst_mult_3_18_q ))) ) + ( Xd_0__inst_mult_3_74  ) + ( Xd_0__inst_mult_3_73  ))
// Xd_0__inst_mult_3_77  = CARRY(( !Xd_0__inst_mult_3_20_q  $ (((!Xd_0__inst_mult_3_19_q ) # (!Xd_0__inst_mult_3_18_q ))) ) + ( Xd_0__inst_mult_3_74  ) + ( Xd_0__inst_mult_3_73  ))
// Xd_0__inst_mult_3_78  = SHARE((Xd_0__inst_mult_3_19_q  & (Xd_0__inst_mult_3_18_q  & Xd_0__inst_mult_3_20_q )))

	.dataa(!Xd_0__inst_mult_3_19_q ),
	.datab(!Xd_0__inst_mult_3_18_q ),
	.datac(!Xd_0__inst_mult_3_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_73 ),
	.sharein(Xd_0__inst_mult_3_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_76 ),
	.cout(Xd_0__inst_mult_3_77 ),
	.shareout(Xd_0__inst_mult_3_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_26 (
// Equation(s):
// Xd_0__inst_mult_0_76  = SUM(( !Xd_0__inst_mult_0_20_q  $ (((!Xd_0__inst_mult_0_19_q ) # (!Xd_0__inst_mult_0_18_q ))) ) + ( Xd_0__inst_mult_0_74  ) + ( Xd_0__inst_mult_0_73  ))
// Xd_0__inst_mult_0_77  = CARRY(( !Xd_0__inst_mult_0_20_q  $ (((!Xd_0__inst_mult_0_19_q ) # (!Xd_0__inst_mult_0_18_q ))) ) + ( Xd_0__inst_mult_0_74  ) + ( Xd_0__inst_mult_0_73  ))
// Xd_0__inst_mult_0_78  = SHARE((Xd_0__inst_mult_0_19_q  & (Xd_0__inst_mult_0_18_q  & Xd_0__inst_mult_0_20_q )))

	.dataa(!Xd_0__inst_mult_0_19_q ),
	.datab(!Xd_0__inst_mult_0_18_q ),
	.datac(!Xd_0__inst_mult_0_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_73 ),
	.sharein(Xd_0__inst_mult_0_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_76 ),
	.cout(Xd_0__inst_mult_0_77 ),
	.shareout(Xd_0__inst_mult_0_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_26 (
// Equation(s):
// Xd_0__inst_mult_1_76  = SUM(( !Xd_0__inst_mult_1_20_q  $ (((!Xd_0__inst_mult_1_19_q ) # (!Xd_0__inst_mult_1_18_q ))) ) + ( Xd_0__inst_mult_1_74  ) + ( Xd_0__inst_mult_1_73  ))
// Xd_0__inst_mult_1_77  = CARRY(( !Xd_0__inst_mult_1_20_q  $ (((!Xd_0__inst_mult_1_19_q ) # (!Xd_0__inst_mult_1_18_q ))) ) + ( Xd_0__inst_mult_1_74  ) + ( Xd_0__inst_mult_1_73  ))
// Xd_0__inst_mult_1_78  = SHARE((Xd_0__inst_mult_1_19_q  & (Xd_0__inst_mult_1_18_q  & Xd_0__inst_mult_1_20_q )))

	.dataa(!Xd_0__inst_mult_1_19_q ),
	.datab(!Xd_0__inst_mult_1_18_q ),
	.datac(!Xd_0__inst_mult_1_20_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_73 ),
	.sharein(Xd_0__inst_mult_1_74 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_76 ),
	.cout(Xd_0__inst_mult_1_77 ),
	.shareout(Xd_0__inst_mult_1_78 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_27 (
// Equation(s):
// Xd_0__inst_mult_28_80  = SUM(( GND ) + ( Xd_0__inst_mult_28_78  ) + ( Xd_0__inst_mult_28_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_77 ),
	.sharein(Xd_0__inst_mult_28_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_27 (
// Equation(s):
// Xd_0__inst_mult_29_80  = SUM(( GND ) + ( Xd_0__inst_mult_29_78  ) + ( Xd_0__inst_mult_29_77  ))
// Xd_0__inst_mult_29_81  = CARRY(( GND ) + ( Xd_0__inst_mult_29_78  ) + ( Xd_0__inst_mult_29_77  ))
// Xd_0__inst_mult_29_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_77 ),
	.sharein(Xd_0__inst_mult_29_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_80 ),
	.cout(Xd_0__inst_mult_29_81 ),
	.shareout(Xd_0__inst_mult_29_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_27 (
// Equation(s):
// Xd_0__inst_mult_26_80  = SUM(( GND ) + ( Xd_0__inst_mult_26_78  ) + ( Xd_0__inst_mult_26_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_77 ),
	.sharein(Xd_0__inst_mult_26_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_27 (
// Equation(s):
// Xd_0__inst_mult_27_80  = SUM(( GND ) + ( Xd_0__inst_mult_27_78  ) + ( Xd_0__inst_mult_27_77  ))
// Xd_0__inst_mult_27_81  = CARRY(( GND ) + ( Xd_0__inst_mult_27_78  ) + ( Xd_0__inst_mult_27_77  ))
// Xd_0__inst_mult_27_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_77 ),
	.sharein(Xd_0__inst_mult_27_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_80 ),
	.cout(Xd_0__inst_mult_27_81 ),
	.shareout(Xd_0__inst_mult_27_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_27 (
// Equation(s):
// Xd_0__inst_mult_24_80  = SUM(( GND ) + ( Xd_0__inst_mult_24_78  ) + ( Xd_0__inst_mult_24_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_77 ),
	.sharein(Xd_0__inst_mult_24_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_27 (
// Equation(s):
// Xd_0__inst_mult_25_80  = SUM(( GND ) + ( Xd_0__inst_mult_25_78  ) + ( Xd_0__inst_mult_25_77  ))
// Xd_0__inst_mult_25_81  = CARRY(( GND ) + ( Xd_0__inst_mult_25_78  ) + ( Xd_0__inst_mult_25_77  ))
// Xd_0__inst_mult_25_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_77 ),
	.sharein(Xd_0__inst_mult_25_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_80 ),
	.cout(Xd_0__inst_mult_25_81 ),
	.shareout(Xd_0__inst_mult_25_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_27 (
// Equation(s):
// Xd_0__inst_mult_22_80  = SUM(( GND ) + ( Xd_0__inst_mult_22_78  ) + ( Xd_0__inst_mult_22_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_77 ),
	.sharein(Xd_0__inst_mult_22_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_27 (
// Equation(s):
// Xd_0__inst_mult_23_80  = SUM(( GND ) + ( Xd_0__inst_mult_23_78  ) + ( Xd_0__inst_mult_23_77  ))
// Xd_0__inst_mult_23_81  = CARRY(( GND ) + ( Xd_0__inst_mult_23_78  ) + ( Xd_0__inst_mult_23_77  ))
// Xd_0__inst_mult_23_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_77 ),
	.sharein(Xd_0__inst_mult_23_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_80 ),
	.cout(Xd_0__inst_mult_23_81 ),
	.shareout(Xd_0__inst_mult_23_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_27 (
// Equation(s):
// Xd_0__inst_mult_20_80  = SUM(( GND ) + ( Xd_0__inst_mult_20_78  ) + ( Xd_0__inst_mult_20_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_77 ),
	.sharein(Xd_0__inst_mult_20_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_27 (
// Equation(s):
// Xd_0__inst_mult_21_80  = SUM(( GND ) + ( Xd_0__inst_mult_21_78  ) + ( Xd_0__inst_mult_21_77  ))
// Xd_0__inst_mult_21_81  = CARRY(( GND ) + ( Xd_0__inst_mult_21_78  ) + ( Xd_0__inst_mult_21_77  ))
// Xd_0__inst_mult_21_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_77 ),
	.sharein(Xd_0__inst_mult_21_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_80 ),
	.cout(Xd_0__inst_mult_21_81 ),
	.shareout(Xd_0__inst_mult_21_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_27 (
// Equation(s):
// Xd_0__inst_mult_18_80  = SUM(( GND ) + ( Xd_0__inst_mult_18_78  ) + ( Xd_0__inst_mult_18_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_77 ),
	.sharein(Xd_0__inst_mult_18_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_27 (
// Equation(s):
// Xd_0__inst_mult_19_80  = SUM(( GND ) + ( Xd_0__inst_mult_19_78  ) + ( Xd_0__inst_mult_19_77  ))
// Xd_0__inst_mult_19_81  = CARRY(( GND ) + ( Xd_0__inst_mult_19_78  ) + ( Xd_0__inst_mult_19_77  ))
// Xd_0__inst_mult_19_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_77 ),
	.sharein(Xd_0__inst_mult_19_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_80 ),
	.cout(Xd_0__inst_mult_19_81 ),
	.shareout(Xd_0__inst_mult_19_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_27 (
// Equation(s):
// Xd_0__inst_mult_16_80  = SUM(( GND ) + ( Xd_0__inst_mult_16_78  ) + ( Xd_0__inst_mult_16_77  ))
// Xd_0__inst_mult_16_81  = CARRY(( GND ) + ( Xd_0__inst_mult_16_78  ) + ( Xd_0__inst_mult_16_77  ))
// Xd_0__inst_mult_16_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_77 ),
	.sharein(Xd_0__inst_mult_16_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_80 ),
	.cout(Xd_0__inst_mult_16_81 ),
	.shareout(Xd_0__inst_mult_16_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_27 (
// Equation(s):
// Xd_0__inst_mult_17_80  = SUM(( GND ) + ( Xd_0__inst_mult_17_78  ) + ( Xd_0__inst_mult_17_77  ))
// Xd_0__inst_mult_17_81  = CARRY(( GND ) + ( Xd_0__inst_mult_17_78  ) + ( Xd_0__inst_mult_17_77  ))
// Xd_0__inst_mult_17_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_77 ),
	.sharein(Xd_0__inst_mult_17_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_80 ),
	.cout(Xd_0__inst_mult_17_81 ),
	.shareout(Xd_0__inst_mult_17_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_27 (
// Equation(s):
// Xd_0__inst_mult_14_80  = SUM(( GND ) + ( Xd_0__inst_mult_14_78  ) + ( Xd_0__inst_mult_14_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_77 ),
	.sharein(Xd_0__inst_mult_14_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_27 (
// Equation(s):
// Xd_0__inst_mult_15_80  = SUM(( GND ) + ( Xd_0__inst_mult_15_78  ) + ( Xd_0__inst_mult_15_77  ))
// Xd_0__inst_mult_15_81  = CARRY(( GND ) + ( Xd_0__inst_mult_15_78  ) + ( Xd_0__inst_mult_15_77  ))
// Xd_0__inst_mult_15_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_77 ),
	.sharein(Xd_0__inst_mult_15_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_80 ),
	.cout(Xd_0__inst_mult_15_81 ),
	.shareout(Xd_0__inst_mult_15_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_27 (
// Equation(s):
// Xd_0__inst_mult_12_80  = SUM(( GND ) + ( Xd_0__inst_mult_12_78  ) + ( Xd_0__inst_mult_12_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_77 ),
	.sharein(Xd_0__inst_mult_12_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_27 (
// Equation(s):
// Xd_0__inst_mult_13_80  = SUM(( GND ) + ( Xd_0__inst_mult_13_78  ) + ( Xd_0__inst_mult_13_77  ))
// Xd_0__inst_mult_13_81  = CARRY(( GND ) + ( Xd_0__inst_mult_13_78  ) + ( Xd_0__inst_mult_13_77  ))
// Xd_0__inst_mult_13_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_77 ),
	.sharein(Xd_0__inst_mult_13_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_80 ),
	.cout(Xd_0__inst_mult_13_81 ),
	.shareout(Xd_0__inst_mult_13_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_27 (
// Equation(s):
// Xd_0__inst_mult_10_80  = SUM(( GND ) + ( Xd_0__inst_mult_10_78  ) + ( Xd_0__inst_mult_10_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_77 ),
	.sharein(Xd_0__inst_mult_10_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_27 (
// Equation(s):
// Xd_0__inst_mult_11_80  = SUM(( GND ) + ( Xd_0__inst_mult_11_78  ) + ( Xd_0__inst_mult_11_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_77 ),
	.sharein(Xd_0__inst_mult_11_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_27 (
// Equation(s):
// Xd_0__inst_mult_8_80  = SUM(( GND ) + ( Xd_0__inst_mult_8_78  ) + ( Xd_0__inst_mult_8_77  ))
// Xd_0__inst_mult_8_81  = CARRY(( GND ) + ( Xd_0__inst_mult_8_78  ) + ( Xd_0__inst_mult_8_77  ))
// Xd_0__inst_mult_8_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_77 ),
	.sharein(Xd_0__inst_mult_8_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_80 ),
	.cout(Xd_0__inst_mult_8_81 ),
	.shareout(Xd_0__inst_mult_8_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_27 (
// Equation(s):
// Xd_0__inst_mult_9_80  = SUM(( GND ) + ( Xd_0__inst_mult_9_78  ) + ( Xd_0__inst_mult_9_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_77 ),
	.sharein(Xd_0__inst_mult_9_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_27 (
// Equation(s):
// Xd_0__inst_mult_6_80  = SUM(( GND ) + ( Xd_0__inst_mult_6_78  ) + ( Xd_0__inst_mult_6_77  ))
// Xd_0__inst_mult_6_81  = CARRY(( GND ) + ( Xd_0__inst_mult_6_78  ) + ( Xd_0__inst_mult_6_77  ))
// Xd_0__inst_mult_6_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_77 ),
	.sharein(Xd_0__inst_mult_6_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_80 ),
	.cout(Xd_0__inst_mult_6_81 ),
	.shareout(Xd_0__inst_mult_6_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_27 (
// Equation(s):
// Xd_0__inst_mult_7_80  = SUM(( GND ) + ( Xd_0__inst_mult_7_78  ) + ( Xd_0__inst_mult_7_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_77 ),
	.sharein(Xd_0__inst_mult_7_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_27 (
// Equation(s):
// Xd_0__inst_mult_4_80  = SUM(( GND ) + ( Xd_0__inst_mult_4_78  ) + ( Xd_0__inst_mult_4_77  ))
// Xd_0__inst_mult_4_81  = CARRY(( GND ) + ( Xd_0__inst_mult_4_78  ) + ( Xd_0__inst_mult_4_77  ))
// Xd_0__inst_mult_4_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_77 ),
	.sharein(Xd_0__inst_mult_4_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_80 ),
	.cout(Xd_0__inst_mult_4_81 ),
	.shareout(Xd_0__inst_mult_4_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_27 (
// Equation(s):
// Xd_0__inst_mult_5_80  = SUM(( GND ) + ( Xd_0__inst_mult_5_78  ) + ( Xd_0__inst_mult_5_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_77 ),
	.sharein(Xd_0__inst_mult_5_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_27 (
// Equation(s):
// Xd_0__inst_mult_2_80  = SUM(( GND ) + ( Xd_0__inst_mult_2_78  ) + ( Xd_0__inst_mult_2_77  ))
// Xd_0__inst_mult_2_81  = CARRY(( GND ) + ( Xd_0__inst_mult_2_78  ) + ( Xd_0__inst_mult_2_77  ))
// Xd_0__inst_mult_2_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_77 ),
	.sharein(Xd_0__inst_mult_2_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_80 ),
	.cout(Xd_0__inst_mult_2_81 ),
	.shareout(Xd_0__inst_mult_2_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_27 (
// Equation(s):
// Xd_0__inst_mult_3_80  = SUM(( GND ) + ( Xd_0__inst_mult_3_78  ) + ( Xd_0__inst_mult_3_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_77 ),
	.sharein(Xd_0__inst_mult_3_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_27 (
// Equation(s):
// Xd_0__inst_mult_0_80  = SUM(( GND ) + ( Xd_0__inst_mult_0_78  ) + ( Xd_0__inst_mult_0_77  ))
// Xd_0__inst_mult_0_81  = CARRY(( GND ) + ( Xd_0__inst_mult_0_78  ) + ( Xd_0__inst_mult_0_77  ))
// Xd_0__inst_mult_0_82  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_77 ),
	.sharein(Xd_0__inst_mult_0_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_80 ),
	.cout(Xd_0__inst_mult_0_81 ),
	.shareout(Xd_0__inst_mult_0_82 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_27 (
// Equation(s):
// Xd_0__inst_mult_1_80  = SUM(( GND ) + ( Xd_0__inst_mult_1_78  ) + ( Xd_0__inst_mult_1_77  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_77 ),
	.sharein(Xd_0__inst_mult_1_78 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_80 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_28 (
// Equation(s):
// Xd_0__inst_mult_28_84  = SUM(( (din_a[196] & din_b[196]) ) + ( Xd_0__inst_mult_14_102  ) + ( Xd_0__inst_mult_14_101  ))
// Xd_0__inst_mult_28_85  = CARRY(( (din_a[196] & din_b[196]) ) + ( Xd_0__inst_mult_14_102  ) + ( Xd_0__inst_mult_14_101  ))
// Xd_0__inst_mult_28_86  = SHARE((din_a[196] & din_b[197]))

	.dataa(!din_a[196]),
	.datab(!din_b[196]),
	.datac(!din_b[197]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_101 ),
	.sharein(Xd_0__inst_mult_14_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_84 ),
	.cout(Xd_0__inst_mult_28_85 ),
	.shareout(Xd_0__inst_mult_28_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_28 (
// Equation(s):
// Xd_0__inst_mult_29_84  = SUM(( (din_a[203] & din_b[203]) ) + ( Xd_0__inst_mult_19_102  ) + ( Xd_0__inst_mult_19_101  ))
// Xd_0__inst_mult_29_85  = CARRY(( (din_a[203] & din_b[203]) ) + ( Xd_0__inst_mult_19_102  ) + ( Xd_0__inst_mult_19_101  ))
// Xd_0__inst_mult_29_86  = SHARE((din_a[203] & din_b[204]))

	.dataa(!din_a[203]),
	.datab(!din_b[203]),
	.datac(!din_b[204]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_101 ),
	.sharein(Xd_0__inst_mult_19_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_84 ),
	.cout(Xd_0__inst_mult_29_85 ),
	.shareout(Xd_0__inst_mult_29_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_28 (
// Equation(s):
// Xd_0__inst_mult_26_84  = SUM(( (din_a[182] & din_b[182]) ) + ( Xd_0__inst_mult_21_102  ) + ( Xd_0__inst_mult_21_101  ))
// Xd_0__inst_mult_26_85  = CARRY(( (din_a[182] & din_b[182]) ) + ( Xd_0__inst_mult_21_102  ) + ( Xd_0__inst_mult_21_101  ))
// Xd_0__inst_mult_26_86  = SHARE((din_a[182] & din_b[183]))

	.dataa(!din_a[182]),
	.datab(!din_b[182]),
	.datac(!din_b[183]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_101 ),
	.sharein(Xd_0__inst_mult_21_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_84 ),
	.cout(Xd_0__inst_mult_26_85 ),
	.shareout(Xd_0__inst_mult_26_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_28 (
// Equation(s):
// Xd_0__inst_mult_27_84  = SUM(( (din_a[189] & din_b[189]) ) + ( Xd_0__inst_mult_18_102  ) + ( Xd_0__inst_mult_18_101  ))
// Xd_0__inst_mult_27_85  = CARRY(( (din_a[189] & din_b[189]) ) + ( Xd_0__inst_mult_18_102  ) + ( Xd_0__inst_mult_18_101  ))
// Xd_0__inst_mult_27_86  = SHARE((din_a[189] & din_b[190]))

	.dataa(!din_a[189]),
	.datab(!din_b[189]),
	.datac(!din_b[190]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_101 ),
	.sharein(Xd_0__inst_mult_18_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_84 ),
	.cout(Xd_0__inst_mult_27_85 ),
	.shareout(Xd_0__inst_mult_27_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_28 (
// Equation(s):
// Xd_0__inst_mult_24_84  = SUM(( (din_a[168] & din_b[168]) ) + ( Xd_0__inst_mult_17_102  ) + ( Xd_0__inst_mult_17_101  ))
// Xd_0__inst_mult_24_85  = CARRY(( (din_a[168] & din_b[168]) ) + ( Xd_0__inst_mult_17_102  ) + ( Xd_0__inst_mult_17_101  ))
// Xd_0__inst_mult_24_86  = SHARE((din_a[168] & din_b[169]))

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(!din_b[169]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_101 ),
	.sharein(Xd_0__inst_mult_17_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_84 ),
	.cout(Xd_0__inst_mult_24_85 ),
	.shareout(Xd_0__inst_mult_24_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_28 (
// Equation(s):
// Xd_0__inst_mult_25_84  = SUM(( (din_a[175] & din_b[175]) ) + ( Xd_0__inst_mult_16_102  ) + ( Xd_0__inst_mult_16_101  ))
// Xd_0__inst_mult_25_85  = CARRY(( (din_a[175] & din_b[175]) ) + ( Xd_0__inst_mult_16_102  ) + ( Xd_0__inst_mult_16_101  ))
// Xd_0__inst_mult_25_86  = SHARE((din_a[175] & din_b[176]))

	.dataa(!din_a[175]),
	.datab(!din_b[175]),
	.datac(!din_b[176]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_101 ),
	.sharein(Xd_0__inst_mult_16_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_84 ),
	.cout(Xd_0__inst_mult_25_85 ),
	.shareout(Xd_0__inst_mult_25_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_28 (
// Equation(s):
// Xd_0__inst_mult_22_84  = SUM(( (din_a[154] & din_b[154]) ) + ( Xd_0__inst_mult_20_102  ) + ( Xd_0__inst_mult_20_101  ))
// Xd_0__inst_mult_22_85  = CARRY(( (din_a[154] & din_b[154]) ) + ( Xd_0__inst_mult_20_102  ) + ( Xd_0__inst_mult_20_101  ))
// Xd_0__inst_mult_22_86  = SHARE((din_a[154] & din_b[155]))

	.dataa(!din_a[154]),
	.datab(!din_b[154]),
	.datac(!din_b[155]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_101 ),
	.sharein(Xd_0__inst_mult_20_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_84 ),
	.cout(Xd_0__inst_mult_22_85 ),
	.shareout(Xd_0__inst_mult_22_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_28 (
// Equation(s):
// Xd_0__inst_mult_23_84  = SUM(( (din_a[161] & din_b[161]) ) + ( Xd_0__inst_mult_28_102  ) + ( Xd_0__inst_mult_28_101  ))
// Xd_0__inst_mult_23_85  = CARRY(( (din_a[161] & din_b[161]) ) + ( Xd_0__inst_mult_28_102  ) + ( Xd_0__inst_mult_28_101  ))
// Xd_0__inst_mult_23_86  = SHARE((din_a[161] & din_b[162]))

	.dataa(!din_a[161]),
	.datab(!din_b[161]),
	.datac(!din_b[162]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_101 ),
	.sharein(Xd_0__inst_mult_28_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_84 ),
	.cout(Xd_0__inst_mult_23_85 ),
	.shareout(Xd_0__inst_mult_23_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_28 (
// Equation(s):
// Xd_0__inst_mult_20_84  = SUM(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_12_102  ) + ( Xd_0__inst_mult_12_101  ))
// Xd_0__inst_mult_20_85  = CARRY(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_12_102  ) + ( Xd_0__inst_mult_12_101  ))
// Xd_0__inst_mult_20_86  = SHARE((din_a[140] & din_b[141]))

	.dataa(!din_a[140]),
	.datab(!din_b[140]),
	.datac(!din_b[141]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_101 ),
	.sharein(Xd_0__inst_mult_12_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_84 ),
	.cout(Xd_0__inst_mult_20_85 ),
	.shareout(Xd_0__inst_mult_20_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_28 (
// Equation(s):
// Xd_0__inst_mult_21_84  = SUM(( (din_a[147] & din_b[147]) ) + ( Xd_0__inst_mult_5_102  ) + ( Xd_0__inst_mult_5_101  ))
// Xd_0__inst_mult_21_85  = CARRY(( (din_a[147] & din_b[147]) ) + ( Xd_0__inst_mult_5_102  ) + ( Xd_0__inst_mult_5_101  ))
// Xd_0__inst_mult_21_86  = SHARE((din_a[147] & din_b[148]))

	.dataa(!din_a[147]),
	.datab(!din_b[147]),
	.datac(!din_b[148]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_101 ),
	.sharein(Xd_0__inst_mult_5_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_84 ),
	.cout(Xd_0__inst_mult_21_85 ),
	.shareout(Xd_0__inst_mult_21_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_28 (
// Equation(s):
// Xd_0__inst_mult_18_84  = SUM(( (din_a[126] & din_b[126]) ) + ( Xd_0__inst_mult_15_102  ) + ( Xd_0__inst_mult_15_101  ))
// Xd_0__inst_mult_18_85  = CARRY(( (din_a[126] & din_b[126]) ) + ( Xd_0__inst_mult_15_102  ) + ( Xd_0__inst_mult_15_101  ))
// Xd_0__inst_mult_18_86  = SHARE((din_a[126] & din_b[127]))

	.dataa(!din_a[126]),
	.datab(!din_b[126]),
	.datac(!din_b[127]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_101 ),
	.sharein(Xd_0__inst_mult_15_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_84 ),
	.cout(Xd_0__inst_mult_18_85 ),
	.shareout(Xd_0__inst_mult_18_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_28 (
// Equation(s):
// Xd_0__inst_mult_19_84  = SUM(( (din_a[133] & din_b[133]) ) + ( Xd_0__inst_mult_7_102  ) + ( Xd_0__inst_mult_7_101  ))
// Xd_0__inst_mult_19_85  = CARRY(( (din_a[133] & din_b[133]) ) + ( Xd_0__inst_mult_7_102  ) + ( Xd_0__inst_mult_7_101  ))
// Xd_0__inst_mult_19_86  = SHARE((din_a[133] & din_b[134]))

	.dataa(!din_a[133]),
	.datab(!din_b[133]),
	.datac(!din_b[134]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_101 ),
	.sharein(Xd_0__inst_mult_7_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_84 ),
	.cout(Xd_0__inst_mult_19_85 ),
	.shareout(Xd_0__inst_mult_19_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_29 (
// Equation(s):
// Xd_0__inst_mult_25_88  = SUM(( GND ) + ( Xd_0__inst_mult_25_106  ) + ( Xd_0__inst_mult_25_105  ))
// Xd_0__inst_mult_25_89  = CARRY(( GND ) + ( Xd_0__inst_mult_25_106  ) + ( Xd_0__inst_mult_25_105  ))
// Xd_0__inst_mult_25_90  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_105 ),
	.sharein(Xd_0__inst_mult_25_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_88 ),
	.cout(Xd_0__inst_mult_25_89 ),
	.shareout(Xd_0__inst_mult_25_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_29 (
// Equation(s):
// Xd_0__inst_mult_22_88  = SUM(( GND ) + ( Xd_0__inst_mult_22_106  ) + ( Xd_0__inst_mult_22_105  ))
// Xd_0__inst_mult_22_89  = CARRY(( GND ) + ( Xd_0__inst_mult_22_106  ) + ( Xd_0__inst_mult_22_105  ))
// Xd_0__inst_mult_22_90  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_105 ),
	.sharein(Xd_0__inst_mult_22_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_88 ),
	.cout(Xd_0__inst_mult_22_89 ),
	.shareout(Xd_0__inst_mult_22_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_28 (
// Equation(s):
// Xd_0__inst_mult_16_84  = SUM(( (din_a[112] & din_b[112]) ) + ( Xd_0__inst_mult_6_102  ) + ( Xd_0__inst_mult_6_101  ))
// Xd_0__inst_mult_16_85  = CARRY(( (din_a[112] & din_b[112]) ) + ( Xd_0__inst_mult_6_102  ) + ( Xd_0__inst_mult_6_101  ))
// Xd_0__inst_mult_16_86  = SHARE((din_a[112] & din_b[113]))

	.dataa(!din_a[112]),
	.datab(!din_b[112]),
	.datac(!din_b[113]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_101 ),
	.sharein(Xd_0__inst_mult_6_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_84 ),
	.cout(Xd_0__inst_mult_16_85 ),
	.shareout(Xd_0__inst_mult_16_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_28 (
// Equation(s):
// Xd_0__inst_mult_17_84  = SUM(( (din_a[119] & din_b[119]) ) + ( Xd_0__inst_mult_9_102  ) + ( Xd_0__inst_mult_9_101  ))
// Xd_0__inst_mult_17_85  = CARRY(( (din_a[119] & din_b[119]) ) + ( Xd_0__inst_mult_9_102  ) + ( Xd_0__inst_mult_9_101  ))
// Xd_0__inst_mult_17_86  = SHARE((din_a[119] & din_b[120]))

	.dataa(!din_a[119]),
	.datab(!din_b[119]),
	.datac(!din_b[120]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_101 ),
	.sharein(Xd_0__inst_mult_9_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_84 ),
	.cout(Xd_0__inst_mult_17_85 ),
	.shareout(Xd_0__inst_mult_17_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_28 (
// Equation(s):
// Xd_0__inst_mult_14_84  = SUM(( (din_a[98] & din_b[98]) ) + ( Xd_0__inst_mult_8_102  ) + ( Xd_0__inst_mult_8_101  ))
// Xd_0__inst_mult_14_85  = CARRY(( (din_a[98] & din_b[98]) ) + ( Xd_0__inst_mult_8_102  ) + ( Xd_0__inst_mult_8_101  ))
// Xd_0__inst_mult_14_86  = SHARE((din_a[98] & din_b[99]))

	.dataa(!din_a[98]),
	.datab(!din_b[98]),
	.datac(!din_b[99]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_101 ),
	.sharein(Xd_0__inst_mult_8_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_84 ),
	.cout(Xd_0__inst_mult_14_85 ),
	.shareout(Xd_0__inst_mult_14_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_28 (
// Equation(s):
// Xd_0__inst_mult_15_84  = SUM(( (din_a[105] & din_b[105]) ) + ( Xd_0__inst_mult_11_102  ) + ( Xd_0__inst_mult_11_101  ))
// Xd_0__inst_mult_15_85  = CARRY(( (din_a[105] & din_b[105]) ) + ( Xd_0__inst_mult_11_102  ) + ( Xd_0__inst_mult_11_101  ))
// Xd_0__inst_mult_15_86  = SHARE((din_a[105] & din_b[106]))

	.dataa(!din_a[105]),
	.datab(!din_b[105]),
	.datac(!din_b[106]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_101 ),
	.sharein(Xd_0__inst_mult_11_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_84 ),
	.cout(Xd_0__inst_mult_15_85 ),
	.shareout(Xd_0__inst_mult_15_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_28 (
// Equation(s):
// Xd_0__inst_mult_12_84  = SUM(( (din_a[84] & din_b[84]) ) + ( Xd_0__inst_mult_10_102  ) + ( Xd_0__inst_mult_10_101  ))
// Xd_0__inst_mult_12_85  = CARRY(( (din_a[84] & din_b[84]) ) + ( Xd_0__inst_mult_10_102  ) + ( Xd_0__inst_mult_10_101  ))
// Xd_0__inst_mult_12_86  = SHARE((din_a[84] & din_b[85]))

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_101 ),
	.sharein(Xd_0__inst_mult_10_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_84 ),
	.cout(Xd_0__inst_mult_12_85 ),
	.shareout(Xd_0__inst_mult_12_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_28 (
// Equation(s):
// Xd_0__inst_mult_13_84  = SUM(( (din_a[91] & din_b[91]) ) + ( Xd_0__inst_mult_13_102  ) + ( Xd_0__inst_mult_13_101  ))
// Xd_0__inst_mult_13_85  = CARRY(( (din_a[91] & din_b[91]) ) + ( Xd_0__inst_mult_13_102  ) + ( Xd_0__inst_mult_13_101  ))
// Xd_0__inst_mult_13_86  = SHARE((din_a[91] & din_b[92]))

	.dataa(!din_a[91]),
	.datab(!din_b[91]),
	.datac(!din_b[92]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_101 ),
	.sharein(Xd_0__inst_mult_13_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_84 ),
	.cout(Xd_0__inst_mult_13_85 ),
	.shareout(Xd_0__inst_mult_13_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_28 (
// Equation(s):
// Xd_0__inst_mult_10_84  = SUM(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_4_102  ) + ( Xd_0__inst_mult_4_101  ))
// Xd_0__inst_mult_10_85  = CARRY(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_4_102  ) + ( Xd_0__inst_mult_4_101  ))
// Xd_0__inst_mult_10_86  = SHARE((din_a[70] & din_b[71]))

	.dataa(!din_a[70]),
	.datab(!din_b[70]),
	.datac(!din_b[71]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_101 ),
	.sharein(Xd_0__inst_mult_4_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_84 ),
	.cout(Xd_0__inst_mult_10_85 ),
	.shareout(Xd_0__inst_mult_10_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_28 (
// Equation(s):
// Xd_0__inst_mult_11_84  = SUM(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_2_102  ) + ( Xd_0__inst_mult_2_101  ))
// Xd_0__inst_mult_11_85  = CARRY(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_2_102  ) + ( Xd_0__inst_mult_2_101  ))
// Xd_0__inst_mult_11_86  = SHARE((din_a[77] & din_b[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_101 ),
	.sharein(Xd_0__inst_mult_2_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_84 ),
	.cout(Xd_0__inst_mult_11_85 ),
	.shareout(Xd_0__inst_mult_11_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_28 (
// Equation(s):
// Xd_0__inst_mult_8_84  = SUM(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_3_102  ) + ( Xd_0__inst_mult_3_101  ))
// Xd_0__inst_mult_8_85  = CARRY(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_3_102  ) + ( Xd_0__inst_mult_3_101  ))
// Xd_0__inst_mult_8_86  = SHARE((din_a[56] & din_b[57]))

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(!din_b[57]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_101 ),
	.sharein(Xd_0__inst_mult_3_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_84 ),
	.cout(Xd_0__inst_mult_8_85 ),
	.shareout(Xd_0__inst_mult_8_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_28 (
// Equation(s):
// Xd_0__inst_mult_9_84  = SUM(( (din_a[63] & din_b[63]) ) + ( Xd_0__inst_mult_0_102  ) + ( Xd_0__inst_mult_0_101  ))
// Xd_0__inst_mult_9_85  = CARRY(( (din_a[63] & din_b[63]) ) + ( Xd_0__inst_mult_0_102  ) + ( Xd_0__inst_mult_0_101  ))
// Xd_0__inst_mult_9_86  = SHARE((din_a[63] & din_b[64]))

	.dataa(!din_a[63]),
	.datab(!din_b[63]),
	.datac(!din_b[64]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_101 ),
	.sharein(Xd_0__inst_mult_0_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_84 ),
	.cout(Xd_0__inst_mult_9_85 ),
	.shareout(Xd_0__inst_mult_9_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_28 (
// Equation(s):
// Xd_0__inst_mult_6_84  = SUM(( (din_a[42] & din_b[42]) ) + ( Xd_0__inst_mult_1_102  ) + ( Xd_0__inst_mult_1_101  ))
// Xd_0__inst_mult_6_85  = CARRY(( (din_a[42] & din_b[42]) ) + ( Xd_0__inst_mult_1_102  ) + ( Xd_0__inst_mult_1_101  ))
// Xd_0__inst_mult_6_86  = SHARE((din_a[42] & din_b[43]))

	.dataa(!din_a[42]),
	.datab(!din_b[42]),
	.datac(!din_b[43]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_101 ),
	.sharein(Xd_0__inst_mult_1_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_84 ),
	.cout(Xd_0__inst_mult_6_85 ),
	.shareout(Xd_0__inst_mult_6_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_28 (
// Equation(s):
// Xd_0__inst_mult_7_84  = SUM(( (din_a[49] & din_b[49]) ) + ( Xd_0__inst_mult_23_102  ) + ( Xd_0__inst_mult_23_101  ))
// Xd_0__inst_mult_7_85  = CARRY(( (din_a[49] & din_b[49]) ) + ( Xd_0__inst_mult_23_102  ) + ( Xd_0__inst_mult_23_101  ))
// Xd_0__inst_mult_7_86  = SHARE((din_a[49] & din_b[50]))

	.dataa(!din_a[49]),
	.datab(!din_b[49]),
	.datac(!din_b[50]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_101 ),
	.sharein(Xd_0__inst_mult_23_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_84 ),
	.cout(Xd_0__inst_mult_7_85 ),
	.shareout(Xd_0__inst_mult_7_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_28 (
// Equation(s):
// Xd_0__inst_mult_4_84  = SUM(( (din_a[28] & din_b[28]) ) + ( Xd_0__inst_mult_29_102  ) + ( Xd_0__inst_mult_29_101  ))
// Xd_0__inst_mult_4_85  = CARRY(( (din_a[28] & din_b[28]) ) + ( Xd_0__inst_mult_29_102  ) + ( Xd_0__inst_mult_29_101  ))
// Xd_0__inst_mult_4_86  = SHARE((din_a[28] & din_b[29]))

	.dataa(!din_a[28]),
	.datab(!din_b[28]),
	.datac(!din_b[29]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_101 ),
	.sharein(Xd_0__inst_mult_29_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_84 ),
	.cout(Xd_0__inst_mult_4_85 ),
	.shareout(Xd_0__inst_mult_4_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_28 (
// Equation(s):
// Xd_0__inst_mult_5_84  = SUM(( (din_a[35] & din_b[35]) ) + ( Xd_0__inst_mult_31_150  ) + ( Xd_0__inst_mult_31_149  ))
// Xd_0__inst_mult_5_85  = CARRY(( (din_a[35] & din_b[35]) ) + ( Xd_0__inst_mult_31_150  ) + ( Xd_0__inst_mult_31_149  ))
// Xd_0__inst_mult_5_86  = SHARE((din_a[35] & din_b[36]))

	.dataa(!din_a[35]),
	.datab(!din_b[35]),
	.datac(!din_b[36]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_149 ),
	.sharein(Xd_0__inst_mult_31_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_84 ),
	.cout(Xd_0__inst_mult_5_85 ),
	.shareout(Xd_0__inst_mult_5_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_113 (
// Equation(s):
// Xd_0__inst_i19_113_sumout  = SUM(( !din_a[34] $ (!din_b[34]) ) + ( Xd_0__inst_i19_119  ) + ( Xd_0__inst_i19_118  ))
// Xd_0__inst_i19_114  = CARRY(( !din_a[34] $ (!din_b[34]) ) + ( Xd_0__inst_i19_119  ) + ( Xd_0__inst_i19_118  ))
// Xd_0__inst_i19_115  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_118 ),
	.sharein(Xd_0__inst_i19_119 ),
	.combout(),
	.sumout(Xd_0__inst_i19_113_sumout ),
	.cout(Xd_0__inst_i19_114 ),
	.shareout(Xd_0__inst_i19_115 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_117 (
// Equation(s):
// Xd_0__inst_i19_117_sumout  = SUM(( !din_a[41] $ (!din_b[41]) ) + ( Xd_0__inst_i19_123  ) + ( Xd_0__inst_i19_122  ))
// Xd_0__inst_i19_118  = CARRY(( !din_a[41] $ (!din_b[41]) ) + ( Xd_0__inst_i19_123  ) + ( Xd_0__inst_i19_122  ))
// Xd_0__inst_i19_119  = SHARE(GND)

	.dataa(!din_a[41]),
	.datab(!din_b[41]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_122 ),
	.sharein(Xd_0__inst_i19_123 ),
	.combout(),
	.sumout(Xd_0__inst_i19_117_sumout ),
	.cout(Xd_0__inst_i19_118 ),
	.shareout(Xd_0__inst_i19_119 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_28 (
// Equation(s):
// Xd_0__inst_mult_2_84  = SUM(( (din_a[14] & din_b[14]) ) + ( Xd_0__inst_mult_30_150  ) + ( Xd_0__inst_mult_30_149  ))
// Xd_0__inst_mult_2_85  = CARRY(( (din_a[14] & din_b[14]) ) + ( Xd_0__inst_mult_30_150  ) + ( Xd_0__inst_mult_30_149  ))
// Xd_0__inst_mult_2_86  = SHARE((din_a[14] & din_b[15]))

	.dataa(!din_a[14]),
	.datab(!din_b[14]),
	.datac(!din_b[15]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_149 ),
	.sharein(Xd_0__inst_mult_30_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_84 ),
	.cout(Xd_0__inst_mult_2_85 ),
	.shareout(Xd_0__inst_mult_2_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_28 (
// Equation(s):
// Xd_0__inst_mult_3_84  = SUM(( (din_a[21] & din_b[21]) ) + ( Xd_0__inst_mult_26_102  ) + ( Xd_0__inst_mult_26_101  ))
// Xd_0__inst_mult_3_85  = CARRY(( (din_a[21] & din_b[21]) ) + ( Xd_0__inst_mult_26_102  ) + ( Xd_0__inst_mult_26_101  ))
// Xd_0__inst_mult_3_86  = SHARE((din_a[21] & din_b[22]))

	.dataa(!din_a[21]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_101 ),
	.sharein(Xd_0__inst_mult_26_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_84 ),
	.cout(Xd_0__inst_mult_3_85 ),
	.shareout(Xd_0__inst_mult_3_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_121 (
// Equation(s):
// Xd_0__inst_i19_121_sumout  = SUM(( !din_a[20] $ (!din_b[20]) ) + ( Xd_0__inst_i19_127  ) + ( Xd_0__inst_i19_126  ))
// Xd_0__inst_i19_122  = CARRY(( !din_a[20] $ (!din_b[20]) ) + ( Xd_0__inst_i19_127  ) + ( Xd_0__inst_i19_126  ))
// Xd_0__inst_i19_123  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i19_126 ),
	.sharein(Xd_0__inst_i19_127 ),
	.combout(),
	.sumout(Xd_0__inst_i19_121_sumout ),
	.cout(Xd_0__inst_i19_122 ),
	.shareout(Xd_0__inst_i19_123 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i19_125 (
// Equation(s):
// Xd_0__inst_i19_125_sumout  = SUM(( !din_a[27] $ (!din_b[27]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_126  = CARRY(( !din_a[27] $ (!din_b[27]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i19_127  = SHARE(GND)

	.dataa(!din_a[27]),
	.datab(!din_b[27]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i19_125_sumout ),
	.cout(Xd_0__inst_i19_126 ),
	.shareout(Xd_0__inst_i19_127 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_28 (
// Equation(s):
// Xd_0__inst_mult_0_84  = SUM(( (din_a[0] & din_b[0]) ) + ( Xd_0__inst_mult_24_102  ) + ( Xd_0__inst_mult_24_101  ))
// Xd_0__inst_mult_0_85  = CARRY(( (din_a[0] & din_b[0]) ) + ( Xd_0__inst_mult_24_102  ) + ( Xd_0__inst_mult_24_101  ))
// Xd_0__inst_mult_0_86  = SHARE((din_a[0] & din_b[1]))

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_101 ),
	.sharein(Xd_0__inst_mult_24_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_84 ),
	.cout(Xd_0__inst_mult_0_85 ),
	.shareout(Xd_0__inst_mult_0_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_28 (
// Equation(s):
// Xd_0__inst_mult_1_84  = SUM(( (din_a[7] & din_b[7]) ) + ( Xd_0__inst_mult_27_102  ) + ( Xd_0__inst_mult_27_101  ))
// Xd_0__inst_mult_1_85  = CARRY(( (din_a[7] & din_b[7]) ) + ( Xd_0__inst_mult_27_102  ) + ( Xd_0__inst_mult_27_101  ))
// Xd_0__inst_mult_1_86  = SHARE((din_a[7] & din_b[8]))

	.dataa(!din_a[7]),
	.datab(!din_b[7]),
	.datac(!din_b[8]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_101 ),
	.sharein(Xd_0__inst_mult_27_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_84 ),
	.cout(Xd_0__inst_mult_1_85 ),
	.shareout(Xd_0__inst_mult_1_86 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_29 (
// Equation(s):
// Xd_0__inst_mult_28_88  = SUM(( (din_a[197] & din_b[196]) ) + ( Xd_0__inst_mult_28_86  ) + ( Xd_0__inst_mult_28_85  ))
// Xd_0__inst_mult_28_89  = CARRY(( (din_a[197] & din_b[196]) ) + ( Xd_0__inst_mult_28_86  ) + ( Xd_0__inst_mult_28_85  ))
// Xd_0__inst_mult_28_90  = SHARE((din_a[196] & din_b[198]))

	.dataa(!din_a[197]),
	.datab(!din_b[196]),
	.datac(!din_a[196]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_85 ),
	.sharein(Xd_0__inst_mult_28_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_88 ),
	.cout(Xd_0__inst_mult_28_89 ),
	.shareout(Xd_0__inst_mult_28_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_29 (
// Equation(s):
// Xd_0__inst_mult_29_88  = SUM(( (din_a[204] & din_b[203]) ) + ( Xd_0__inst_mult_29_86  ) + ( Xd_0__inst_mult_29_85  ))
// Xd_0__inst_mult_29_89  = CARRY(( (din_a[204] & din_b[203]) ) + ( Xd_0__inst_mult_29_86  ) + ( Xd_0__inst_mult_29_85  ))
// Xd_0__inst_mult_29_90  = SHARE((din_a[203] & din_b[205]))

	.dataa(!din_a[204]),
	.datab(!din_b[203]),
	.datac(!din_a[203]),
	.datad(!din_b[205]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_85 ),
	.sharein(Xd_0__inst_mult_29_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_88 ),
	.cout(Xd_0__inst_mult_29_89 ),
	.shareout(Xd_0__inst_mult_29_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_29 (
// Equation(s):
// Xd_0__inst_mult_26_88  = SUM(( (din_a[183] & din_b[182]) ) + ( Xd_0__inst_mult_26_86  ) + ( Xd_0__inst_mult_26_85  ))
// Xd_0__inst_mult_26_89  = CARRY(( (din_a[183] & din_b[182]) ) + ( Xd_0__inst_mult_26_86  ) + ( Xd_0__inst_mult_26_85  ))
// Xd_0__inst_mult_26_90  = SHARE((din_a[182] & din_b[184]))

	.dataa(!din_a[183]),
	.datab(!din_b[182]),
	.datac(!din_a[182]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_85 ),
	.sharein(Xd_0__inst_mult_26_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_88 ),
	.cout(Xd_0__inst_mult_26_89 ),
	.shareout(Xd_0__inst_mult_26_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_29 (
// Equation(s):
// Xd_0__inst_mult_27_88  = SUM(( (din_a[190] & din_b[189]) ) + ( Xd_0__inst_mult_27_86  ) + ( Xd_0__inst_mult_27_85  ))
// Xd_0__inst_mult_27_89  = CARRY(( (din_a[190] & din_b[189]) ) + ( Xd_0__inst_mult_27_86  ) + ( Xd_0__inst_mult_27_85  ))
// Xd_0__inst_mult_27_90  = SHARE((din_a[189] & din_b[191]))

	.dataa(!din_a[190]),
	.datab(!din_b[189]),
	.datac(!din_a[189]),
	.datad(!din_b[191]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_85 ),
	.sharein(Xd_0__inst_mult_27_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_88 ),
	.cout(Xd_0__inst_mult_27_89 ),
	.shareout(Xd_0__inst_mult_27_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_29 (
// Equation(s):
// Xd_0__inst_mult_24_88  = SUM(( (din_a[169] & din_b[168]) ) + ( Xd_0__inst_mult_24_86  ) + ( Xd_0__inst_mult_24_85  ))
// Xd_0__inst_mult_24_89  = CARRY(( (din_a[169] & din_b[168]) ) + ( Xd_0__inst_mult_24_86  ) + ( Xd_0__inst_mult_24_85  ))
// Xd_0__inst_mult_24_90  = SHARE((din_a[168] & din_b[170]))

	.dataa(!din_a[169]),
	.datab(!din_b[168]),
	.datac(!din_a[168]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_85 ),
	.sharein(Xd_0__inst_mult_24_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_88 ),
	.cout(Xd_0__inst_mult_24_89 ),
	.shareout(Xd_0__inst_mult_24_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_30 (
// Equation(s):
// Xd_0__inst_mult_25_92  = SUM(( (din_a[176] & din_b[175]) ) + ( Xd_0__inst_mult_25_86  ) + ( Xd_0__inst_mult_25_85  ))
// Xd_0__inst_mult_25_93  = CARRY(( (din_a[176] & din_b[175]) ) + ( Xd_0__inst_mult_25_86  ) + ( Xd_0__inst_mult_25_85  ))
// Xd_0__inst_mult_25_94  = SHARE((din_a[175] & din_b[177]))

	.dataa(!din_a[176]),
	.datab(!din_b[175]),
	.datac(!din_a[175]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_85 ),
	.sharein(Xd_0__inst_mult_25_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_92 ),
	.cout(Xd_0__inst_mult_25_93 ),
	.shareout(Xd_0__inst_mult_25_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_30 (
// Equation(s):
// Xd_0__inst_mult_22_92  = SUM(( (din_a[155] & din_b[154]) ) + ( Xd_0__inst_mult_22_86  ) + ( Xd_0__inst_mult_22_85  ))
// Xd_0__inst_mult_22_93  = CARRY(( (din_a[155] & din_b[154]) ) + ( Xd_0__inst_mult_22_86  ) + ( Xd_0__inst_mult_22_85  ))
// Xd_0__inst_mult_22_94  = SHARE((din_a[154] & din_b[156]))

	.dataa(!din_a[155]),
	.datab(!din_b[154]),
	.datac(!din_a[154]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_85 ),
	.sharein(Xd_0__inst_mult_22_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_92 ),
	.cout(Xd_0__inst_mult_22_93 ),
	.shareout(Xd_0__inst_mult_22_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_29 (
// Equation(s):
// Xd_0__inst_mult_23_88  = SUM(( (din_a[162] & din_b[161]) ) + ( Xd_0__inst_mult_23_86  ) + ( Xd_0__inst_mult_23_85  ))
// Xd_0__inst_mult_23_89  = CARRY(( (din_a[162] & din_b[161]) ) + ( Xd_0__inst_mult_23_86  ) + ( Xd_0__inst_mult_23_85  ))
// Xd_0__inst_mult_23_90  = SHARE((din_a[161] & din_b[163]))

	.dataa(!din_a[162]),
	.datab(!din_b[161]),
	.datac(!din_a[161]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_85 ),
	.sharein(Xd_0__inst_mult_23_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_88 ),
	.cout(Xd_0__inst_mult_23_89 ),
	.shareout(Xd_0__inst_mult_23_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_29 (
// Equation(s):
// Xd_0__inst_mult_20_88  = SUM(( (din_a[141] & din_b[140]) ) + ( Xd_0__inst_mult_20_86  ) + ( Xd_0__inst_mult_20_85  ))
// Xd_0__inst_mult_20_89  = CARRY(( (din_a[141] & din_b[140]) ) + ( Xd_0__inst_mult_20_86  ) + ( Xd_0__inst_mult_20_85  ))
// Xd_0__inst_mult_20_90  = SHARE((din_a[140] & din_b[142]))

	.dataa(!din_a[141]),
	.datab(!din_b[140]),
	.datac(!din_a[140]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_85 ),
	.sharein(Xd_0__inst_mult_20_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_88 ),
	.cout(Xd_0__inst_mult_20_89 ),
	.shareout(Xd_0__inst_mult_20_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_29 (
// Equation(s):
// Xd_0__inst_mult_21_88  = SUM(( (din_a[148] & din_b[147]) ) + ( Xd_0__inst_mult_21_86  ) + ( Xd_0__inst_mult_21_85  ))
// Xd_0__inst_mult_21_89  = CARRY(( (din_a[148] & din_b[147]) ) + ( Xd_0__inst_mult_21_86  ) + ( Xd_0__inst_mult_21_85  ))
// Xd_0__inst_mult_21_90  = SHARE((din_a[147] & din_b[149]))

	.dataa(!din_a[148]),
	.datab(!din_b[147]),
	.datac(!din_a[147]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_85 ),
	.sharein(Xd_0__inst_mult_21_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_88 ),
	.cout(Xd_0__inst_mult_21_89 ),
	.shareout(Xd_0__inst_mult_21_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_29 (
// Equation(s):
// Xd_0__inst_mult_18_88  = SUM(( (din_a[127] & din_b[126]) ) + ( Xd_0__inst_mult_18_86  ) + ( Xd_0__inst_mult_18_85  ))
// Xd_0__inst_mult_18_89  = CARRY(( (din_a[127] & din_b[126]) ) + ( Xd_0__inst_mult_18_86  ) + ( Xd_0__inst_mult_18_85  ))
// Xd_0__inst_mult_18_90  = SHARE((din_a[126] & din_b[128]))

	.dataa(!din_a[127]),
	.datab(!din_b[126]),
	.datac(!din_a[126]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_85 ),
	.sharein(Xd_0__inst_mult_18_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_88 ),
	.cout(Xd_0__inst_mult_18_89 ),
	.shareout(Xd_0__inst_mult_18_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_29 (
// Equation(s):
// Xd_0__inst_mult_19_88  = SUM(( (din_a[134] & din_b[133]) ) + ( Xd_0__inst_mult_19_86  ) + ( Xd_0__inst_mult_19_85  ))
// Xd_0__inst_mult_19_89  = CARRY(( (din_a[134] & din_b[133]) ) + ( Xd_0__inst_mult_19_86  ) + ( Xd_0__inst_mult_19_85  ))
// Xd_0__inst_mult_19_90  = SHARE((din_a[133] & din_b[135]))

	.dataa(!din_a[134]),
	.datab(!din_b[133]),
	.datac(!din_a[133]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_85 ),
	.sharein(Xd_0__inst_mult_19_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_88 ),
	.cout(Xd_0__inst_mult_19_89 ),
	.shareout(Xd_0__inst_mult_19_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_29 (
// Equation(s):
// Xd_0__inst_mult_16_88  = SUM(( (din_a[113] & din_b[112]) ) + ( Xd_0__inst_mult_16_86  ) + ( Xd_0__inst_mult_16_85  ))
// Xd_0__inst_mult_16_89  = CARRY(( (din_a[113] & din_b[112]) ) + ( Xd_0__inst_mult_16_86  ) + ( Xd_0__inst_mult_16_85  ))
// Xd_0__inst_mult_16_90  = SHARE((din_a[112] & din_b[114]))

	.dataa(!din_a[113]),
	.datab(!din_b[112]),
	.datac(!din_a[112]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_85 ),
	.sharein(Xd_0__inst_mult_16_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_88 ),
	.cout(Xd_0__inst_mult_16_89 ),
	.shareout(Xd_0__inst_mult_16_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_29 (
// Equation(s):
// Xd_0__inst_mult_17_88  = SUM(( (din_a[120] & din_b[119]) ) + ( Xd_0__inst_mult_17_86  ) + ( Xd_0__inst_mult_17_85  ))
// Xd_0__inst_mult_17_89  = CARRY(( (din_a[120] & din_b[119]) ) + ( Xd_0__inst_mult_17_86  ) + ( Xd_0__inst_mult_17_85  ))
// Xd_0__inst_mult_17_90  = SHARE((din_a[119] & din_b[121]))

	.dataa(!din_a[120]),
	.datab(!din_b[119]),
	.datac(!din_a[119]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_85 ),
	.sharein(Xd_0__inst_mult_17_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_88 ),
	.cout(Xd_0__inst_mult_17_89 ),
	.shareout(Xd_0__inst_mult_17_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_29 (
// Equation(s):
// Xd_0__inst_mult_14_88  = SUM(( (din_a[99] & din_b[98]) ) + ( Xd_0__inst_mult_14_86  ) + ( Xd_0__inst_mult_14_85  ))
// Xd_0__inst_mult_14_89  = CARRY(( (din_a[99] & din_b[98]) ) + ( Xd_0__inst_mult_14_86  ) + ( Xd_0__inst_mult_14_85  ))
// Xd_0__inst_mult_14_90  = SHARE((din_a[98] & din_b[100]))

	.dataa(!din_a[99]),
	.datab(!din_b[98]),
	.datac(!din_a[98]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_85 ),
	.sharein(Xd_0__inst_mult_14_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_88 ),
	.cout(Xd_0__inst_mult_14_89 ),
	.shareout(Xd_0__inst_mult_14_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_29 (
// Equation(s):
// Xd_0__inst_mult_15_88  = SUM(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_15_86  ) + ( Xd_0__inst_mult_15_85  ))
// Xd_0__inst_mult_15_89  = CARRY(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_15_86  ) + ( Xd_0__inst_mult_15_85  ))
// Xd_0__inst_mult_15_90  = SHARE((din_a[105] & din_b[107]))

	.dataa(!din_a[106]),
	.datab(!din_b[105]),
	.datac(!din_a[105]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_85 ),
	.sharein(Xd_0__inst_mult_15_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_88 ),
	.cout(Xd_0__inst_mult_15_89 ),
	.shareout(Xd_0__inst_mult_15_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_29 (
// Equation(s):
// Xd_0__inst_mult_12_88  = SUM(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_12_86  ) + ( Xd_0__inst_mult_12_85  ))
// Xd_0__inst_mult_12_89  = CARRY(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_12_86  ) + ( Xd_0__inst_mult_12_85  ))
// Xd_0__inst_mult_12_90  = SHARE((din_a[84] & din_b[86]))

	.dataa(!din_a[85]),
	.datab(!din_b[84]),
	.datac(!din_a[84]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_85 ),
	.sharein(Xd_0__inst_mult_12_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_88 ),
	.cout(Xd_0__inst_mult_12_89 ),
	.shareout(Xd_0__inst_mult_12_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_29 (
// Equation(s):
// Xd_0__inst_mult_13_88  = SUM(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_13_86  ) + ( Xd_0__inst_mult_13_85  ))
// Xd_0__inst_mult_13_89  = CARRY(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_13_86  ) + ( Xd_0__inst_mult_13_85  ))
// Xd_0__inst_mult_13_90  = SHARE((din_a[91] & din_b[93]))

	.dataa(!din_a[92]),
	.datab(!din_b[91]),
	.datac(!din_a[91]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_85 ),
	.sharein(Xd_0__inst_mult_13_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_88 ),
	.cout(Xd_0__inst_mult_13_89 ),
	.shareout(Xd_0__inst_mult_13_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_29 (
// Equation(s):
// Xd_0__inst_mult_10_88  = SUM(( (din_a[71] & din_b[70]) ) + ( Xd_0__inst_mult_10_86  ) + ( Xd_0__inst_mult_10_85  ))
// Xd_0__inst_mult_10_89  = CARRY(( (din_a[71] & din_b[70]) ) + ( Xd_0__inst_mult_10_86  ) + ( Xd_0__inst_mult_10_85  ))
// Xd_0__inst_mult_10_90  = SHARE((din_a[70] & din_b[72]))

	.dataa(!din_a[71]),
	.datab(!din_b[70]),
	.datac(!din_a[70]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_85 ),
	.sharein(Xd_0__inst_mult_10_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_88 ),
	.cout(Xd_0__inst_mult_10_89 ),
	.shareout(Xd_0__inst_mult_10_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_29 (
// Equation(s):
// Xd_0__inst_mult_11_88  = SUM(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_11_86  ) + ( Xd_0__inst_mult_11_85  ))
// Xd_0__inst_mult_11_89  = CARRY(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_11_86  ) + ( Xd_0__inst_mult_11_85  ))
// Xd_0__inst_mult_11_90  = SHARE((din_a[77] & din_b[79]))

	.dataa(!din_a[78]),
	.datab(!din_b[77]),
	.datac(!din_a[77]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_85 ),
	.sharein(Xd_0__inst_mult_11_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_88 ),
	.cout(Xd_0__inst_mult_11_89 ),
	.shareout(Xd_0__inst_mult_11_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_29 (
// Equation(s):
// Xd_0__inst_mult_8_88  = SUM(( (din_a[57] & din_b[56]) ) + ( Xd_0__inst_mult_8_86  ) + ( Xd_0__inst_mult_8_85  ))
// Xd_0__inst_mult_8_89  = CARRY(( (din_a[57] & din_b[56]) ) + ( Xd_0__inst_mult_8_86  ) + ( Xd_0__inst_mult_8_85  ))
// Xd_0__inst_mult_8_90  = SHARE((din_a[56] & din_b[58]))

	.dataa(!din_a[57]),
	.datab(!din_b[56]),
	.datac(!din_a[56]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_85 ),
	.sharein(Xd_0__inst_mult_8_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_88 ),
	.cout(Xd_0__inst_mult_8_89 ),
	.shareout(Xd_0__inst_mult_8_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_29 (
// Equation(s):
// Xd_0__inst_mult_9_88  = SUM(( (din_a[64] & din_b[63]) ) + ( Xd_0__inst_mult_9_86  ) + ( Xd_0__inst_mult_9_85  ))
// Xd_0__inst_mult_9_89  = CARRY(( (din_a[64] & din_b[63]) ) + ( Xd_0__inst_mult_9_86  ) + ( Xd_0__inst_mult_9_85  ))
// Xd_0__inst_mult_9_90  = SHARE((din_a[63] & din_b[65]))

	.dataa(!din_a[64]),
	.datab(!din_b[63]),
	.datac(!din_a[63]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_85 ),
	.sharein(Xd_0__inst_mult_9_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_88 ),
	.cout(Xd_0__inst_mult_9_89 ),
	.shareout(Xd_0__inst_mult_9_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_29 (
// Equation(s):
// Xd_0__inst_mult_6_88  = SUM(( (din_a[43] & din_b[42]) ) + ( Xd_0__inst_mult_6_86  ) + ( Xd_0__inst_mult_6_85  ))
// Xd_0__inst_mult_6_89  = CARRY(( (din_a[43] & din_b[42]) ) + ( Xd_0__inst_mult_6_86  ) + ( Xd_0__inst_mult_6_85  ))
// Xd_0__inst_mult_6_90  = SHARE((din_a[42] & din_b[44]))

	.dataa(!din_a[43]),
	.datab(!din_b[42]),
	.datac(!din_a[42]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_85 ),
	.sharein(Xd_0__inst_mult_6_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_88 ),
	.cout(Xd_0__inst_mult_6_89 ),
	.shareout(Xd_0__inst_mult_6_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_29 (
// Equation(s):
// Xd_0__inst_mult_7_88  = SUM(( (din_a[50] & din_b[49]) ) + ( Xd_0__inst_mult_7_86  ) + ( Xd_0__inst_mult_7_85  ))
// Xd_0__inst_mult_7_89  = CARRY(( (din_a[50] & din_b[49]) ) + ( Xd_0__inst_mult_7_86  ) + ( Xd_0__inst_mult_7_85  ))
// Xd_0__inst_mult_7_90  = SHARE((din_a[49] & din_b[51]))

	.dataa(!din_a[50]),
	.datab(!din_b[49]),
	.datac(!din_a[49]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_85 ),
	.sharein(Xd_0__inst_mult_7_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_88 ),
	.cout(Xd_0__inst_mult_7_89 ),
	.shareout(Xd_0__inst_mult_7_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_29 (
// Equation(s):
// Xd_0__inst_mult_4_88  = SUM(( (din_a[29] & din_b[28]) ) + ( Xd_0__inst_mult_4_86  ) + ( Xd_0__inst_mult_4_85  ))
// Xd_0__inst_mult_4_89  = CARRY(( (din_a[29] & din_b[28]) ) + ( Xd_0__inst_mult_4_86  ) + ( Xd_0__inst_mult_4_85  ))
// Xd_0__inst_mult_4_90  = SHARE((din_a[28] & din_b[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[28]),
	.datac(!din_a[28]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_85 ),
	.sharein(Xd_0__inst_mult_4_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_88 ),
	.cout(Xd_0__inst_mult_4_89 ),
	.shareout(Xd_0__inst_mult_4_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_29 (
// Equation(s):
// Xd_0__inst_mult_5_88  = SUM(( (din_a[36] & din_b[35]) ) + ( Xd_0__inst_mult_5_86  ) + ( Xd_0__inst_mult_5_85  ))
// Xd_0__inst_mult_5_89  = CARRY(( (din_a[36] & din_b[35]) ) + ( Xd_0__inst_mult_5_86  ) + ( Xd_0__inst_mult_5_85  ))
// Xd_0__inst_mult_5_90  = SHARE((din_a[35] & din_b[37]))

	.dataa(!din_a[36]),
	.datab(!din_b[35]),
	.datac(!din_a[35]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_85 ),
	.sharein(Xd_0__inst_mult_5_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_88 ),
	.cout(Xd_0__inst_mult_5_89 ),
	.shareout(Xd_0__inst_mult_5_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_29 (
// Equation(s):
// Xd_0__inst_mult_2_88  = SUM(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_2_86  ) + ( Xd_0__inst_mult_2_85  ))
// Xd_0__inst_mult_2_89  = CARRY(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_2_86  ) + ( Xd_0__inst_mult_2_85  ))
// Xd_0__inst_mult_2_90  = SHARE((din_a[14] & din_b[16]))

	.dataa(!din_a[15]),
	.datab(!din_b[14]),
	.datac(!din_a[14]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_85 ),
	.sharein(Xd_0__inst_mult_2_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_88 ),
	.cout(Xd_0__inst_mult_2_89 ),
	.shareout(Xd_0__inst_mult_2_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_29 (
// Equation(s):
// Xd_0__inst_mult_3_88  = SUM(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_3_86  ) + ( Xd_0__inst_mult_3_85  ))
// Xd_0__inst_mult_3_89  = CARRY(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_3_86  ) + ( Xd_0__inst_mult_3_85  ))
// Xd_0__inst_mult_3_90  = SHARE((din_a[21] & din_b[23]))

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(!din_a[21]),
	.datad(!din_b[23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_85 ),
	.sharein(Xd_0__inst_mult_3_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_88 ),
	.cout(Xd_0__inst_mult_3_89 ),
	.shareout(Xd_0__inst_mult_3_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_29 (
// Equation(s):
// Xd_0__inst_mult_0_88  = SUM(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_86  ) + ( Xd_0__inst_mult_0_85  ))
// Xd_0__inst_mult_0_89  = CARRY(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_86  ) + ( Xd_0__inst_mult_0_85  ))
// Xd_0__inst_mult_0_90  = SHARE((din_a[0] & din_b[2]))

	.dataa(!din_a[1]),
	.datab(!din_b[0]),
	.datac(!din_a[0]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_85 ),
	.sharein(Xd_0__inst_mult_0_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_88 ),
	.cout(Xd_0__inst_mult_0_89 ),
	.shareout(Xd_0__inst_mult_0_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_29 (
// Equation(s):
// Xd_0__inst_mult_1_88  = SUM(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_1_86  ) + ( Xd_0__inst_mult_1_85  ))
// Xd_0__inst_mult_1_89  = CARRY(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_1_86  ) + ( Xd_0__inst_mult_1_85  ))
// Xd_0__inst_mult_1_90  = SHARE((din_a[7] & din_b[9]))

	.dataa(!din_a[8]),
	.datab(!din_b[7]),
	.datac(!din_a[7]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_85 ),
	.sharein(Xd_0__inst_mult_1_86 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_88 ),
	.cout(Xd_0__inst_mult_1_89 ),
	.shareout(Xd_0__inst_mult_1_90 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_30 (
// Equation(s):
// Xd_0__inst_mult_28_92  = SUM(( (!din_a[197] & (((din_a[198] & din_b[196])))) # (din_a[197] & (!din_b[197] $ (((!din_a[198]) # (!din_b[196]))))) ) + ( Xd_0__inst_mult_28_90  ) + ( Xd_0__inst_mult_28_89  ))
// Xd_0__inst_mult_28_93  = CARRY(( (!din_a[197] & (((din_a[198] & din_b[196])))) # (din_a[197] & (!din_b[197] $ (((!din_a[198]) # (!din_b[196]))))) ) + ( Xd_0__inst_mult_28_90  ) + ( Xd_0__inst_mult_28_89  ))
// Xd_0__inst_mult_28_94  = SHARE((din_a[197] & (din_b[197] & (din_a[198] & din_b[196]))))

	.dataa(!din_a[197]),
	.datab(!din_b[197]),
	.datac(!din_a[198]),
	.datad(!din_b[196]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_89 ),
	.sharein(Xd_0__inst_mult_28_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_92 ),
	.cout(Xd_0__inst_mult_28_93 ),
	.shareout(Xd_0__inst_mult_28_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_30 (
// Equation(s):
// Xd_0__inst_mult_29_92  = SUM(( (!din_a[204] & (((din_a[205] & din_b[203])))) # (din_a[204] & (!din_b[204] $ (((!din_a[205]) # (!din_b[203]))))) ) + ( Xd_0__inst_mult_29_90  ) + ( Xd_0__inst_mult_29_89  ))
// Xd_0__inst_mult_29_93  = CARRY(( (!din_a[204] & (((din_a[205] & din_b[203])))) # (din_a[204] & (!din_b[204] $ (((!din_a[205]) # (!din_b[203]))))) ) + ( Xd_0__inst_mult_29_90  ) + ( Xd_0__inst_mult_29_89  ))
// Xd_0__inst_mult_29_94  = SHARE((din_a[204] & (din_b[204] & (din_a[205] & din_b[203]))))

	.dataa(!din_a[204]),
	.datab(!din_b[204]),
	.datac(!din_a[205]),
	.datad(!din_b[203]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_89 ),
	.sharein(Xd_0__inst_mult_29_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_92 ),
	.cout(Xd_0__inst_mult_29_93 ),
	.shareout(Xd_0__inst_mult_29_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_30 (
// Equation(s):
// Xd_0__inst_mult_26_92  = SUM(( (!din_a[183] & (((din_a[184] & din_b[182])))) # (din_a[183] & (!din_b[183] $ (((!din_a[184]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_26_90  ) + ( Xd_0__inst_mult_26_89  ))
// Xd_0__inst_mult_26_93  = CARRY(( (!din_a[183] & (((din_a[184] & din_b[182])))) # (din_a[183] & (!din_b[183] $ (((!din_a[184]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_26_90  ) + ( Xd_0__inst_mult_26_89  ))
// Xd_0__inst_mult_26_94  = SHARE((din_a[183] & (din_b[183] & (din_a[184] & din_b[182]))))

	.dataa(!din_a[183]),
	.datab(!din_b[183]),
	.datac(!din_a[184]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_89 ),
	.sharein(Xd_0__inst_mult_26_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_92 ),
	.cout(Xd_0__inst_mult_26_93 ),
	.shareout(Xd_0__inst_mult_26_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_30 (
// Equation(s):
// Xd_0__inst_mult_27_92  = SUM(( (!din_a[190] & (((din_a[191] & din_b[189])))) # (din_a[190] & (!din_b[190] $ (((!din_a[191]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_27_90  ) + ( Xd_0__inst_mult_27_89  ))
// Xd_0__inst_mult_27_93  = CARRY(( (!din_a[190] & (((din_a[191] & din_b[189])))) # (din_a[190] & (!din_b[190] $ (((!din_a[191]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_27_90  ) + ( Xd_0__inst_mult_27_89  ))
// Xd_0__inst_mult_27_94  = SHARE((din_a[190] & (din_b[190] & (din_a[191] & din_b[189]))))

	.dataa(!din_a[190]),
	.datab(!din_b[190]),
	.datac(!din_a[191]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_89 ),
	.sharein(Xd_0__inst_mult_27_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_92 ),
	.cout(Xd_0__inst_mult_27_93 ),
	.shareout(Xd_0__inst_mult_27_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_30 (
// Equation(s):
// Xd_0__inst_mult_24_92  = SUM(( (!din_a[169] & (((din_a[170] & din_b[168])))) # (din_a[169] & (!din_b[169] $ (((!din_a[170]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_24_90  ) + ( Xd_0__inst_mult_24_89  ))
// Xd_0__inst_mult_24_93  = CARRY(( (!din_a[169] & (((din_a[170] & din_b[168])))) # (din_a[169] & (!din_b[169] $ (((!din_a[170]) # (!din_b[168]))))) ) + ( Xd_0__inst_mult_24_90  ) + ( Xd_0__inst_mult_24_89  ))
// Xd_0__inst_mult_24_94  = SHARE((din_a[169] & (din_b[169] & (din_a[170] & din_b[168]))))

	.dataa(!din_a[169]),
	.datab(!din_b[169]),
	.datac(!din_a[170]),
	.datad(!din_b[168]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_89 ),
	.sharein(Xd_0__inst_mult_24_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_92 ),
	.cout(Xd_0__inst_mult_24_93 ),
	.shareout(Xd_0__inst_mult_24_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_31 (
// Equation(s):
// Xd_0__inst_mult_25_96  = SUM(( (!din_a[176] & (((din_a[177] & din_b[175])))) # (din_a[176] & (!din_b[176] $ (((!din_a[177]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_25_94  ) + ( Xd_0__inst_mult_25_93  ))
// Xd_0__inst_mult_25_97  = CARRY(( (!din_a[176] & (((din_a[177] & din_b[175])))) # (din_a[176] & (!din_b[176] $ (((!din_a[177]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_25_94  ) + ( Xd_0__inst_mult_25_93  ))
// Xd_0__inst_mult_25_98  = SHARE((din_a[176] & (din_b[176] & (din_a[177] & din_b[175]))))

	.dataa(!din_a[176]),
	.datab(!din_b[176]),
	.datac(!din_a[177]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_93 ),
	.sharein(Xd_0__inst_mult_25_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_96 ),
	.cout(Xd_0__inst_mult_25_97 ),
	.shareout(Xd_0__inst_mult_25_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_31 (
// Equation(s):
// Xd_0__inst_mult_22_96  = SUM(( (!din_a[155] & (((din_a[156] & din_b[154])))) # (din_a[155] & (!din_b[155] $ (((!din_a[156]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_22_94  ) + ( Xd_0__inst_mult_22_93  ))
// Xd_0__inst_mult_22_97  = CARRY(( (!din_a[155] & (((din_a[156] & din_b[154])))) # (din_a[155] & (!din_b[155] $ (((!din_a[156]) # (!din_b[154]))))) ) + ( Xd_0__inst_mult_22_94  ) + ( Xd_0__inst_mult_22_93  ))
// Xd_0__inst_mult_22_98  = SHARE((din_a[155] & (din_b[155] & (din_a[156] & din_b[154]))))

	.dataa(!din_a[155]),
	.datab(!din_b[155]),
	.datac(!din_a[156]),
	.datad(!din_b[154]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_93 ),
	.sharein(Xd_0__inst_mult_22_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_96 ),
	.cout(Xd_0__inst_mult_22_97 ),
	.shareout(Xd_0__inst_mult_22_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_30 (
// Equation(s):
// Xd_0__inst_mult_23_92  = SUM(( (!din_a[162] & (((din_a[163] & din_b[161])))) # (din_a[162] & (!din_b[162] $ (((!din_a[163]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_23_90  ) + ( Xd_0__inst_mult_23_89  ))
// Xd_0__inst_mult_23_93  = CARRY(( (!din_a[162] & (((din_a[163] & din_b[161])))) # (din_a[162] & (!din_b[162] $ (((!din_a[163]) # (!din_b[161]))))) ) + ( Xd_0__inst_mult_23_90  ) + ( Xd_0__inst_mult_23_89  ))
// Xd_0__inst_mult_23_94  = SHARE((din_a[162] & (din_b[162] & (din_a[163] & din_b[161]))))

	.dataa(!din_a[162]),
	.datab(!din_b[162]),
	.datac(!din_a[163]),
	.datad(!din_b[161]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_89 ),
	.sharein(Xd_0__inst_mult_23_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_92 ),
	.cout(Xd_0__inst_mult_23_93 ),
	.shareout(Xd_0__inst_mult_23_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_30 (
// Equation(s):
// Xd_0__inst_mult_20_92  = SUM(( (!din_a[141] & (((din_a[142] & din_b[140])))) # (din_a[141] & (!din_b[141] $ (((!din_a[142]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_20_90  ) + ( Xd_0__inst_mult_20_89  ))
// Xd_0__inst_mult_20_93  = CARRY(( (!din_a[141] & (((din_a[142] & din_b[140])))) # (din_a[141] & (!din_b[141] $ (((!din_a[142]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_20_90  ) + ( Xd_0__inst_mult_20_89  ))
// Xd_0__inst_mult_20_94  = SHARE((din_a[141] & (din_b[141] & (din_a[142] & din_b[140]))))

	.dataa(!din_a[141]),
	.datab(!din_b[141]),
	.datac(!din_a[142]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_89 ),
	.sharein(Xd_0__inst_mult_20_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_92 ),
	.cout(Xd_0__inst_mult_20_93 ),
	.shareout(Xd_0__inst_mult_20_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_30 (
// Equation(s):
// Xd_0__inst_mult_21_92  = SUM(( (!din_a[148] & (((din_a[149] & din_b[147])))) # (din_a[148] & (!din_b[148] $ (((!din_a[149]) # (!din_b[147]))))) ) + ( Xd_0__inst_mult_21_90  ) + ( Xd_0__inst_mult_21_89  ))
// Xd_0__inst_mult_21_93  = CARRY(( (!din_a[148] & (((din_a[149] & din_b[147])))) # (din_a[148] & (!din_b[148] $ (((!din_a[149]) # (!din_b[147]))))) ) + ( Xd_0__inst_mult_21_90  ) + ( Xd_0__inst_mult_21_89  ))
// Xd_0__inst_mult_21_94  = SHARE((din_a[148] & (din_b[148] & (din_a[149] & din_b[147]))))

	.dataa(!din_a[148]),
	.datab(!din_b[148]),
	.datac(!din_a[149]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_89 ),
	.sharein(Xd_0__inst_mult_21_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_92 ),
	.cout(Xd_0__inst_mult_21_93 ),
	.shareout(Xd_0__inst_mult_21_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_30 (
// Equation(s):
// Xd_0__inst_mult_18_92  = SUM(( (!din_a[127] & (((din_a[128] & din_b[126])))) # (din_a[127] & (!din_b[127] $ (((!din_a[128]) # (!din_b[126]))))) ) + ( Xd_0__inst_mult_18_90  ) + ( Xd_0__inst_mult_18_89  ))
// Xd_0__inst_mult_18_93  = CARRY(( (!din_a[127] & (((din_a[128] & din_b[126])))) # (din_a[127] & (!din_b[127] $ (((!din_a[128]) # (!din_b[126]))))) ) + ( Xd_0__inst_mult_18_90  ) + ( Xd_0__inst_mult_18_89  ))
// Xd_0__inst_mult_18_94  = SHARE((din_a[127] & (din_b[127] & (din_a[128] & din_b[126]))))

	.dataa(!din_a[127]),
	.datab(!din_b[127]),
	.datac(!din_a[128]),
	.datad(!din_b[126]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_89 ),
	.sharein(Xd_0__inst_mult_18_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_92 ),
	.cout(Xd_0__inst_mult_18_93 ),
	.shareout(Xd_0__inst_mult_18_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_30 (
// Equation(s):
// Xd_0__inst_mult_19_92  = SUM(( (!din_a[134] & (((din_a[135] & din_b[133])))) # (din_a[134] & (!din_b[134] $ (((!din_a[135]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_19_90  ) + ( Xd_0__inst_mult_19_89  ))
// Xd_0__inst_mult_19_93  = CARRY(( (!din_a[134] & (((din_a[135] & din_b[133])))) # (din_a[134] & (!din_b[134] $ (((!din_a[135]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_19_90  ) + ( Xd_0__inst_mult_19_89  ))
// Xd_0__inst_mult_19_94  = SHARE((din_a[134] & (din_b[134] & (din_a[135] & din_b[133]))))

	.dataa(!din_a[134]),
	.datab(!din_b[134]),
	.datac(!din_a[135]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_89 ),
	.sharein(Xd_0__inst_mult_19_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_92 ),
	.cout(Xd_0__inst_mult_19_93 ),
	.shareout(Xd_0__inst_mult_19_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_30 (
// Equation(s):
// Xd_0__inst_mult_16_92  = SUM(( (!din_a[113] & (((din_a[114] & din_b[112])))) # (din_a[113] & (!din_b[113] $ (((!din_a[114]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_16_90  ) + ( Xd_0__inst_mult_16_89  ))
// Xd_0__inst_mult_16_93  = CARRY(( (!din_a[113] & (((din_a[114] & din_b[112])))) # (din_a[113] & (!din_b[113] $ (((!din_a[114]) # (!din_b[112]))))) ) + ( Xd_0__inst_mult_16_90  ) + ( Xd_0__inst_mult_16_89  ))
// Xd_0__inst_mult_16_94  = SHARE((din_a[113] & (din_b[113] & (din_a[114] & din_b[112]))))

	.dataa(!din_a[113]),
	.datab(!din_b[113]),
	.datac(!din_a[114]),
	.datad(!din_b[112]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_89 ),
	.sharein(Xd_0__inst_mult_16_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_92 ),
	.cout(Xd_0__inst_mult_16_93 ),
	.shareout(Xd_0__inst_mult_16_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_30 (
// Equation(s):
// Xd_0__inst_mult_17_92  = SUM(( (!din_a[120] & (((din_a[121] & din_b[119])))) # (din_a[120] & (!din_b[120] $ (((!din_a[121]) # (!din_b[119]))))) ) + ( Xd_0__inst_mult_17_90  ) + ( Xd_0__inst_mult_17_89  ))
// Xd_0__inst_mult_17_93  = CARRY(( (!din_a[120] & (((din_a[121] & din_b[119])))) # (din_a[120] & (!din_b[120] $ (((!din_a[121]) # (!din_b[119]))))) ) + ( Xd_0__inst_mult_17_90  ) + ( Xd_0__inst_mult_17_89  ))
// Xd_0__inst_mult_17_94  = SHARE((din_a[120] & (din_b[120] & (din_a[121] & din_b[119]))))

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(!din_a[121]),
	.datad(!din_b[119]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_89 ),
	.sharein(Xd_0__inst_mult_17_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_92 ),
	.cout(Xd_0__inst_mult_17_93 ),
	.shareout(Xd_0__inst_mult_17_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_30 (
// Equation(s):
// Xd_0__inst_mult_14_92  = SUM(( (!din_a[99] & (((din_a[100] & din_b[98])))) # (din_a[99] & (!din_b[99] $ (((!din_a[100]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_14_90  ) + ( Xd_0__inst_mult_14_89  ))
// Xd_0__inst_mult_14_93  = CARRY(( (!din_a[99] & (((din_a[100] & din_b[98])))) # (din_a[99] & (!din_b[99] $ (((!din_a[100]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_14_90  ) + ( Xd_0__inst_mult_14_89  ))
// Xd_0__inst_mult_14_94  = SHARE((din_a[99] & (din_b[99] & (din_a[100] & din_b[98]))))

	.dataa(!din_a[99]),
	.datab(!din_b[99]),
	.datac(!din_a[100]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_89 ),
	.sharein(Xd_0__inst_mult_14_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_92 ),
	.cout(Xd_0__inst_mult_14_93 ),
	.shareout(Xd_0__inst_mult_14_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_30 (
// Equation(s):
// Xd_0__inst_mult_15_92  = SUM(( (!din_a[106] & (((din_a[107] & din_b[105])))) # (din_a[106] & (!din_b[106] $ (((!din_a[107]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_15_90  ) + ( Xd_0__inst_mult_15_89  ))
// Xd_0__inst_mult_15_93  = CARRY(( (!din_a[106] & (((din_a[107] & din_b[105])))) # (din_a[106] & (!din_b[106] $ (((!din_a[107]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_15_90  ) + ( Xd_0__inst_mult_15_89  ))
// Xd_0__inst_mult_15_94  = SHARE((din_a[106] & (din_b[106] & (din_a[107] & din_b[105]))))

	.dataa(!din_a[106]),
	.datab(!din_b[106]),
	.datac(!din_a[107]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_89 ),
	.sharein(Xd_0__inst_mult_15_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_92 ),
	.cout(Xd_0__inst_mult_15_93 ),
	.shareout(Xd_0__inst_mult_15_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_30 (
// Equation(s):
// Xd_0__inst_mult_12_92  = SUM(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_12_90  ) + ( Xd_0__inst_mult_12_89  ))
// Xd_0__inst_mult_12_93  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_12_90  ) + ( Xd_0__inst_mult_12_89  ))
// Xd_0__inst_mult_12_94  = SHARE((din_a[85] & (din_b[85] & (din_a[86] & din_b[84]))))

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_89 ),
	.sharein(Xd_0__inst_mult_12_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_92 ),
	.cout(Xd_0__inst_mult_12_93 ),
	.shareout(Xd_0__inst_mult_12_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_30 (
// Equation(s):
// Xd_0__inst_mult_13_92  = SUM(( (!din_a[92] & (((din_a[93] & din_b[91])))) # (din_a[92] & (!din_b[92] $ (((!din_a[93]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_13_90  ) + ( Xd_0__inst_mult_13_89  ))
// Xd_0__inst_mult_13_93  = CARRY(( (!din_a[92] & (((din_a[93] & din_b[91])))) # (din_a[92] & (!din_b[92] $ (((!din_a[93]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_13_90  ) + ( Xd_0__inst_mult_13_89  ))
// Xd_0__inst_mult_13_94  = SHARE((din_a[92] & (din_b[92] & (din_a[93] & din_b[91]))))

	.dataa(!din_a[92]),
	.datab(!din_b[92]),
	.datac(!din_a[93]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_89 ),
	.sharein(Xd_0__inst_mult_13_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_92 ),
	.cout(Xd_0__inst_mult_13_93 ),
	.shareout(Xd_0__inst_mult_13_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_30 (
// Equation(s):
// Xd_0__inst_mult_10_92  = SUM(( (!din_a[71] & (((din_a[72] & din_b[70])))) # (din_a[71] & (!din_b[71] $ (((!din_a[72]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_10_90  ) + ( Xd_0__inst_mult_10_89  ))
// Xd_0__inst_mult_10_93  = CARRY(( (!din_a[71] & (((din_a[72] & din_b[70])))) # (din_a[71] & (!din_b[71] $ (((!din_a[72]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_10_90  ) + ( Xd_0__inst_mult_10_89  ))
// Xd_0__inst_mult_10_94  = SHARE((din_a[71] & (din_b[71] & (din_a[72] & din_b[70]))))

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(!din_a[72]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_89 ),
	.sharein(Xd_0__inst_mult_10_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_92 ),
	.cout(Xd_0__inst_mult_10_93 ),
	.shareout(Xd_0__inst_mult_10_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_30 (
// Equation(s):
// Xd_0__inst_mult_11_92  = SUM(( (!din_a[78] & (((din_a[79] & din_b[77])))) # (din_a[78] & (!din_b[78] $ (((!din_a[79]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_11_90  ) + ( Xd_0__inst_mult_11_89  ))
// Xd_0__inst_mult_11_93  = CARRY(( (!din_a[78] & (((din_a[79] & din_b[77])))) # (din_a[78] & (!din_b[78] $ (((!din_a[79]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_11_90  ) + ( Xd_0__inst_mult_11_89  ))
// Xd_0__inst_mult_11_94  = SHARE((din_a[78] & (din_b[78] & (din_a[79] & din_b[77]))))

	.dataa(!din_a[78]),
	.datab(!din_b[78]),
	.datac(!din_a[79]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_89 ),
	.sharein(Xd_0__inst_mult_11_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_92 ),
	.cout(Xd_0__inst_mult_11_93 ),
	.shareout(Xd_0__inst_mult_11_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_30 (
// Equation(s):
// Xd_0__inst_mult_8_92  = SUM(( (!din_a[57] & (((din_a[58] & din_b[56])))) # (din_a[57] & (!din_b[57] $ (((!din_a[58]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_8_90  ) + ( Xd_0__inst_mult_8_89  ))
// Xd_0__inst_mult_8_93  = CARRY(( (!din_a[57] & (((din_a[58] & din_b[56])))) # (din_a[57] & (!din_b[57] $ (((!din_a[58]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_8_90  ) + ( Xd_0__inst_mult_8_89  ))
// Xd_0__inst_mult_8_94  = SHARE((din_a[57] & (din_b[57] & (din_a[58] & din_b[56]))))

	.dataa(!din_a[57]),
	.datab(!din_b[57]),
	.datac(!din_a[58]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_89 ),
	.sharein(Xd_0__inst_mult_8_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_92 ),
	.cout(Xd_0__inst_mult_8_93 ),
	.shareout(Xd_0__inst_mult_8_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_30 (
// Equation(s):
// Xd_0__inst_mult_9_92  = SUM(( (!din_a[64] & (((din_a[65] & din_b[63])))) # (din_a[64] & (!din_b[64] $ (((!din_a[65]) # (!din_b[63]))))) ) + ( Xd_0__inst_mult_9_90  ) + ( Xd_0__inst_mult_9_89  ))
// Xd_0__inst_mult_9_93  = CARRY(( (!din_a[64] & (((din_a[65] & din_b[63])))) # (din_a[64] & (!din_b[64] $ (((!din_a[65]) # (!din_b[63]))))) ) + ( Xd_0__inst_mult_9_90  ) + ( Xd_0__inst_mult_9_89  ))
// Xd_0__inst_mult_9_94  = SHARE((din_a[64] & (din_b[64] & (din_a[65] & din_b[63]))))

	.dataa(!din_a[64]),
	.datab(!din_b[64]),
	.datac(!din_a[65]),
	.datad(!din_b[63]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_89 ),
	.sharein(Xd_0__inst_mult_9_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_92 ),
	.cout(Xd_0__inst_mult_9_93 ),
	.shareout(Xd_0__inst_mult_9_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_30 (
// Equation(s):
// Xd_0__inst_mult_6_92  = SUM(( (!din_a[43] & (((din_a[44] & din_b[42])))) # (din_a[43] & (!din_b[43] $ (((!din_a[44]) # (!din_b[42]))))) ) + ( Xd_0__inst_mult_6_90  ) + ( Xd_0__inst_mult_6_89  ))
// Xd_0__inst_mult_6_93  = CARRY(( (!din_a[43] & (((din_a[44] & din_b[42])))) # (din_a[43] & (!din_b[43] $ (((!din_a[44]) # (!din_b[42]))))) ) + ( Xd_0__inst_mult_6_90  ) + ( Xd_0__inst_mult_6_89  ))
// Xd_0__inst_mult_6_94  = SHARE((din_a[43] & (din_b[43] & (din_a[44] & din_b[42]))))

	.dataa(!din_a[43]),
	.datab(!din_b[43]),
	.datac(!din_a[44]),
	.datad(!din_b[42]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_89 ),
	.sharein(Xd_0__inst_mult_6_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_92 ),
	.cout(Xd_0__inst_mult_6_93 ),
	.shareout(Xd_0__inst_mult_6_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_30 (
// Equation(s):
// Xd_0__inst_mult_7_92  = SUM(( (!din_a[50] & (((din_a[51] & din_b[49])))) # (din_a[50] & (!din_b[50] $ (((!din_a[51]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_7_90  ) + ( Xd_0__inst_mult_7_89  ))
// Xd_0__inst_mult_7_93  = CARRY(( (!din_a[50] & (((din_a[51] & din_b[49])))) # (din_a[50] & (!din_b[50] $ (((!din_a[51]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_7_90  ) + ( Xd_0__inst_mult_7_89  ))
// Xd_0__inst_mult_7_94  = SHARE((din_a[50] & (din_b[50] & (din_a[51] & din_b[49]))))

	.dataa(!din_a[50]),
	.datab(!din_b[50]),
	.datac(!din_a[51]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_89 ),
	.sharein(Xd_0__inst_mult_7_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_92 ),
	.cout(Xd_0__inst_mult_7_93 ),
	.shareout(Xd_0__inst_mult_7_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_30 (
// Equation(s):
// Xd_0__inst_mult_4_92  = SUM(( (!din_a[29] & (((din_a[30] & din_b[28])))) # (din_a[29] & (!din_b[29] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_4_90  ) + ( Xd_0__inst_mult_4_89  ))
// Xd_0__inst_mult_4_93  = CARRY(( (!din_a[29] & (((din_a[30] & din_b[28])))) # (din_a[29] & (!din_b[29] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_4_90  ) + ( Xd_0__inst_mult_4_89  ))
// Xd_0__inst_mult_4_94  = SHARE((din_a[29] & (din_b[29] & (din_a[30] & din_b[28]))))

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(!din_a[30]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_89 ),
	.sharein(Xd_0__inst_mult_4_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_92 ),
	.cout(Xd_0__inst_mult_4_93 ),
	.shareout(Xd_0__inst_mult_4_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_30 (
// Equation(s):
// Xd_0__inst_mult_5_92  = SUM(( (!din_a[36] & (((din_a[37] & din_b[35])))) # (din_a[36] & (!din_b[36] $ (((!din_a[37]) # (!din_b[35]))))) ) + ( Xd_0__inst_mult_5_90  ) + ( Xd_0__inst_mult_5_89  ))
// Xd_0__inst_mult_5_93  = CARRY(( (!din_a[36] & (((din_a[37] & din_b[35])))) # (din_a[36] & (!din_b[36] $ (((!din_a[37]) # (!din_b[35]))))) ) + ( Xd_0__inst_mult_5_90  ) + ( Xd_0__inst_mult_5_89  ))
// Xd_0__inst_mult_5_94  = SHARE((din_a[36] & (din_b[36] & (din_a[37] & din_b[35]))))

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(!din_a[37]),
	.datad(!din_b[35]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_89 ),
	.sharein(Xd_0__inst_mult_5_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_92 ),
	.cout(Xd_0__inst_mult_5_93 ),
	.shareout(Xd_0__inst_mult_5_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_30 (
// Equation(s):
// Xd_0__inst_mult_2_92  = SUM(( (!din_a[15] & (((din_a[16] & din_b[14])))) # (din_a[15] & (!din_b[15] $ (((!din_a[16]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_90  ) + ( Xd_0__inst_mult_2_89  ))
// Xd_0__inst_mult_2_93  = CARRY(( (!din_a[15] & (((din_a[16] & din_b[14])))) # (din_a[15] & (!din_b[15] $ (((!din_a[16]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_90  ) + ( Xd_0__inst_mult_2_89  ))
// Xd_0__inst_mult_2_94  = SHARE((din_a[15] & (din_b[15] & (din_a[16] & din_b[14]))))

	.dataa(!din_a[15]),
	.datab(!din_b[15]),
	.datac(!din_a[16]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_89 ),
	.sharein(Xd_0__inst_mult_2_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_92 ),
	.cout(Xd_0__inst_mult_2_93 ),
	.shareout(Xd_0__inst_mult_2_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_30 (
// Equation(s):
// Xd_0__inst_mult_3_92  = SUM(( (!din_a[22] & (((din_a[23] & din_b[21])))) # (din_a[22] & (!din_b[22] $ (((!din_a[23]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_3_90  ) + ( Xd_0__inst_mult_3_89  ))
// Xd_0__inst_mult_3_93  = CARRY(( (!din_a[22] & (((din_a[23] & din_b[21])))) # (din_a[22] & (!din_b[22] $ (((!din_a[23]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_3_90  ) + ( Xd_0__inst_mult_3_89  ))
// Xd_0__inst_mult_3_94  = SHARE((din_a[22] & (din_b[22] & (din_a[23] & din_b[21]))))

	.dataa(!din_a[22]),
	.datab(!din_b[22]),
	.datac(!din_a[23]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_89 ),
	.sharein(Xd_0__inst_mult_3_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_92 ),
	.cout(Xd_0__inst_mult_3_93 ),
	.shareout(Xd_0__inst_mult_3_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_30 (
// Equation(s):
// Xd_0__inst_mult_0_92  = SUM(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_90  ) + ( Xd_0__inst_mult_0_89  ))
// Xd_0__inst_mult_0_93  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_90  ) + ( Xd_0__inst_mult_0_89  ))
// Xd_0__inst_mult_0_94  = SHARE((din_a[1] & (din_b[1] & (din_a[2] & din_b[0]))))

	.dataa(!din_a[1]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_89 ),
	.sharein(Xd_0__inst_mult_0_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_92 ),
	.cout(Xd_0__inst_mult_0_93 ),
	.shareout(Xd_0__inst_mult_0_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_30 (
// Equation(s):
// Xd_0__inst_mult_1_92  = SUM(( (!din_a[8] & (((din_a[9] & din_b[7])))) # (din_a[8] & (!din_b[8] $ (((!din_a[9]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_90  ) + ( Xd_0__inst_mult_1_89  ))
// Xd_0__inst_mult_1_93  = CARRY(( (!din_a[8] & (((din_a[9] & din_b[7])))) # (din_a[8] & (!din_b[8] $ (((!din_a[9]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_90  ) + ( Xd_0__inst_mult_1_89  ))
// Xd_0__inst_mult_1_94  = SHARE((din_a[8] & (din_b[8] & (din_a[9] & din_b[7]))))

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(!din_a[9]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_89 ),
	.sharein(Xd_0__inst_mult_1_90 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_92 ),
	.cout(Xd_0__inst_mult_1_93 ),
	.shareout(Xd_0__inst_mult_1_94 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_31 (
// Equation(s):
// Xd_0__inst_mult_28_97  = CARRY(( GND ) + ( Xd_0__inst_mult_0_82  ) + ( Xd_0__inst_mult_0_81  ))
// Xd_0__inst_mult_28_98  = SHARE((Xd_0__inst_mult_28_0_q  & Xd_0__inst_mult_28_1_q ))

	.dataa(!Xd_0__inst_mult_28_0_q ),
	.datab(!Xd_0__inst_mult_28_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_81 ),
	.sharein(Xd_0__inst_mult_0_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_97 ),
	.shareout(Xd_0__inst_mult_28_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_31 (
// Equation(s):
// Xd_0__inst_mult_29_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_29_98  = SHARE((Xd_0__inst_mult_29_0_q  & Xd_0__inst_mult_29_1_q ))

	.dataa(!Xd_0__inst_mult_29_0_q ),
	.datab(!Xd_0__inst_mult_29_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_97 ),
	.shareout(Xd_0__inst_mult_29_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_31 (
// Equation(s):
// Xd_0__inst_mult_26_97  = CARRY(( GND ) + ( Xd_0__inst_mult_4_82  ) + ( Xd_0__inst_mult_4_81  ))
// Xd_0__inst_mult_26_98  = SHARE((Xd_0__inst_mult_26_0_q  & Xd_0__inst_mult_26_1_q ))

	.dataa(!Xd_0__inst_mult_26_0_q ),
	.datab(!Xd_0__inst_mult_26_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_81 ),
	.sharein(Xd_0__inst_mult_4_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_97 ),
	.shareout(Xd_0__inst_mult_26_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_31 (
// Equation(s):
// Xd_0__inst_mult_27_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_27_98  = SHARE((Xd_0__inst_mult_27_0_q  & Xd_0__inst_mult_27_1_q ))

	.dataa(!Xd_0__inst_mult_27_0_q ),
	.datab(!Xd_0__inst_mult_27_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_97 ),
	.shareout(Xd_0__inst_mult_27_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_31 (
// Equation(s):
// Xd_0__inst_mult_24_97  = CARRY(( GND ) + ( Xd_0__inst_mult_27_82  ) + ( Xd_0__inst_mult_27_81  ))
// Xd_0__inst_mult_24_98  = SHARE((Xd_0__inst_mult_24_0_q  & Xd_0__inst_mult_24_1_q ))

	.dataa(!Xd_0__inst_mult_24_0_q ),
	.datab(!Xd_0__inst_mult_24_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_81 ),
	.sharein(Xd_0__inst_mult_27_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_97 ),
	.shareout(Xd_0__inst_mult_24_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_32 (
// Equation(s):
// Xd_0__inst_mult_25_101  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_25_102  = SHARE((Xd_0__inst_mult_25_0_q  & Xd_0__inst_mult_25_1_q ))

	.dataa(!Xd_0__inst_mult_25_0_q ),
	.datab(!Xd_0__inst_mult_25_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_101 ),
	.shareout(Xd_0__inst_mult_25_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_32 (
// Equation(s):
// Xd_0__inst_mult_22_101  = CARRY(( GND ) + ( Xd_0__inst_mult_19_82  ) + ( Xd_0__inst_mult_19_81  ))
// Xd_0__inst_mult_22_102  = SHARE((Xd_0__inst_mult_22_0_q  & Xd_0__inst_mult_22_1_q ))

	.dataa(!Xd_0__inst_mult_22_0_q ),
	.datab(!Xd_0__inst_mult_22_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_81 ),
	.sharein(Xd_0__inst_mult_19_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_101 ),
	.shareout(Xd_0__inst_mult_22_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_31 (
// Equation(s):
// Xd_0__inst_mult_23_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_23_98  = SHARE((Xd_0__inst_mult_23_0_q  & Xd_0__inst_mult_23_1_q ))

	.dataa(!Xd_0__inst_mult_23_0_q ),
	.datab(!Xd_0__inst_mult_23_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_97 ),
	.shareout(Xd_0__inst_mult_23_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_31 (
// Equation(s):
// Xd_0__inst_mult_20_97  = CARRY(( GND ) + ( Xd_0__inst_mult_23_82  ) + ( Xd_0__inst_mult_23_81  ))
// Xd_0__inst_mult_20_98  = SHARE((Xd_0__inst_mult_20_0_q  & Xd_0__inst_mult_20_1_q ))

	.dataa(!Xd_0__inst_mult_20_0_q ),
	.datab(!Xd_0__inst_mult_20_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_81 ),
	.sharein(Xd_0__inst_mult_23_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_97 ),
	.shareout(Xd_0__inst_mult_20_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_31 (
// Equation(s):
// Xd_0__inst_mult_21_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_21_98  = SHARE((Xd_0__inst_mult_21_0_q  & Xd_0__inst_mult_21_1_q ))

	.dataa(!Xd_0__inst_mult_21_0_q ),
	.datab(!Xd_0__inst_mult_21_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_97 ),
	.shareout(Xd_0__inst_mult_21_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_31 (
// Equation(s):
// Xd_0__inst_mult_18_97  = CARRY(( GND ) + ( Xd_0__inst_mult_6_82  ) + ( Xd_0__inst_mult_6_81  ))
// Xd_0__inst_mult_18_98  = SHARE((Xd_0__inst_mult_18_0_q  & Xd_0__inst_mult_18_1_q ))

	.dataa(!Xd_0__inst_mult_18_0_q ),
	.datab(!Xd_0__inst_mult_18_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_81 ),
	.sharein(Xd_0__inst_mult_6_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_97 ),
	.shareout(Xd_0__inst_mult_18_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_31 (
// Equation(s):
// Xd_0__inst_mult_19_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_19_98  = SHARE((Xd_0__inst_mult_19_0_q  & Xd_0__inst_mult_19_1_q ))

	.dataa(!Xd_0__inst_mult_19_0_q ),
	.datab(!Xd_0__inst_mult_19_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_97 ),
	.shareout(Xd_0__inst_mult_19_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_32 (
// Equation(s):
// Xd_0__inst_mult_30_100  = SUM(( (!din_a[212] & (((din_a[211] & din_b[212])))) # (din_a[212] & (!din_b[211] $ (((!din_a[211]) # (!din_b[212]))))) ) + ( Xd_0__inst_mult_30_94  ) + ( Xd_0__inst_mult_30_93  ))
// Xd_0__inst_mult_30_101  = CARRY(( (!din_a[212] & (((din_a[211] & din_b[212])))) # (din_a[212] & (!din_b[211] $ (((!din_a[211]) # (!din_b[212]))))) ) + ( Xd_0__inst_mult_30_94  ) + ( Xd_0__inst_mult_30_93  ))
// Xd_0__inst_mult_30_102  = SHARE((din_a[212] & (din_b[211] & (din_a[211] & din_b[212]))))

	.dataa(!din_a[212]),
	.datab(!din_b[211]),
	.datac(!din_a[211]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_93 ),
	.sharein(Xd_0__inst_mult_30_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_100 ),
	.cout(Xd_0__inst_mult_30_101 ),
	.shareout(Xd_0__inst_mult_30_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_32 (
// Equation(s):
// Xd_0__inst_mult_31_100  = SUM(( (!din_a[219] & (((din_a[218] & din_b[219])))) # (din_a[219] & (!din_b[218] $ (((!din_a[218]) # (!din_b[219]))))) ) + ( Xd_0__inst_mult_31_94  ) + ( Xd_0__inst_mult_31_93  ))
// Xd_0__inst_mult_31_101  = CARRY(( (!din_a[219] & (((din_a[218] & din_b[219])))) # (din_a[219] & (!din_b[218] $ (((!din_a[218]) # (!din_b[219]))))) ) + ( Xd_0__inst_mult_31_94  ) + ( Xd_0__inst_mult_31_93  ))
// Xd_0__inst_mult_31_102  = SHARE((din_a[219] & (din_b[218] & (din_a[218] & din_b[219]))))

	.dataa(!din_a[219]),
	.datab(!din_b[218]),
	.datac(!din_a[218]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_93 ),
	.sharein(Xd_0__inst_mult_31_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_100 ),
	.cout(Xd_0__inst_mult_31_101 ),
	.shareout(Xd_0__inst_mult_31_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_31 (
// Equation(s):
// Xd_0__inst_mult_16_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_16_98  = SHARE((Xd_0__inst_mult_16_0_q  & Xd_0__inst_mult_16_1_q ))

	.dataa(!Xd_0__inst_mult_16_0_q ),
	.datab(!Xd_0__inst_mult_16_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_97 ),
	.shareout(Xd_0__inst_mult_16_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_31 (
// Equation(s):
// Xd_0__inst_mult_17_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_17_98  = SHARE((Xd_0__inst_mult_17_0_q  & Xd_0__inst_mult_17_1_q ))

	.dataa(!Xd_0__inst_mult_17_0_q ),
	.datab(!Xd_0__inst_mult_17_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_97 ),
	.shareout(Xd_0__inst_mult_17_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_31 (
// Equation(s):
// Xd_0__inst_mult_14_97  = CARRY(( GND ) + ( Xd_0__inst_mult_8_82  ) + ( Xd_0__inst_mult_8_81  ))
// Xd_0__inst_mult_14_98  = SHARE((Xd_0__inst_mult_14_0_q  & Xd_0__inst_mult_14_1_q ))

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_81 ),
	.sharein(Xd_0__inst_mult_8_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_97 ),
	.shareout(Xd_0__inst_mult_14_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_31 (
// Equation(s):
// Xd_0__inst_mult_15_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_98  = SHARE((Xd_0__inst_mult_15_0_q  & Xd_0__inst_mult_15_1_q ))

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_97 ),
	.shareout(Xd_0__inst_mult_15_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_31 (
// Equation(s):
// Xd_0__inst_mult_12_97  = CARRY(( GND ) + ( Xd_0__inst_mult_15_82  ) + ( Xd_0__inst_mult_15_81  ))
// Xd_0__inst_mult_12_98  = SHARE((Xd_0__inst_mult_12_0_q  & Xd_0__inst_mult_12_1_q ))

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_81 ),
	.sharein(Xd_0__inst_mult_15_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_97 ),
	.shareout(Xd_0__inst_mult_12_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_31 (
// Equation(s):
// Xd_0__inst_mult_13_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_98  = SHARE((Xd_0__inst_mult_13_0_q  & Xd_0__inst_mult_13_1_q ))

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_97 ),
	.shareout(Xd_0__inst_mult_13_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_31 (
// Equation(s):
// Xd_0__inst_mult_10_97  = CARRY(( GND ) + ( Xd_0__inst_mult_16_82  ) + ( Xd_0__inst_mult_16_81  ))
// Xd_0__inst_mult_10_98  = SHARE((Xd_0__inst_mult_10_0_q  & Xd_0__inst_mult_10_1_q ))

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_81 ),
	.sharein(Xd_0__inst_mult_16_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_97 ),
	.shareout(Xd_0__inst_mult_10_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_31 (
// Equation(s):
// Xd_0__inst_mult_11_97  = CARRY(( GND ) + ( Xd_0__inst_mult_13_82  ) + ( Xd_0__inst_mult_13_81  ))
// Xd_0__inst_mult_11_98  = SHARE((Xd_0__inst_mult_11_0_q  & Xd_0__inst_mult_11_1_q ))

	.dataa(!Xd_0__inst_mult_11_0_q ),
	.datab(!Xd_0__inst_mult_11_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_81 ),
	.sharein(Xd_0__inst_mult_13_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_97 ),
	.shareout(Xd_0__inst_mult_11_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_31 (
// Equation(s):
// Xd_0__inst_mult_8_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_98  = SHARE((Xd_0__inst_mult_8_0_q  & Xd_0__inst_mult_8_1_q ))

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_97 ),
	.shareout(Xd_0__inst_mult_8_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_31 (
// Equation(s):
// Xd_0__inst_mult_9_97  = CARRY(( GND ) + ( Xd_0__inst_mult_17_82  ) + ( Xd_0__inst_mult_17_81  ))
// Xd_0__inst_mult_9_98  = SHARE((Xd_0__inst_mult_9_0_q  & Xd_0__inst_mult_9_1_q ))

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_81 ),
	.sharein(Xd_0__inst_mult_17_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_97 ),
	.shareout(Xd_0__inst_mult_9_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_31 (
// Equation(s):
// Xd_0__inst_mult_6_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_98  = SHARE((Xd_0__inst_mult_6_0_q  & Xd_0__inst_mult_6_1_q ))

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_97 ),
	.shareout(Xd_0__inst_mult_6_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_31 (
// Equation(s):
// Xd_0__inst_mult_7_97  = CARRY(( GND ) + ( Xd_0__inst_mult_21_82  ) + ( Xd_0__inst_mult_21_81  ))
// Xd_0__inst_mult_7_98  = SHARE((Xd_0__inst_mult_7_0_q  & Xd_0__inst_mult_7_1_q ))

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_81 ),
	.sharein(Xd_0__inst_mult_21_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_97 ),
	.shareout(Xd_0__inst_mult_7_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_31 (
// Equation(s):
// Xd_0__inst_mult_4_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_98  = SHARE((Xd_0__inst_mult_4_0_q  & Xd_0__inst_mult_4_1_q ))

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_97 ),
	.shareout(Xd_0__inst_mult_4_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_31 (
// Equation(s):
// Xd_0__inst_mult_5_97  = CARRY(( GND ) + ( Xd_0__inst_mult_25_82  ) + ( Xd_0__inst_mult_25_81  ))
// Xd_0__inst_mult_5_98  = SHARE((Xd_0__inst_mult_5_0_q  & Xd_0__inst_mult_5_1_q ))

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_81 ),
	.sharein(Xd_0__inst_mult_25_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_97 ),
	.shareout(Xd_0__inst_mult_5_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_31 (
// Equation(s):
// Xd_0__inst_mult_2_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_98  = SHARE((Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_1_q ))

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_97 ),
	.shareout(Xd_0__inst_mult_2_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_31 (
// Equation(s):
// Xd_0__inst_mult_3_97  = CARRY(( GND ) + ( Xd_0__inst_mult_29_82  ) + ( Xd_0__inst_mult_29_81  ))
// Xd_0__inst_mult_3_98  = SHARE((Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_1_q ))

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_81 ),
	.sharein(Xd_0__inst_mult_29_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_97 ),
	.shareout(Xd_0__inst_mult_3_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_31 (
// Equation(s):
// Xd_0__inst_mult_0_97  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_98  = SHARE((Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_1_q ))

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_97 ),
	.shareout(Xd_0__inst_mult_0_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_31 (
// Equation(s):
// Xd_0__inst_mult_1_97  = CARRY(( GND ) + ( Xd_0__inst_mult_2_82  ) + ( Xd_0__inst_mult_2_81  ))
// Xd_0__inst_mult_1_98  = SHARE((Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_1_q ))

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_81 ),
	.sharein(Xd_0__inst_mult_2_82 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_97 ),
	.shareout(Xd_0__inst_mult_1_98 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_33 (
// Equation(s):
// Xd_0__inst_mult_30_104  = SUM(( (din_a[213] & din_b[211]) ) + ( Xd_0__inst_mult_30_102  ) + ( Xd_0__inst_mult_30_101  ))
// Xd_0__inst_mult_30_105  = CARRY(( (din_a[213] & din_b[211]) ) + ( Xd_0__inst_mult_30_102  ) + ( Xd_0__inst_mult_30_101  ))
// Xd_0__inst_mult_30_106  = SHARE((din_a[213] & din_b[212]))

	.dataa(!din_a[213]),
	.datab(!din_b[211]),
	.datac(!din_b[212]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_101 ),
	.sharein(Xd_0__inst_mult_30_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_104 ),
	.cout(Xd_0__inst_mult_30_105 ),
	.shareout(Xd_0__inst_mult_30_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_34 (
// Equation(s):
// Xd_0__inst_mult_30_108  = SUM(( (din_a[210] & din_b[214]) ) + ( Xd_0__inst_mult_30_158  ) + ( Xd_0__inst_mult_30_157  ))
// Xd_0__inst_mult_30_109  = CARRY(( (din_a[210] & din_b[214]) ) + ( Xd_0__inst_mult_30_158  ) + ( Xd_0__inst_mult_30_157  ))
// Xd_0__inst_mult_30_110  = SHARE((din_a[212] & din_b[213]))

	.dataa(!din_a[210]),
	.datab(!din_b[214]),
	.datac(!din_a[212]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_157 ),
	.sharein(Xd_0__inst_mult_30_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_108 ),
	.cout(Xd_0__inst_mult_30_109 ),
	.shareout(Xd_0__inst_mult_30_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_33 (
// Equation(s):
// Xd_0__inst_mult_31_104  = SUM(( (din_a[220] & din_b[218]) ) + ( Xd_0__inst_mult_31_102  ) + ( Xd_0__inst_mult_31_101  ))
// Xd_0__inst_mult_31_105  = CARRY(( (din_a[220] & din_b[218]) ) + ( Xd_0__inst_mult_31_102  ) + ( Xd_0__inst_mult_31_101  ))
// Xd_0__inst_mult_31_106  = SHARE((din_a[220] & din_b[219]))

	.dataa(!din_a[220]),
	.datab(!din_b[218]),
	.datac(!din_b[219]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_101 ),
	.sharein(Xd_0__inst_mult_31_102 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_104 ),
	.cout(Xd_0__inst_mult_31_105 ),
	.shareout(Xd_0__inst_mult_31_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_34 (
// Equation(s):
// Xd_0__inst_mult_31_108  = SUM(( (din_a[217] & din_b[221]) ) + ( Xd_0__inst_mult_31_158  ) + ( Xd_0__inst_mult_31_157  ))
// Xd_0__inst_mult_31_109  = CARRY(( (din_a[217] & din_b[221]) ) + ( Xd_0__inst_mult_31_158  ) + ( Xd_0__inst_mult_31_157  ))
// Xd_0__inst_mult_31_110  = SHARE((din_a[219] & din_b[220]))

	.dataa(!din_a[217]),
	.datab(!din_b[221]),
	.datac(!din_a[219]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_157 ),
	.sharein(Xd_0__inst_mult_31_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_108 ),
	.cout(Xd_0__inst_mult_31_109 ),
	.shareout(Xd_0__inst_mult_31_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_35 (
// Equation(s):
// Xd_0__inst_mult_30_112  = SUM(( (!din_a[215] & (((din_a[214] & din_b[211])))) # (din_a[215] & (!din_b[210] $ (((!din_a[214]) # (!din_b[211]))))) ) + ( Xd_0__inst_mult_30_106  ) + ( Xd_0__inst_mult_30_105  ))
// Xd_0__inst_mult_30_113  = CARRY(( (!din_a[215] & (((din_a[214] & din_b[211])))) # (din_a[215] & (!din_b[210] $ (((!din_a[214]) # (!din_b[211]))))) ) + ( Xd_0__inst_mult_30_106  ) + ( Xd_0__inst_mult_30_105  ))
// Xd_0__inst_mult_30_114  = SHARE((din_a[215] & (din_b[210] & (din_a[214] & din_b[211]))))

	.dataa(!din_a[215]),
	.datab(!din_b[210]),
	.datac(!din_a[214]),
	.datad(!din_b[211]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_105 ),
	.sharein(Xd_0__inst_mult_30_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_112 ),
	.cout(Xd_0__inst_mult_30_113 ),
	.shareout(Xd_0__inst_mult_30_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_36 (
// Equation(s):
// Xd_0__inst_mult_30_116  = SUM(( (!din_a[211] & (((din_a[210] & din_b[215])))) # (din_a[211] & (!din_b[214] $ (((!din_a[210]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_110  ) + ( Xd_0__inst_mult_30_109  ))
// Xd_0__inst_mult_30_117  = CARRY(( (!din_a[211] & (((din_a[210] & din_b[215])))) # (din_a[211] & (!din_b[214] $ (((!din_a[210]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_110  ) + ( Xd_0__inst_mult_30_109  ))
// Xd_0__inst_mult_30_118  = SHARE((din_a[211] & (din_b[214] & (din_a[210] & din_b[215]))))

	.dataa(!din_a[211]),
	.datab(!din_b[214]),
	.datac(!din_a[210]),
	.datad(!din_b[215]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_109 ),
	.sharein(Xd_0__inst_mult_30_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_116 ),
	.cout(Xd_0__inst_mult_30_117 ),
	.shareout(Xd_0__inst_mult_30_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_35 (
// Equation(s):
// Xd_0__inst_mult_31_112  = SUM(( (!din_a[222] & (((din_a[221] & din_b[218])))) # (din_a[222] & (!din_b[217] $ (((!din_a[221]) # (!din_b[218]))))) ) + ( Xd_0__inst_mult_31_106  ) + ( Xd_0__inst_mult_31_105  ))
// Xd_0__inst_mult_31_113  = CARRY(( (!din_a[222] & (((din_a[221] & din_b[218])))) # (din_a[222] & (!din_b[217] $ (((!din_a[221]) # (!din_b[218]))))) ) + ( Xd_0__inst_mult_31_106  ) + ( Xd_0__inst_mult_31_105  ))
// Xd_0__inst_mult_31_114  = SHARE((din_a[222] & (din_b[217] & (din_a[221] & din_b[218]))))

	.dataa(!din_a[222]),
	.datab(!din_b[217]),
	.datac(!din_a[221]),
	.datad(!din_b[218]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_105 ),
	.sharein(Xd_0__inst_mult_31_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_112 ),
	.cout(Xd_0__inst_mult_31_113 ),
	.shareout(Xd_0__inst_mult_31_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_36 (
// Equation(s):
// Xd_0__inst_mult_31_116  = SUM(( (!din_a[218] & (((din_a[217] & din_b[222])))) # (din_a[218] & (!din_b[221] $ (((!din_a[217]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_110  ) + ( Xd_0__inst_mult_31_109  ))
// Xd_0__inst_mult_31_117  = CARRY(( (!din_a[218] & (((din_a[217] & din_b[222])))) # (din_a[218] & (!din_b[221] $ (((!din_a[217]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_110  ) + ( Xd_0__inst_mult_31_109  ))
// Xd_0__inst_mult_31_118  = SHARE((din_a[218] & (din_b[221] & (din_a[217] & din_b[222]))))

	.dataa(!din_a[218]),
	.datab(!din_b[221]),
	.datac(!din_a[217]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_109 ),
	.sharein(Xd_0__inst_mult_31_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_116 ),
	.cout(Xd_0__inst_mult_31_117 ),
	.shareout(Xd_0__inst_mult_31_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_37 (
// Equation(s):
// Xd_0__inst_mult_30_120  = SUM(( (!din_a[215] & (((din_a[214] & din_b[212])))) # (din_a[215] & (!din_b[211] $ (((!din_a[214]) # (!din_b[212]))))) ) + ( Xd_0__inst_mult_30_114  ) + ( Xd_0__inst_mult_30_113  ))
// Xd_0__inst_mult_30_121  = CARRY(( (!din_a[215] & (((din_a[214] & din_b[212])))) # (din_a[215] & (!din_b[211] $ (((!din_a[214]) # (!din_b[212]))))) ) + ( Xd_0__inst_mult_30_114  ) + ( Xd_0__inst_mult_30_113  ))
// Xd_0__inst_mult_30_122  = SHARE((din_a[215] & (din_b[211] & (din_a[214] & din_b[212]))))

	.dataa(!din_a[215]),
	.datab(!din_b[211]),
	.datac(!din_a[214]),
	.datad(!din_b[212]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_113 ),
	.sharein(Xd_0__inst_mult_30_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_120 ),
	.cout(Xd_0__inst_mult_30_121 ),
	.shareout(Xd_0__inst_mult_30_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_38 (
// Equation(s):
// Xd_0__inst_mult_30_124  = SUM(( (!din_a[212] & (((din_a[211] & din_b[215])))) # (din_a[212] & (!din_b[214] $ (((!din_a[211]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_118  ) + ( Xd_0__inst_mult_30_117  ))
// Xd_0__inst_mult_30_125  = CARRY(( (!din_a[212] & (((din_a[211] & din_b[215])))) # (din_a[212] & (!din_b[214] $ (((!din_a[211]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_118  ) + ( Xd_0__inst_mult_30_117  ))
// Xd_0__inst_mult_30_126  = SHARE((din_a[212] & (din_b[214] & (din_a[211] & din_b[215]))))

	.dataa(!din_a[212]),
	.datab(!din_b[214]),
	.datac(!din_a[211]),
	.datad(!din_b[215]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_117 ),
	.sharein(Xd_0__inst_mult_30_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_124 ),
	.cout(Xd_0__inst_mult_30_125 ),
	.shareout(Xd_0__inst_mult_30_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_37 (
// Equation(s):
// Xd_0__inst_mult_31_120  = SUM(( (!din_a[222] & (((din_a[221] & din_b[219])))) # (din_a[222] & (!din_b[218] $ (((!din_a[221]) # (!din_b[219]))))) ) + ( Xd_0__inst_mult_31_114  ) + ( Xd_0__inst_mult_31_113  ))
// Xd_0__inst_mult_31_121  = CARRY(( (!din_a[222] & (((din_a[221] & din_b[219])))) # (din_a[222] & (!din_b[218] $ (((!din_a[221]) # (!din_b[219]))))) ) + ( Xd_0__inst_mult_31_114  ) + ( Xd_0__inst_mult_31_113  ))
// Xd_0__inst_mult_31_122  = SHARE((din_a[222] & (din_b[218] & (din_a[221] & din_b[219]))))

	.dataa(!din_a[222]),
	.datab(!din_b[218]),
	.datac(!din_a[221]),
	.datad(!din_b[219]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_113 ),
	.sharein(Xd_0__inst_mult_31_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_120 ),
	.cout(Xd_0__inst_mult_31_121 ),
	.shareout(Xd_0__inst_mult_31_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_38 (
// Equation(s):
// Xd_0__inst_mult_31_124  = SUM(( (!din_a[219] & (((din_a[218] & din_b[222])))) # (din_a[219] & (!din_b[221] $ (((!din_a[218]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_118  ) + ( Xd_0__inst_mult_31_117  ))
// Xd_0__inst_mult_31_125  = CARRY(( (!din_a[219] & (((din_a[218] & din_b[222])))) # (din_a[219] & (!din_b[221] $ (((!din_a[218]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_118  ) + ( Xd_0__inst_mult_31_117  ))
// Xd_0__inst_mult_31_126  = SHARE((din_a[219] & (din_b[221] & (din_a[218] & din_b[222]))))

	.dataa(!din_a[219]),
	.datab(!din_b[221]),
	.datac(!din_a[218]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_117 ),
	.sharein(Xd_0__inst_mult_31_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_124 ),
	.cout(Xd_0__inst_mult_31_125 ),
	.shareout(Xd_0__inst_mult_31_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_39 (
// Equation(s):
// Xd_0__inst_mult_30_128  = SUM(( (!din_a[215] & (((din_a[214] & din_b[213])))) # (din_a[215] & (!din_b[212] $ (((!din_a[214]) # (!din_b[213]))))) ) + ( Xd_0__inst_mult_30_122  ) + ( Xd_0__inst_mult_30_121  ))
// Xd_0__inst_mult_30_129  = CARRY(( (!din_a[215] & (((din_a[214] & din_b[213])))) # (din_a[215] & (!din_b[212] $ (((!din_a[214]) # (!din_b[213]))))) ) + ( Xd_0__inst_mult_30_122  ) + ( Xd_0__inst_mult_30_121  ))
// Xd_0__inst_mult_30_130  = SHARE((din_a[215] & (din_b[212] & (din_a[214] & din_b[213]))))

	.dataa(!din_a[215]),
	.datab(!din_b[212]),
	.datac(!din_a[214]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_121 ),
	.sharein(Xd_0__inst_mult_30_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_128 ),
	.cout(Xd_0__inst_mult_30_129 ),
	.shareout(Xd_0__inst_mult_30_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_40 (
// Equation(s):
// Xd_0__inst_mult_30_132  = SUM(( (!din_a[213] & (((din_a[212] & din_b[215])))) # (din_a[213] & (!din_b[214] $ (((!din_a[212]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_126  ) + ( Xd_0__inst_mult_30_125  ))
// Xd_0__inst_mult_30_133  = CARRY(( (!din_a[213] & (((din_a[212] & din_b[215])))) # (din_a[213] & (!din_b[214] $ (((!din_a[212]) # (!din_b[215]))))) ) + ( Xd_0__inst_mult_30_126  ) + ( Xd_0__inst_mult_30_125  ))
// Xd_0__inst_mult_30_134  = SHARE((din_a[213] & (din_b[214] & (din_a[212] & din_b[215]))))

	.dataa(!din_a[213]),
	.datab(!din_b[214]),
	.datac(!din_a[212]),
	.datad(!din_b[215]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_125 ),
	.sharein(Xd_0__inst_mult_30_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_132 ),
	.cout(Xd_0__inst_mult_30_133 ),
	.shareout(Xd_0__inst_mult_30_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_39 (
// Equation(s):
// Xd_0__inst_mult_31_128  = SUM(( (!din_a[222] & (((din_a[221] & din_b[220])))) # (din_a[222] & (!din_b[219] $ (((!din_a[221]) # (!din_b[220]))))) ) + ( Xd_0__inst_mult_31_122  ) + ( Xd_0__inst_mult_31_121  ))
// Xd_0__inst_mult_31_129  = CARRY(( (!din_a[222] & (((din_a[221] & din_b[220])))) # (din_a[222] & (!din_b[219] $ (((!din_a[221]) # (!din_b[220]))))) ) + ( Xd_0__inst_mult_31_122  ) + ( Xd_0__inst_mult_31_121  ))
// Xd_0__inst_mult_31_130  = SHARE((din_a[222] & (din_b[219] & (din_a[221] & din_b[220]))))

	.dataa(!din_a[222]),
	.datab(!din_b[219]),
	.datac(!din_a[221]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_121 ),
	.sharein(Xd_0__inst_mult_31_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_128 ),
	.cout(Xd_0__inst_mult_31_129 ),
	.shareout(Xd_0__inst_mult_31_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_40 (
// Equation(s):
// Xd_0__inst_mult_31_132  = SUM(( (!din_a[220] & (((din_a[219] & din_b[222])))) # (din_a[220] & (!din_b[221] $ (((!din_a[219]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_126  ) + ( Xd_0__inst_mult_31_125  ))
// Xd_0__inst_mult_31_133  = CARRY(( (!din_a[220] & (((din_a[219] & din_b[222])))) # (din_a[220] & (!din_b[221] $ (((!din_a[219]) # (!din_b[222]))))) ) + ( Xd_0__inst_mult_31_126  ) + ( Xd_0__inst_mult_31_125  ))
// Xd_0__inst_mult_31_134  = SHARE((din_a[220] & (din_b[221] & (din_a[219] & din_b[222]))))

	.dataa(!din_a[220]),
	.datab(!din_b[221]),
	.datac(!din_a[219]),
	.datad(!din_b[222]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_125 ),
	.sharein(Xd_0__inst_mult_31_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_132 ),
	.cout(Xd_0__inst_mult_31_133 ),
	.shareout(Xd_0__inst_mult_31_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_41 (
// Equation(s):
// Xd_0__inst_mult_30_136  = SUM(( (!din_a[215] & (((din_a[214] & din_b[214])))) # (din_a[215] & (!din_b[213] $ (((!din_a[214]) # (!din_b[214]))))) ) + ( Xd_0__inst_mult_30_130  ) + ( Xd_0__inst_mult_30_129  ))
// Xd_0__inst_mult_30_137  = CARRY(( (!din_a[215] & (((din_a[214] & din_b[214])))) # (din_a[215] & (!din_b[213] $ (((!din_a[214]) # (!din_b[214]))))) ) + ( Xd_0__inst_mult_30_130  ) + ( Xd_0__inst_mult_30_129  ))
// Xd_0__inst_mult_30_138  = SHARE((din_a[215] & (din_b[213] & (din_a[214] & din_b[214]))))

	.dataa(!din_a[215]),
	.datab(!din_b[213]),
	.datac(!din_a[214]),
	.datad(!din_b[214]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_129 ),
	.sharein(Xd_0__inst_mult_30_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_136 ),
	.cout(Xd_0__inst_mult_30_137 ),
	.shareout(Xd_0__inst_mult_30_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_42 (
// Equation(s):
// Xd_0__inst_mult_30_140  = SUM(( (din_a[213] & din_b[215]) ) + ( Xd_0__inst_mult_30_134  ) + ( Xd_0__inst_mult_30_133  ))
// Xd_0__inst_mult_30_141  = CARRY(( (din_a[213] & din_b[215]) ) + ( Xd_0__inst_mult_30_134  ) + ( Xd_0__inst_mult_30_133  ))
// Xd_0__inst_mult_30_142  = SHARE(GND)

	.dataa(!din_a[213]),
	.datab(!din_b[215]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_133 ),
	.sharein(Xd_0__inst_mult_30_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_140 ),
	.cout(Xd_0__inst_mult_30_141 ),
	.shareout(Xd_0__inst_mult_30_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_41 (
// Equation(s):
// Xd_0__inst_mult_31_136  = SUM(( (!din_a[222] & (((din_a[221] & din_b[221])))) # (din_a[222] & (!din_b[220] $ (((!din_a[221]) # (!din_b[221]))))) ) + ( Xd_0__inst_mult_31_130  ) + ( Xd_0__inst_mult_31_129  ))
// Xd_0__inst_mult_31_137  = CARRY(( (!din_a[222] & (((din_a[221] & din_b[221])))) # (din_a[222] & (!din_b[220] $ (((!din_a[221]) # (!din_b[221]))))) ) + ( Xd_0__inst_mult_31_130  ) + ( Xd_0__inst_mult_31_129  ))
// Xd_0__inst_mult_31_138  = SHARE((din_a[222] & (din_b[220] & (din_a[221] & din_b[221]))))

	.dataa(!din_a[222]),
	.datab(!din_b[220]),
	.datac(!din_a[221]),
	.datad(!din_b[221]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_129 ),
	.sharein(Xd_0__inst_mult_31_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_136 ),
	.cout(Xd_0__inst_mult_31_137 ),
	.shareout(Xd_0__inst_mult_31_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_42 (
// Equation(s):
// Xd_0__inst_mult_31_140  = SUM(( (din_a[220] & din_b[222]) ) + ( Xd_0__inst_mult_31_134  ) + ( Xd_0__inst_mult_31_133  ))
// Xd_0__inst_mult_31_141  = CARRY(( (din_a[220] & din_b[222]) ) + ( Xd_0__inst_mult_31_134  ) + ( Xd_0__inst_mult_31_133  ))
// Xd_0__inst_mult_31_142  = SHARE(GND)

	.dataa(!din_a[220]),
	.datab(!din_b[222]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_133 ),
	.sharein(Xd_0__inst_mult_31_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_140 ),
	.cout(Xd_0__inst_mult_31_141 ),
	.shareout(Xd_0__inst_mult_31_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_43 (
// Equation(s):
// Xd_0__inst_mult_30_144  = SUM(( (din_a[215] & din_b[214]) ) + ( Xd_0__inst_mult_30_138  ) + ( Xd_0__inst_mult_30_137  ))
// Xd_0__inst_mult_30_145  = CARRY(( (din_a[215] & din_b[214]) ) + ( Xd_0__inst_mult_30_138  ) + ( Xd_0__inst_mult_30_137  ))
// Xd_0__inst_mult_30_146  = SHARE(GND)

	.dataa(!din_a[215]),
	.datab(!din_b[214]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_137 ),
	.sharein(Xd_0__inst_mult_30_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_144 ),
	.cout(Xd_0__inst_mult_30_145 ),
	.shareout(Xd_0__inst_mult_30_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_44 (
// Equation(s):
// Xd_0__inst_mult_30_148  = SUM(( GND ) + ( Xd_0__inst_mult_30_142  ) + ( Xd_0__inst_mult_30_141  ))
// Xd_0__inst_mult_30_149  = CARRY(( GND ) + ( Xd_0__inst_mult_30_142  ) + ( Xd_0__inst_mult_30_141  ))
// Xd_0__inst_mult_30_150  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_141 ),
	.sharein(Xd_0__inst_mult_30_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_148 ),
	.cout(Xd_0__inst_mult_30_149 ),
	.shareout(Xd_0__inst_mult_30_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_43 (
// Equation(s):
// Xd_0__inst_mult_31_144  = SUM(( (din_a[222] & din_b[221]) ) + ( Xd_0__inst_mult_31_138  ) + ( Xd_0__inst_mult_31_137  ))
// Xd_0__inst_mult_31_145  = CARRY(( (din_a[222] & din_b[221]) ) + ( Xd_0__inst_mult_31_138  ) + ( Xd_0__inst_mult_31_137  ))
// Xd_0__inst_mult_31_146  = SHARE(GND)

	.dataa(!din_a[222]),
	.datab(!din_b[221]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_137 ),
	.sharein(Xd_0__inst_mult_31_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_144 ),
	.cout(Xd_0__inst_mult_31_145 ),
	.shareout(Xd_0__inst_mult_31_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_44 (
// Equation(s):
// Xd_0__inst_mult_31_148  = SUM(( GND ) + ( Xd_0__inst_mult_31_142  ) + ( Xd_0__inst_mult_31_141  ))
// Xd_0__inst_mult_31_149  = CARRY(( GND ) + ( Xd_0__inst_mult_31_142  ) + ( Xd_0__inst_mult_31_141  ))
// Xd_0__inst_mult_31_150  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_141 ),
	.sharein(Xd_0__inst_mult_31_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_148 ),
	.cout(Xd_0__inst_mult_31_149 ),
	.shareout(Xd_0__inst_mult_31_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_45 (
// Equation(s):
// Xd_0__inst_mult_30_152  = SUM(( GND ) + ( Xd_0__inst_mult_30_146  ) + ( Xd_0__inst_mult_30_145  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_145 ),
	.sharein(Xd_0__inst_mult_30_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_45 (
// Equation(s):
// Xd_0__inst_mult_31_152  = SUM(( GND ) + ( Xd_0__inst_mult_31_146  ) + ( Xd_0__inst_mult_31_145  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_145 ),
	.sharein(Xd_0__inst_mult_31_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_32 (
// Equation(s):
// Xd_0__inst_mult_14_100  = SUM(( GND ) + ( Xd_0__inst_mult_14_146  ) + ( Xd_0__inst_mult_14_145  ))
// Xd_0__inst_mult_14_101  = CARRY(( GND ) + ( Xd_0__inst_mult_14_146  ) + ( Xd_0__inst_mult_14_145  ))
// Xd_0__inst_mult_14_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_145 ),
	.sharein(Xd_0__inst_mult_14_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_100 ),
	.cout(Xd_0__inst_mult_14_101 ),
	.shareout(Xd_0__inst_mult_14_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_32 (
// Equation(s):
// Xd_0__inst_mult_19_100  = SUM(( GND ) + ( Xd_0__inst_mult_19_146  ) + ( Xd_0__inst_mult_19_145  ))
// Xd_0__inst_mult_19_101  = CARRY(( GND ) + ( Xd_0__inst_mult_19_146  ) + ( Xd_0__inst_mult_19_145  ))
// Xd_0__inst_mult_19_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_145 ),
	.sharein(Xd_0__inst_mult_19_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_100 ),
	.cout(Xd_0__inst_mult_19_101 ),
	.shareout(Xd_0__inst_mult_19_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_32 (
// Equation(s):
// Xd_0__inst_mult_21_100  = SUM(( GND ) + ( Xd_0__inst_mult_21_146  ) + ( Xd_0__inst_mult_21_145  ))
// Xd_0__inst_mult_21_101  = CARRY(( GND ) + ( Xd_0__inst_mult_21_146  ) + ( Xd_0__inst_mult_21_145  ))
// Xd_0__inst_mult_21_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_145 ),
	.sharein(Xd_0__inst_mult_21_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_100 ),
	.cout(Xd_0__inst_mult_21_101 ),
	.shareout(Xd_0__inst_mult_21_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_32 (
// Equation(s):
// Xd_0__inst_mult_18_100  = SUM(( GND ) + ( Xd_0__inst_mult_18_146  ) + ( Xd_0__inst_mult_18_145  ))
// Xd_0__inst_mult_18_101  = CARRY(( GND ) + ( Xd_0__inst_mult_18_146  ) + ( Xd_0__inst_mult_18_145  ))
// Xd_0__inst_mult_18_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_145 ),
	.sharein(Xd_0__inst_mult_18_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_100 ),
	.cout(Xd_0__inst_mult_18_101 ),
	.shareout(Xd_0__inst_mult_18_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_32 (
// Equation(s):
// Xd_0__inst_mult_17_100  = SUM(( GND ) + ( Xd_0__inst_mult_17_146  ) + ( Xd_0__inst_mult_17_145  ))
// Xd_0__inst_mult_17_101  = CARRY(( GND ) + ( Xd_0__inst_mult_17_146  ) + ( Xd_0__inst_mult_17_145  ))
// Xd_0__inst_mult_17_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_145 ),
	.sharein(Xd_0__inst_mult_17_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_100 ),
	.cout(Xd_0__inst_mult_17_101 ),
	.shareout(Xd_0__inst_mult_17_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_32 (
// Equation(s):
// Xd_0__inst_mult_16_100  = SUM(( GND ) + ( Xd_0__inst_mult_16_146  ) + ( Xd_0__inst_mult_16_145  ))
// Xd_0__inst_mult_16_101  = CARRY(( GND ) + ( Xd_0__inst_mult_16_146  ) + ( Xd_0__inst_mult_16_145  ))
// Xd_0__inst_mult_16_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_145 ),
	.sharein(Xd_0__inst_mult_16_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_100 ),
	.cout(Xd_0__inst_mult_16_101 ),
	.shareout(Xd_0__inst_mult_16_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_32 (
// Equation(s):
// Xd_0__inst_mult_20_100  = SUM(( GND ) + ( Xd_0__inst_mult_20_146  ) + ( Xd_0__inst_mult_20_145  ))
// Xd_0__inst_mult_20_101  = CARRY(( GND ) + ( Xd_0__inst_mult_20_146  ) + ( Xd_0__inst_mult_20_145  ))
// Xd_0__inst_mult_20_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_145 ),
	.sharein(Xd_0__inst_mult_20_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_100 ),
	.cout(Xd_0__inst_mult_20_101 ),
	.shareout(Xd_0__inst_mult_20_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_32 (
// Equation(s):
// Xd_0__inst_mult_28_100  = SUM(( GND ) + ( Xd_0__inst_mult_28_146  ) + ( Xd_0__inst_mult_28_145  ))
// Xd_0__inst_mult_28_101  = CARRY(( GND ) + ( Xd_0__inst_mult_28_146  ) + ( Xd_0__inst_mult_28_145  ))
// Xd_0__inst_mult_28_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_145 ),
	.sharein(Xd_0__inst_mult_28_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_100 ),
	.cout(Xd_0__inst_mult_28_101 ),
	.shareout(Xd_0__inst_mult_28_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_32 (
// Equation(s):
// Xd_0__inst_mult_12_100  = SUM(( GND ) + ( Xd_0__inst_mult_12_146  ) + ( Xd_0__inst_mult_12_145  ))
// Xd_0__inst_mult_12_101  = CARRY(( GND ) + ( Xd_0__inst_mult_12_146  ) + ( Xd_0__inst_mult_12_145  ))
// Xd_0__inst_mult_12_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_145 ),
	.sharein(Xd_0__inst_mult_12_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_100 ),
	.cout(Xd_0__inst_mult_12_101 ),
	.shareout(Xd_0__inst_mult_12_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_32 (
// Equation(s):
// Xd_0__inst_mult_5_100  = SUM(( GND ) + ( Xd_0__inst_mult_5_146  ) + ( Xd_0__inst_mult_5_145  ))
// Xd_0__inst_mult_5_101  = CARRY(( GND ) + ( Xd_0__inst_mult_5_146  ) + ( Xd_0__inst_mult_5_145  ))
// Xd_0__inst_mult_5_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_145 ),
	.sharein(Xd_0__inst_mult_5_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_100 ),
	.cout(Xd_0__inst_mult_5_101 ),
	.shareout(Xd_0__inst_mult_5_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_32 (
// Equation(s):
// Xd_0__inst_mult_15_100  = SUM(( GND ) + ( Xd_0__inst_mult_15_146  ) + ( Xd_0__inst_mult_15_145  ))
// Xd_0__inst_mult_15_101  = CARRY(( GND ) + ( Xd_0__inst_mult_15_146  ) + ( Xd_0__inst_mult_15_145  ))
// Xd_0__inst_mult_15_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_145 ),
	.sharein(Xd_0__inst_mult_15_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_100 ),
	.cout(Xd_0__inst_mult_15_101 ),
	.shareout(Xd_0__inst_mult_15_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_32 (
// Equation(s):
// Xd_0__inst_mult_7_100  = SUM(( GND ) + ( Xd_0__inst_mult_7_146  ) + ( Xd_0__inst_mult_7_145  ))
// Xd_0__inst_mult_7_101  = CARRY(( GND ) + ( Xd_0__inst_mult_7_146  ) + ( Xd_0__inst_mult_7_145  ))
// Xd_0__inst_mult_7_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_145 ),
	.sharein(Xd_0__inst_mult_7_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_100 ),
	.cout(Xd_0__inst_mult_7_101 ),
	.shareout(Xd_0__inst_mult_7_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_33 (
// Equation(s):
// Xd_0__inst_mult_25_104  = SUM(( (din_a[178] & din_b[180]) ) + ( Xd_0__inst_mult_25_142  ) + ( Xd_0__inst_mult_25_141  ))
// Xd_0__inst_mult_25_105  = CARRY(( (din_a[178] & din_b[180]) ) + ( Xd_0__inst_mult_25_142  ) + ( Xd_0__inst_mult_25_141  ))
// Xd_0__inst_mult_25_106  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[180]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_141 ),
	.sharein(Xd_0__inst_mult_25_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_104 ),
	.cout(Xd_0__inst_mult_25_105 ),
	.shareout(Xd_0__inst_mult_25_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_33 (
// Equation(s):
// Xd_0__inst_mult_22_104  = SUM(( (din_a[157] & din_b[159]) ) + ( Xd_0__inst_mult_22_142  ) + ( Xd_0__inst_mult_22_141  ))
// Xd_0__inst_mult_22_105  = CARRY(( (din_a[157] & din_b[159]) ) + ( Xd_0__inst_mult_22_142  ) + ( Xd_0__inst_mult_22_141  ))
// Xd_0__inst_mult_22_106  = SHARE(GND)

	.dataa(!din_a[157]),
	.datab(!din_b[159]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_141 ),
	.sharein(Xd_0__inst_mult_22_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_104 ),
	.cout(Xd_0__inst_mult_22_105 ),
	.shareout(Xd_0__inst_mult_22_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_32 (
// Equation(s):
// Xd_0__inst_mult_6_100  = SUM(( GND ) + ( Xd_0__inst_mult_6_146  ) + ( Xd_0__inst_mult_6_145  ))
// Xd_0__inst_mult_6_101  = CARRY(( GND ) + ( Xd_0__inst_mult_6_146  ) + ( Xd_0__inst_mult_6_145  ))
// Xd_0__inst_mult_6_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_145 ),
	.sharein(Xd_0__inst_mult_6_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_100 ),
	.cout(Xd_0__inst_mult_6_101 ),
	.shareout(Xd_0__inst_mult_6_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_32 (
// Equation(s):
// Xd_0__inst_mult_9_100  = SUM(( GND ) + ( Xd_0__inst_mult_9_146  ) + ( Xd_0__inst_mult_9_145  ))
// Xd_0__inst_mult_9_101  = CARRY(( GND ) + ( Xd_0__inst_mult_9_146  ) + ( Xd_0__inst_mult_9_145  ))
// Xd_0__inst_mult_9_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_145 ),
	.sharein(Xd_0__inst_mult_9_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_100 ),
	.cout(Xd_0__inst_mult_9_101 ),
	.shareout(Xd_0__inst_mult_9_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_32 (
// Equation(s):
// Xd_0__inst_mult_8_100  = SUM(( GND ) + ( Xd_0__inst_mult_8_146  ) + ( Xd_0__inst_mult_8_145  ))
// Xd_0__inst_mult_8_101  = CARRY(( GND ) + ( Xd_0__inst_mult_8_146  ) + ( Xd_0__inst_mult_8_145  ))
// Xd_0__inst_mult_8_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_145 ),
	.sharein(Xd_0__inst_mult_8_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_100 ),
	.cout(Xd_0__inst_mult_8_101 ),
	.shareout(Xd_0__inst_mult_8_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_32 (
// Equation(s):
// Xd_0__inst_mult_11_100  = SUM(( GND ) + ( Xd_0__inst_mult_11_146  ) + ( Xd_0__inst_mult_11_145  ))
// Xd_0__inst_mult_11_101  = CARRY(( GND ) + ( Xd_0__inst_mult_11_146  ) + ( Xd_0__inst_mult_11_145  ))
// Xd_0__inst_mult_11_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_145 ),
	.sharein(Xd_0__inst_mult_11_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_100 ),
	.cout(Xd_0__inst_mult_11_101 ),
	.shareout(Xd_0__inst_mult_11_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_32 (
// Equation(s):
// Xd_0__inst_mult_10_100  = SUM(( GND ) + ( Xd_0__inst_mult_10_146  ) + ( Xd_0__inst_mult_10_145  ))
// Xd_0__inst_mult_10_101  = CARRY(( GND ) + ( Xd_0__inst_mult_10_146  ) + ( Xd_0__inst_mult_10_145  ))
// Xd_0__inst_mult_10_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_145 ),
	.sharein(Xd_0__inst_mult_10_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_100 ),
	.cout(Xd_0__inst_mult_10_101 ),
	.shareout(Xd_0__inst_mult_10_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_32 (
// Equation(s):
// Xd_0__inst_mult_13_100  = SUM(( GND ) + ( Xd_0__inst_mult_13_146  ) + ( Xd_0__inst_mult_13_145  ))
// Xd_0__inst_mult_13_101  = CARRY(( GND ) + ( Xd_0__inst_mult_13_146  ) + ( Xd_0__inst_mult_13_145  ))
// Xd_0__inst_mult_13_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_145 ),
	.sharein(Xd_0__inst_mult_13_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_100 ),
	.cout(Xd_0__inst_mult_13_101 ),
	.shareout(Xd_0__inst_mult_13_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_32 (
// Equation(s):
// Xd_0__inst_mult_4_100  = SUM(( GND ) + ( Xd_0__inst_mult_4_146  ) + ( Xd_0__inst_mult_4_145  ))
// Xd_0__inst_mult_4_101  = CARRY(( GND ) + ( Xd_0__inst_mult_4_146  ) + ( Xd_0__inst_mult_4_145  ))
// Xd_0__inst_mult_4_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_145 ),
	.sharein(Xd_0__inst_mult_4_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_100 ),
	.cout(Xd_0__inst_mult_4_101 ),
	.shareout(Xd_0__inst_mult_4_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_32 (
// Equation(s):
// Xd_0__inst_mult_2_100  = SUM(( GND ) + ( Xd_0__inst_mult_2_146  ) + ( Xd_0__inst_mult_2_145  ))
// Xd_0__inst_mult_2_101  = CARRY(( GND ) + ( Xd_0__inst_mult_2_146  ) + ( Xd_0__inst_mult_2_145  ))
// Xd_0__inst_mult_2_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_145 ),
	.sharein(Xd_0__inst_mult_2_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_100 ),
	.cout(Xd_0__inst_mult_2_101 ),
	.shareout(Xd_0__inst_mult_2_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_32 (
// Equation(s):
// Xd_0__inst_mult_3_100  = SUM(( GND ) + ( Xd_0__inst_mult_3_146  ) + ( Xd_0__inst_mult_3_145  ))
// Xd_0__inst_mult_3_101  = CARRY(( GND ) + ( Xd_0__inst_mult_3_146  ) + ( Xd_0__inst_mult_3_145  ))
// Xd_0__inst_mult_3_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_145 ),
	.sharein(Xd_0__inst_mult_3_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_100 ),
	.cout(Xd_0__inst_mult_3_101 ),
	.shareout(Xd_0__inst_mult_3_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_32 (
// Equation(s):
// Xd_0__inst_mult_0_100  = SUM(( GND ) + ( Xd_0__inst_mult_0_146  ) + ( Xd_0__inst_mult_0_145  ))
// Xd_0__inst_mult_0_101  = CARRY(( GND ) + ( Xd_0__inst_mult_0_146  ) + ( Xd_0__inst_mult_0_145  ))
// Xd_0__inst_mult_0_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_145 ),
	.sharein(Xd_0__inst_mult_0_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_100 ),
	.cout(Xd_0__inst_mult_0_101 ),
	.shareout(Xd_0__inst_mult_0_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_32 (
// Equation(s):
// Xd_0__inst_mult_1_100  = SUM(( GND ) + ( Xd_0__inst_mult_1_146  ) + ( Xd_0__inst_mult_1_145  ))
// Xd_0__inst_mult_1_101  = CARRY(( GND ) + ( Xd_0__inst_mult_1_146  ) + ( Xd_0__inst_mult_1_145  ))
// Xd_0__inst_mult_1_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_145 ),
	.sharein(Xd_0__inst_mult_1_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_100 ),
	.cout(Xd_0__inst_mult_1_101 ),
	.shareout(Xd_0__inst_mult_1_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_32 (
// Equation(s):
// Xd_0__inst_mult_23_100  = SUM(( GND ) + ( Xd_0__inst_mult_23_146  ) + ( Xd_0__inst_mult_23_145  ))
// Xd_0__inst_mult_23_101  = CARRY(( GND ) + ( Xd_0__inst_mult_23_146  ) + ( Xd_0__inst_mult_23_145  ))
// Xd_0__inst_mult_23_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_145 ),
	.sharein(Xd_0__inst_mult_23_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_100 ),
	.cout(Xd_0__inst_mult_23_101 ),
	.shareout(Xd_0__inst_mult_23_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_32 (
// Equation(s):
// Xd_0__inst_mult_29_100  = SUM(( GND ) + ( Xd_0__inst_mult_29_146  ) + ( Xd_0__inst_mult_29_145  ))
// Xd_0__inst_mult_29_101  = CARRY(( GND ) + ( Xd_0__inst_mult_29_146  ) + ( Xd_0__inst_mult_29_145  ))
// Xd_0__inst_mult_29_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_145 ),
	.sharein(Xd_0__inst_mult_29_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_100 ),
	.cout(Xd_0__inst_mult_29_101 ),
	.shareout(Xd_0__inst_mult_29_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_32 (
// Equation(s):
// Xd_0__inst_mult_26_100  = SUM(( GND ) + ( Xd_0__inst_mult_26_146  ) + ( Xd_0__inst_mult_26_145  ))
// Xd_0__inst_mult_26_101  = CARRY(( GND ) + ( Xd_0__inst_mult_26_146  ) + ( Xd_0__inst_mult_26_145  ))
// Xd_0__inst_mult_26_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_145 ),
	.sharein(Xd_0__inst_mult_26_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_100 ),
	.cout(Xd_0__inst_mult_26_101 ),
	.shareout(Xd_0__inst_mult_26_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_32 (
// Equation(s):
// Xd_0__inst_mult_24_100  = SUM(( GND ) + ( Xd_0__inst_mult_24_146  ) + ( Xd_0__inst_mult_24_145  ))
// Xd_0__inst_mult_24_101  = CARRY(( GND ) + ( Xd_0__inst_mult_24_146  ) + ( Xd_0__inst_mult_24_145  ))
// Xd_0__inst_mult_24_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_145 ),
	.sharein(Xd_0__inst_mult_24_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_100 ),
	.cout(Xd_0__inst_mult_24_101 ),
	.shareout(Xd_0__inst_mult_24_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_32 (
// Equation(s):
// Xd_0__inst_mult_27_100  = SUM(( GND ) + ( Xd_0__inst_mult_27_146  ) + ( Xd_0__inst_mult_27_145  ))
// Xd_0__inst_mult_27_101  = CARRY(( GND ) + ( Xd_0__inst_mult_27_146  ) + ( Xd_0__inst_mult_27_145  ))
// Xd_0__inst_mult_27_102  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_145 ),
	.sharein(Xd_0__inst_mult_27_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_100 ),
	.cout(Xd_0__inst_mult_27_101 ),
	.shareout(Xd_0__inst_mult_27_102 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_33 (
// Equation(s):
// Xd_0__inst_mult_28_104  = SUM(( (!din_a[198] & (((din_a[197] & din_b[198])))) # (din_a[198] & (!din_b[197] $ (((!din_a[197]) # (!din_b[198]))))) ) + ( Xd_0__inst_mult_28_94  ) + ( Xd_0__inst_mult_28_93  ))
// Xd_0__inst_mult_28_105  = CARRY(( (!din_a[198] & (((din_a[197] & din_b[198])))) # (din_a[198] & (!din_b[197] $ (((!din_a[197]) # (!din_b[198]))))) ) + ( Xd_0__inst_mult_28_94  ) + ( Xd_0__inst_mult_28_93  ))
// Xd_0__inst_mult_28_106  = SHARE((din_a[198] & (din_b[197] & (din_a[197] & din_b[198]))))

	.dataa(!din_a[198]),
	.datab(!din_b[197]),
	.datac(!din_a[197]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_93 ),
	.sharein(Xd_0__inst_mult_28_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_104 ),
	.cout(Xd_0__inst_mult_28_105 ),
	.shareout(Xd_0__inst_mult_28_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_33 (
// Equation(s):
// Xd_0__inst_mult_29_104  = SUM(( (!din_a[205] & (((din_a[204] & din_b[205])))) # (din_a[205] & (!din_b[204] $ (((!din_a[204]) # (!din_b[205]))))) ) + ( Xd_0__inst_mult_29_94  ) + ( Xd_0__inst_mult_29_93  ))
// Xd_0__inst_mult_29_105  = CARRY(( (!din_a[205] & (((din_a[204] & din_b[205])))) # (din_a[205] & (!din_b[204] $ (((!din_a[204]) # (!din_b[205]))))) ) + ( Xd_0__inst_mult_29_94  ) + ( Xd_0__inst_mult_29_93  ))
// Xd_0__inst_mult_29_106  = SHARE((din_a[205] & (din_b[204] & (din_a[204] & din_b[205]))))

	.dataa(!din_a[205]),
	.datab(!din_b[204]),
	.datac(!din_a[204]),
	.datad(!din_b[205]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_93 ),
	.sharein(Xd_0__inst_mult_29_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_104 ),
	.cout(Xd_0__inst_mult_29_105 ),
	.shareout(Xd_0__inst_mult_29_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_33 (
// Equation(s):
// Xd_0__inst_mult_26_104  = SUM(( (!din_a[184] & (((din_a[183] & din_b[184])))) # (din_a[184] & (!din_b[183] $ (((!din_a[183]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_26_94  ) + ( Xd_0__inst_mult_26_93  ))
// Xd_0__inst_mult_26_105  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[184])))) # (din_a[184] & (!din_b[183] $ (((!din_a[183]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_26_94  ) + ( Xd_0__inst_mult_26_93  ))
// Xd_0__inst_mult_26_106  = SHARE((din_a[184] & (din_b[183] & (din_a[183] & din_b[184]))))

	.dataa(!din_a[184]),
	.datab(!din_b[183]),
	.datac(!din_a[183]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_93 ),
	.sharein(Xd_0__inst_mult_26_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_104 ),
	.cout(Xd_0__inst_mult_26_105 ),
	.shareout(Xd_0__inst_mult_26_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_33 (
// Equation(s):
// Xd_0__inst_mult_27_104  = SUM(( (!din_a[191] & (((din_a[190] & din_b[191])))) # (din_a[191] & (!din_b[190] $ (((!din_a[190]) # (!din_b[191]))))) ) + ( Xd_0__inst_mult_27_94  ) + ( Xd_0__inst_mult_27_93  ))
// Xd_0__inst_mult_27_105  = CARRY(( (!din_a[191] & (((din_a[190] & din_b[191])))) # (din_a[191] & (!din_b[190] $ (((!din_a[190]) # (!din_b[191]))))) ) + ( Xd_0__inst_mult_27_94  ) + ( Xd_0__inst_mult_27_93  ))
// Xd_0__inst_mult_27_106  = SHARE((din_a[191] & (din_b[190] & (din_a[190] & din_b[191]))))

	.dataa(!din_a[191]),
	.datab(!din_b[190]),
	.datac(!din_a[190]),
	.datad(!din_b[191]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_93 ),
	.sharein(Xd_0__inst_mult_27_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_104 ),
	.cout(Xd_0__inst_mult_27_105 ),
	.shareout(Xd_0__inst_mult_27_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_33 (
// Equation(s):
// Xd_0__inst_mult_24_104  = SUM(( (!din_a[170] & (((din_a[169] & din_b[170])))) # (din_a[170] & (!din_b[169] $ (((!din_a[169]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_24_94  ) + ( Xd_0__inst_mult_24_93  ))
// Xd_0__inst_mult_24_105  = CARRY(( (!din_a[170] & (((din_a[169] & din_b[170])))) # (din_a[170] & (!din_b[169] $ (((!din_a[169]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_24_94  ) + ( Xd_0__inst_mult_24_93  ))
// Xd_0__inst_mult_24_106  = SHARE((din_a[170] & (din_b[169] & (din_a[169] & din_b[170]))))

	.dataa(!din_a[170]),
	.datab(!din_b[169]),
	.datac(!din_a[169]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_93 ),
	.sharein(Xd_0__inst_mult_24_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_104 ),
	.cout(Xd_0__inst_mult_24_105 ),
	.shareout(Xd_0__inst_mult_24_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_34 (
// Equation(s):
// Xd_0__inst_mult_25_108  = SUM(( (!din_a[177] & (((din_a[176] & din_b[177])))) # (din_a[177] & (!din_b[176] $ (((!din_a[176]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_25_98  ) + ( Xd_0__inst_mult_25_97  ))
// Xd_0__inst_mult_25_109  = CARRY(( (!din_a[177] & (((din_a[176] & din_b[177])))) # (din_a[177] & (!din_b[176] $ (((!din_a[176]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_25_98  ) + ( Xd_0__inst_mult_25_97  ))
// Xd_0__inst_mult_25_110  = SHARE((din_a[177] & (din_b[176] & (din_a[176] & din_b[177]))))

	.dataa(!din_a[177]),
	.datab(!din_b[176]),
	.datac(!din_a[176]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_97 ),
	.sharein(Xd_0__inst_mult_25_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_108 ),
	.cout(Xd_0__inst_mult_25_109 ),
	.shareout(Xd_0__inst_mult_25_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_34 (
// Equation(s):
// Xd_0__inst_mult_22_108  = SUM(( (!din_a[156] & (((din_a[155] & din_b[156])))) # (din_a[156] & (!din_b[155] $ (((!din_a[155]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_22_98  ) + ( Xd_0__inst_mult_22_97  ))
// Xd_0__inst_mult_22_109  = CARRY(( (!din_a[156] & (((din_a[155] & din_b[156])))) # (din_a[156] & (!din_b[155] $ (((!din_a[155]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_22_98  ) + ( Xd_0__inst_mult_22_97  ))
// Xd_0__inst_mult_22_110  = SHARE((din_a[156] & (din_b[155] & (din_a[155] & din_b[156]))))

	.dataa(!din_a[156]),
	.datab(!din_b[155]),
	.datac(!din_a[155]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_97 ),
	.sharein(Xd_0__inst_mult_22_98 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_108 ),
	.cout(Xd_0__inst_mult_22_109 ),
	.shareout(Xd_0__inst_mult_22_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_33 (
// Equation(s):
// Xd_0__inst_mult_23_104  = SUM(( (!din_a[163] & (((din_a[162] & din_b[163])))) # (din_a[163] & (!din_b[162] $ (((!din_a[162]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_23_94  ) + ( Xd_0__inst_mult_23_93  ))
// Xd_0__inst_mult_23_105  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[163])))) # (din_a[163] & (!din_b[162] $ (((!din_a[162]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_23_94  ) + ( Xd_0__inst_mult_23_93  ))
// Xd_0__inst_mult_23_106  = SHARE((din_a[163] & (din_b[162] & (din_a[162] & din_b[163]))))

	.dataa(!din_a[163]),
	.datab(!din_b[162]),
	.datac(!din_a[162]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_93 ),
	.sharein(Xd_0__inst_mult_23_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_104 ),
	.cout(Xd_0__inst_mult_23_105 ),
	.shareout(Xd_0__inst_mult_23_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_33 (
// Equation(s):
// Xd_0__inst_mult_20_104  = SUM(( (!din_a[142] & (((din_a[141] & din_b[142])))) # (din_a[142] & (!din_b[141] $ (((!din_a[141]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_20_94  ) + ( Xd_0__inst_mult_20_93  ))
// Xd_0__inst_mult_20_105  = CARRY(( (!din_a[142] & (((din_a[141] & din_b[142])))) # (din_a[142] & (!din_b[141] $ (((!din_a[141]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_20_94  ) + ( Xd_0__inst_mult_20_93  ))
// Xd_0__inst_mult_20_106  = SHARE((din_a[142] & (din_b[141] & (din_a[141] & din_b[142]))))

	.dataa(!din_a[142]),
	.datab(!din_b[141]),
	.datac(!din_a[141]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_93 ),
	.sharein(Xd_0__inst_mult_20_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_104 ),
	.cout(Xd_0__inst_mult_20_105 ),
	.shareout(Xd_0__inst_mult_20_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_33 (
// Equation(s):
// Xd_0__inst_mult_21_104  = SUM(( (!din_a[149] & (((din_a[148] & din_b[149])))) # (din_a[149] & (!din_b[148] $ (((!din_a[148]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_21_94  ) + ( Xd_0__inst_mult_21_93  ))
// Xd_0__inst_mult_21_105  = CARRY(( (!din_a[149] & (((din_a[148] & din_b[149])))) # (din_a[149] & (!din_b[148] $ (((!din_a[148]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_21_94  ) + ( Xd_0__inst_mult_21_93  ))
// Xd_0__inst_mult_21_106  = SHARE((din_a[149] & (din_b[148] & (din_a[148] & din_b[149]))))

	.dataa(!din_a[149]),
	.datab(!din_b[148]),
	.datac(!din_a[148]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_93 ),
	.sharein(Xd_0__inst_mult_21_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_104 ),
	.cout(Xd_0__inst_mult_21_105 ),
	.shareout(Xd_0__inst_mult_21_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_33 (
// Equation(s):
// Xd_0__inst_mult_18_104  = SUM(( (!din_a[128] & (((din_a[127] & din_b[128])))) # (din_a[128] & (!din_b[127] $ (((!din_a[127]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_18_94  ) + ( Xd_0__inst_mult_18_93  ))
// Xd_0__inst_mult_18_105  = CARRY(( (!din_a[128] & (((din_a[127] & din_b[128])))) # (din_a[128] & (!din_b[127] $ (((!din_a[127]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_18_94  ) + ( Xd_0__inst_mult_18_93  ))
// Xd_0__inst_mult_18_106  = SHARE((din_a[128] & (din_b[127] & (din_a[127] & din_b[128]))))

	.dataa(!din_a[128]),
	.datab(!din_b[127]),
	.datac(!din_a[127]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_93 ),
	.sharein(Xd_0__inst_mult_18_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_104 ),
	.cout(Xd_0__inst_mult_18_105 ),
	.shareout(Xd_0__inst_mult_18_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_33 (
// Equation(s):
// Xd_0__inst_mult_19_104  = SUM(( (!din_a[135] & (((din_a[134] & din_b[135])))) # (din_a[135] & (!din_b[134] $ (((!din_a[134]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_19_94  ) + ( Xd_0__inst_mult_19_93  ))
// Xd_0__inst_mult_19_105  = CARRY(( (!din_a[135] & (((din_a[134] & din_b[135])))) # (din_a[135] & (!din_b[134] $ (((!din_a[134]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_19_94  ) + ( Xd_0__inst_mult_19_93  ))
// Xd_0__inst_mult_19_106  = SHARE((din_a[135] & (din_b[134] & (din_a[134] & din_b[135]))))

	.dataa(!din_a[135]),
	.datab(!din_b[134]),
	.datac(!din_a[134]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_93 ),
	.sharein(Xd_0__inst_mult_19_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_104 ),
	.cout(Xd_0__inst_mult_19_105 ),
	.shareout(Xd_0__inst_mult_19_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_33 (
// Equation(s):
// Xd_0__inst_mult_16_104  = SUM(( (!din_a[114] & (((din_a[113] & din_b[114])))) # (din_a[114] & (!din_b[113] $ (((!din_a[113]) # (!din_b[114]))))) ) + ( Xd_0__inst_mult_16_94  ) + ( Xd_0__inst_mult_16_93  ))
// Xd_0__inst_mult_16_105  = CARRY(( (!din_a[114] & (((din_a[113] & din_b[114])))) # (din_a[114] & (!din_b[113] $ (((!din_a[113]) # (!din_b[114]))))) ) + ( Xd_0__inst_mult_16_94  ) + ( Xd_0__inst_mult_16_93  ))
// Xd_0__inst_mult_16_106  = SHARE((din_a[114] & (din_b[113] & (din_a[113] & din_b[114]))))

	.dataa(!din_a[114]),
	.datab(!din_b[113]),
	.datac(!din_a[113]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_93 ),
	.sharein(Xd_0__inst_mult_16_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_104 ),
	.cout(Xd_0__inst_mult_16_105 ),
	.shareout(Xd_0__inst_mult_16_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_33 (
// Equation(s):
// Xd_0__inst_mult_17_104  = SUM(( (!din_a[121] & (((din_a[120] & din_b[121])))) # (din_a[121] & (!din_b[120] $ (((!din_a[120]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_17_94  ) + ( Xd_0__inst_mult_17_93  ))
// Xd_0__inst_mult_17_105  = CARRY(( (!din_a[121] & (((din_a[120] & din_b[121])))) # (din_a[121] & (!din_b[120] $ (((!din_a[120]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_17_94  ) + ( Xd_0__inst_mult_17_93  ))
// Xd_0__inst_mult_17_106  = SHARE((din_a[121] & (din_b[120] & (din_a[120] & din_b[121]))))

	.dataa(!din_a[121]),
	.datab(!din_b[120]),
	.datac(!din_a[120]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_93 ),
	.sharein(Xd_0__inst_mult_17_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_104 ),
	.cout(Xd_0__inst_mult_17_105 ),
	.shareout(Xd_0__inst_mult_17_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_33 (
// Equation(s):
// Xd_0__inst_mult_14_104  = SUM(( (!din_a[100] & (((din_a[99] & din_b[100])))) # (din_a[100] & (!din_b[99] $ (((!din_a[99]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_14_94  ) + ( Xd_0__inst_mult_14_93  ))
// Xd_0__inst_mult_14_105  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[100])))) # (din_a[100] & (!din_b[99] $ (((!din_a[99]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_14_94  ) + ( Xd_0__inst_mult_14_93  ))
// Xd_0__inst_mult_14_106  = SHARE((din_a[100] & (din_b[99] & (din_a[99] & din_b[100]))))

	.dataa(!din_a[100]),
	.datab(!din_b[99]),
	.datac(!din_a[99]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_93 ),
	.sharein(Xd_0__inst_mult_14_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_104 ),
	.cout(Xd_0__inst_mult_14_105 ),
	.shareout(Xd_0__inst_mult_14_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_33 (
// Equation(s):
// Xd_0__inst_mult_15_104  = SUM(( (!din_a[107] & (((din_a[106] & din_b[107])))) # (din_a[107] & (!din_b[106] $ (((!din_a[106]) # (!din_b[107]))))) ) + ( Xd_0__inst_mult_15_94  ) + ( Xd_0__inst_mult_15_93  ))
// Xd_0__inst_mult_15_105  = CARRY(( (!din_a[107] & (((din_a[106] & din_b[107])))) # (din_a[107] & (!din_b[106] $ (((!din_a[106]) # (!din_b[107]))))) ) + ( Xd_0__inst_mult_15_94  ) + ( Xd_0__inst_mult_15_93  ))
// Xd_0__inst_mult_15_106  = SHARE((din_a[107] & (din_b[106] & (din_a[106] & din_b[107]))))

	.dataa(!din_a[107]),
	.datab(!din_b[106]),
	.datac(!din_a[106]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_93 ),
	.sharein(Xd_0__inst_mult_15_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_104 ),
	.cout(Xd_0__inst_mult_15_105 ),
	.shareout(Xd_0__inst_mult_15_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_33 (
// Equation(s):
// Xd_0__inst_mult_12_104  = SUM(( (!din_a[86] & (((din_a[85] & din_b[86])))) # (din_a[86] & (!din_b[85] $ (((!din_a[85]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_12_94  ) + ( Xd_0__inst_mult_12_93  ))
// Xd_0__inst_mult_12_105  = CARRY(( (!din_a[86] & (((din_a[85] & din_b[86])))) # (din_a[86] & (!din_b[85] $ (((!din_a[85]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_12_94  ) + ( Xd_0__inst_mult_12_93  ))
// Xd_0__inst_mult_12_106  = SHARE((din_a[86] & (din_b[85] & (din_a[85] & din_b[86]))))

	.dataa(!din_a[86]),
	.datab(!din_b[85]),
	.datac(!din_a[85]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_93 ),
	.sharein(Xd_0__inst_mult_12_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_104 ),
	.cout(Xd_0__inst_mult_12_105 ),
	.shareout(Xd_0__inst_mult_12_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_33 (
// Equation(s):
// Xd_0__inst_mult_13_104  = SUM(( (!din_a[93] & (((din_a[92] & din_b[93])))) # (din_a[93] & (!din_b[92] $ (((!din_a[92]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_13_94  ) + ( Xd_0__inst_mult_13_93  ))
// Xd_0__inst_mult_13_105  = CARRY(( (!din_a[93] & (((din_a[92] & din_b[93])))) # (din_a[93] & (!din_b[92] $ (((!din_a[92]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_13_94  ) + ( Xd_0__inst_mult_13_93  ))
// Xd_0__inst_mult_13_106  = SHARE((din_a[93] & (din_b[92] & (din_a[92] & din_b[93]))))

	.dataa(!din_a[93]),
	.datab(!din_b[92]),
	.datac(!din_a[92]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_93 ),
	.sharein(Xd_0__inst_mult_13_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_104 ),
	.cout(Xd_0__inst_mult_13_105 ),
	.shareout(Xd_0__inst_mult_13_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_33 (
// Equation(s):
// Xd_0__inst_mult_10_104  = SUM(( (!din_a[72] & (((din_a[71] & din_b[72])))) # (din_a[72] & (!din_b[71] $ (((!din_a[71]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_10_94  ) + ( Xd_0__inst_mult_10_93  ))
// Xd_0__inst_mult_10_105  = CARRY(( (!din_a[72] & (((din_a[71] & din_b[72])))) # (din_a[72] & (!din_b[71] $ (((!din_a[71]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_10_94  ) + ( Xd_0__inst_mult_10_93  ))
// Xd_0__inst_mult_10_106  = SHARE((din_a[72] & (din_b[71] & (din_a[71] & din_b[72]))))

	.dataa(!din_a[72]),
	.datab(!din_b[71]),
	.datac(!din_a[71]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_93 ),
	.sharein(Xd_0__inst_mult_10_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_104 ),
	.cout(Xd_0__inst_mult_10_105 ),
	.shareout(Xd_0__inst_mult_10_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_33 (
// Equation(s):
// Xd_0__inst_mult_11_104  = SUM(( (!din_a[79] & (((din_a[78] & din_b[79])))) # (din_a[79] & (!din_b[78] $ (((!din_a[78]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_11_94  ) + ( Xd_0__inst_mult_11_93  ))
// Xd_0__inst_mult_11_105  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[79])))) # (din_a[79] & (!din_b[78] $ (((!din_a[78]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_11_94  ) + ( Xd_0__inst_mult_11_93  ))
// Xd_0__inst_mult_11_106  = SHARE((din_a[79] & (din_b[78] & (din_a[78] & din_b[79]))))

	.dataa(!din_a[79]),
	.datab(!din_b[78]),
	.datac(!din_a[78]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_93 ),
	.sharein(Xd_0__inst_mult_11_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_104 ),
	.cout(Xd_0__inst_mult_11_105 ),
	.shareout(Xd_0__inst_mult_11_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_33 (
// Equation(s):
// Xd_0__inst_mult_8_104  = SUM(( (!din_a[58] & (((din_a[57] & din_b[58])))) # (din_a[58] & (!din_b[57] $ (((!din_a[57]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_8_94  ) + ( Xd_0__inst_mult_8_93  ))
// Xd_0__inst_mult_8_105  = CARRY(( (!din_a[58] & (((din_a[57] & din_b[58])))) # (din_a[58] & (!din_b[57] $ (((!din_a[57]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_8_94  ) + ( Xd_0__inst_mult_8_93  ))
// Xd_0__inst_mult_8_106  = SHARE((din_a[58] & (din_b[57] & (din_a[57] & din_b[58]))))

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(!din_a[57]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_93 ),
	.sharein(Xd_0__inst_mult_8_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_104 ),
	.cout(Xd_0__inst_mult_8_105 ),
	.shareout(Xd_0__inst_mult_8_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_33 (
// Equation(s):
// Xd_0__inst_mult_9_104  = SUM(( (!din_a[65] & (((din_a[64] & din_b[65])))) # (din_a[65] & (!din_b[64] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_9_94  ) + ( Xd_0__inst_mult_9_93  ))
// Xd_0__inst_mult_9_105  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[65])))) # (din_a[65] & (!din_b[64] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_9_94  ) + ( Xd_0__inst_mult_9_93  ))
// Xd_0__inst_mult_9_106  = SHARE((din_a[65] & (din_b[64] & (din_a[64] & din_b[65]))))

	.dataa(!din_a[65]),
	.datab(!din_b[64]),
	.datac(!din_a[64]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_93 ),
	.sharein(Xd_0__inst_mult_9_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_104 ),
	.cout(Xd_0__inst_mult_9_105 ),
	.shareout(Xd_0__inst_mult_9_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_33 (
// Equation(s):
// Xd_0__inst_mult_6_104  = SUM(( (!din_a[44] & (((din_a[43] & din_b[44])))) # (din_a[44] & (!din_b[43] $ (((!din_a[43]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_6_94  ) + ( Xd_0__inst_mult_6_93  ))
// Xd_0__inst_mult_6_105  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[44])))) # (din_a[44] & (!din_b[43] $ (((!din_a[43]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_6_94  ) + ( Xd_0__inst_mult_6_93  ))
// Xd_0__inst_mult_6_106  = SHARE((din_a[44] & (din_b[43] & (din_a[43] & din_b[44]))))

	.dataa(!din_a[44]),
	.datab(!din_b[43]),
	.datac(!din_a[43]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_93 ),
	.sharein(Xd_0__inst_mult_6_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_104 ),
	.cout(Xd_0__inst_mult_6_105 ),
	.shareout(Xd_0__inst_mult_6_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_33 (
// Equation(s):
// Xd_0__inst_mult_7_104  = SUM(( (!din_a[51] & (((din_a[50] & din_b[51])))) # (din_a[51] & (!din_b[50] $ (((!din_a[50]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_7_94  ) + ( Xd_0__inst_mult_7_93  ))
// Xd_0__inst_mult_7_105  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[51])))) # (din_a[51] & (!din_b[50] $ (((!din_a[50]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_7_94  ) + ( Xd_0__inst_mult_7_93  ))
// Xd_0__inst_mult_7_106  = SHARE((din_a[51] & (din_b[50] & (din_a[50] & din_b[51]))))

	.dataa(!din_a[51]),
	.datab(!din_b[50]),
	.datac(!din_a[50]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_93 ),
	.sharein(Xd_0__inst_mult_7_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_104 ),
	.cout(Xd_0__inst_mult_7_105 ),
	.shareout(Xd_0__inst_mult_7_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_33 (
// Equation(s):
// Xd_0__inst_mult_4_104  = SUM(( (!din_a[30] & (((din_a[29] & din_b[30])))) # (din_a[30] & (!din_b[29] $ (((!din_a[29]) # (!din_b[30]))))) ) + ( Xd_0__inst_mult_4_94  ) + ( Xd_0__inst_mult_4_93  ))
// Xd_0__inst_mult_4_105  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[30])))) # (din_a[30] & (!din_b[29] $ (((!din_a[29]) # (!din_b[30]))))) ) + ( Xd_0__inst_mult_4_94  ) + ( Xd_0__inst_mult_4_93  ))
// Xd_0__inst_mult_4_106  = SHARE((din_a[30] & (din_b[29] & (din_a[29] & din_b[30]))))

	.dataa(!din_a[30]),
	.datab(!din_b[29]),
	.datac(!din_a[29]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_93 ),
	.sharein(Xd_0__inst_mult_4_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_104 ),
	.cout(Xd_0__inst_mult_4_105 ),
	.shareout(Xd_0__inst_mult_4_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_33 (
// Equation(s):
// Xd_0__inst_mult_5_104  = SUM(( (!din_a[37] & (((din_a[36] & din_b[37])))) # (din_a[37] & (!din_b[36] $ (((!din_a[36]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_5_94  ) + ( Xd_0__inst_mult_5_93  ))
// Xd_0__inst_mult_5_105  = CARRY(( (!din_a[37] & (((din_a[36] & din_b[37])))) # (din_a[37] & (!din_b[36] $ (((!din_a[36]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_5_94  ) + ( Xd_0__inst_mult_5_93  ))
// Xd_0__inst_mult_5_106  = SHARE((din_a[37] & (din_b[36] & (din_a[36] & din_b[37]))))

	.dataa(!din_a[37]),
	.datab(!din_b[36]),
	.datac(!din_a[36]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_93 ),
	.sharein(Xd_0__inst_mult_5_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_104 ),
	.cout(Xd_0__inst_mult_5_105 ),
	.shareout(Xd_0__inst_mult_5_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_33 (
// Equation(s):
// Xd_0__inst_mult_2_104  = SUM(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_2_94  ) + ( Xd_0__inst_mult_2_93  ))
// Xd_0__inst_mult_2_105  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_2_94  ) + ( Xd_0__inst_mult_2_93  ))
// Xd_0__inst_mult_2_106  = SHARE((din_a[16] & (din_b[15] & (din_a[15] & din_b[16]))))

	.dataa(!din_a[16]),
	.datab(!din_b[15]),
	.datac(!din_a[15]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_93 ),
	.sharein(Xd_0__inst_mult_2_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_104 ),
	.cout(Xd_0__inst_mult_2_105 ),
	.shareout(Xd_0__inst_mult_2_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_33 (
// Equation(s):
// Xd_0__inst_mult_3_104  = SUM(( (!din_a[23] & (((din_a[22] & din_b[23])))) # (din_a[23] & (!din_b[22] $ (((!din_a[22]) # (!din_b[23]))))) ) + ( Xd_0__inst_mult_3_94  ) + ( Xd_0__inst_mult_3_93  ))
// Xd_0__inst_mult_3_105  = CARRY(( (!din_a[23] & (((din_a[22] & din_b[23])))) # (din_a[23] & (!din_b[22] $ (((!din_a[22]) # (!din_b[23]))))) ) + ( Xd_0__inst_mult_3_94  ) + ( Xd_0__inst_mult_3_93  ))
// Xd_0__inst_mult_3_106  = SHARE((din_a[23] & (din_b[22] & (din_a[22] & din_b[23]))))

	.dataa(!din_a[23]),
	.datab(!din_b[22]),
	.datac(!din_a[22]),
	.datad(!din_b[23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_93 ),
	.sharein(Xd_0__inst_mult_3_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_104 ),
	.cout(Xd_0__inst_mult_3_105 ),
	.shareout(Xd_0__inst_mult_3_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_33 (
// Equation(s):
// Xd_0__inst_mult_0_104  = SUM(( (!din_a[2] & (((din_a[1] & din_b[2])))) # (din_a[2] & (!din_b[1] $ (((!din_a[1]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_94  ) + ( Xd_0__inst_mult_0_93  ))
// Xd_0__inst_mult_0_105  = CARRY(( (!din_a[2] & (((din_a[1] & din_b[2])))) # (din_a[2] & (!din_b[1] $ (((!din_a[1]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_94  ) + ( Xd_0__inst_mult_0_93  ))
// Xd_0__inst_mult_0_106  = SHARE((din_a[2] & (din_b[1] & (din_a[1] & din_b[2]))))

	.dataa(!din_a[2]),
	.datab(!din_b[1]),
	.datac(!din_a[1]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_93 ),
	.sharein(Xd_0__inst_mult_0_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_104 ),
	.cout(Xd_0__inst_mult_0_105 ),
	.shareout(Xd_0__inst_mult_0_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_33 (
// Equation(s):
// Xd_0__inst_mult_1_104  = SUM(( (!din_a[9] & (((din_a[8] & din_b[9])))) # (din_a[9] & (!din_b[8] $ (((!din_a[8]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_94  ) + ( Xd_0__inst_mult_1_93  ))
// Xd_0__inst_mult_1_105  = CARRY(( (!din_a[9] & (((din_a[8] & din_b[9])))) # (din_a[9] & (!din_b[8] $ (((!din_a[8]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_94  ) + ( Xd_0__inst_mult_1_93  ))
// Xd_0__inst_mult_1_106  = SHARE((din_a[9] & (din_b[8] & (din_a[8] & din_b[9]))))

	.dataa(!din_a[9]),
	.datab(!din_b[8]),
	.datac(!din_a[8]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_93 ),
	.sharein(Xd_0__inst_mult_1_94 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_104 ),
	.cout(Xd_0__inst_mult_1_105 ),
	.shareout(Xd_0__inst_mult_1_106 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_34 (
// Equation(s):
// Xd_0__inst_mult_28_108  = SUM(( (din_a[199] & din_b[197]) ) + ( Xd_0__inst_mult_28_106  ) + ( Xd_0__inst_mult_28_105  ))
// Xd_0__inst_mult_28_109  = CARRY(( (din_a[199] & din_b[197]) ) + ( Xd_0__inst_mult_28_106  ) + ( Xd_0__inst_mult_28_105  ))
// Xd_0__inst_mult_28_110  = SHARE((din_a[199] & din_b[198]))

	.dataa(!din_a[199]),
	.datab(!din_b[197]),
	.datac(!din_b[198]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_105 ),
	.sharein(Xd_0__inst_mult_28_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_108 ),
	.cout(Xd_0__inst_mult_28_109 ),
	.shareout(Xd_0__inst_mult_28_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_35 (
// Equation(s):
// Xd_0__inst_mult_28_112  = SUM(( (din_a[196] & din_b[200]) ) + ( Xd_0__inst_mult_28_158  ) + ( Xd_0__inst_mult_28_157  ))
// Xd_0__inst_mult_28_113  = CARRY(( (din_a[196] & din_b[200]) ) + ( Xd_0__inst_mult_28_158  ) + ( Xd_0__inst_mult_28_157  ))
// Xd_0__inst_mult_28_114  = SHARE((din_a[198] & din_b[199]))

	.dataa(!din_a[196]),
	.datab(!din_b[200]),
	.datac(!din_a[198]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_157 ),
	.sharein(Xd_0__inst_mult_28_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_112 ),
	.cout(Xd_0__inst_mult_28_113 ),
	.shareout(Xd_0__inst_mult_28_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_34 (
// Equation(s):
// Xd_0__inst_mult_29_108  = SUM(( (din_a[206] & din_b[204]) ) + ( Xd_0__inst_mult_29_106  ) + ( Xd_0__inst_mult_29_105  ))
// Xd_0__inst_mult_29_109  = CARRY(( (din_a[206] & din_b[204]) ) + ( Xd_0__inst_mult_29_106  ) + ( Xd_0__inst_mult_29_105  ))
// Xd_0__inst_mult_29_110  = SHARE((din_a[206] & din_b[205]))

	.dataa(!din_a[206]),
	.datab(!din_b[204]),
	.datac(!din_b[205]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_105 ),
	.sharein(Xd_0__inst_mult_29_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_108 ),
	.cout(Xd_0__inst_mult_29_109 ),
	.shareout(Xd_0__inst_mult_29_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_35 (
// Equation(s):
// Xd_0__inst_mult_29_112  = SUM(( (din_a[203] & din_b[207]) ) + ( Xd_0__inst_mult_29_158  ) + ( Xd_0__inst_mult_29_157  ))
// Xd_0__inst_mult_29_113  = CARRY(( (din_a[203] & din_b[207]) ) + ( Xd_0__inst_mult_29_158  ) + ( Xd_0__inst_mult_29_157  ))
// Xd_0__inst_mult_29_114  = SHARE((din_a[205] & din_b[206]))

	.dataa(!din_a[203]),
	.datab(!din_b[207]),
	.datac(!din_a[205]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_157 ),
	.sharein(Xd_0__inst_mult_29_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_112 ),
	.cout(Xd_0__inst_mult_29_113 ),
	.shareout(Xd_0__inst_mult_29_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_34 (
// Equation(s):
// Xd_0__inst_mult_26_108  = SUM(( (din_a[185] & din_b[183]) ) + ( Xd_0__inst_mult_26_106  ) + ( Xd_0__inst_mult_26_105  ))
// Xd_0__inst_mult_26_109  = CARRY(( (din_a[185] & din_b[183]) ) + ( Xd_0__inst_mult_26_106  ) + ( Xd_0__inst_mult_26_105  ))
// Xd_0__inst_mult_26_110  = SHARE((din_a[185] & din_b[184]))

	.dataa(!din_a[185]),
	.datab(!din_b[183]),
	.datac(!din_b[184]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_105 ),
	.sharein(Xd_0__inst_mult_26_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_108 ),
	.cout(Xd_0__inst_mult_26_109 ),
	.shareout(Xd_0__inst_mult_26_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_35 (
// Equation(s):
// Xd_0__inst_mult_26_112  = SUM(( (din_a[182] & din_b[186]) ) + ( Xd_0__inst_mult_26_158  ) + ( Xd_0__inst_mult_26_157  ))
// Xd_0__inst_mult_26_113  = CARRY(( (din_a[182] & din_b[186]) ) + ( Xd_0__inst_mult_26_158  ) + ( Xd_0__inst_mult_26_157  ))
// Xd_0__inst_mult_26_114  = SHARE((din_a[184] & din_b[185]))

	.dataa(!din_a[182]),
	.datab(!din_b[186]),
	.datac(!din_a[184]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_157 ),
	.sharein(Xd_0__inst_mult_26_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_112 ),
	.cout(Xd_0__inst_mult_26_113 ),
	.shareout(Xd_0__inst_mult_26_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_34 (
// Equation(s):
// Xd_0__inst_mult_27_108  = SUM(( (din_a[192] & din_b[190]) ) + ( Xd_0__inst_mult_27_106  ) + ( Xd_0__inst_mult_27_105  ))
// Xd_0__inst_mult_27_109  = CARRY(( (din_a[192] & din_b[190]) ) + ( Xd_0__inst_mult_27_106  ) + ( Xd_0__inst_mult_27_105  ))
// Xd_0__inst_mult_27_110  = SHARE((din_a[192] & din_b[191]))

	.dataa(!din_a[192]),
	.datab(!din_b[190]),
	.datac(!din_b[191]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_105 ),
	.sharein(Xd_0__inst_mult_27_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_108 ),
	.cout(Xd_0__inst_mult_27_109 ),
	.shareout(Xd_0__inst_mult_27_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_35 (
// Equation(s):
// Xd_0__inst_mult_27_112  = SUM(( (din_a[189] & din_b[193]) ) + ( Xd_0__inst_mult_27_158  ) + ( Xd_0__inst_mult_27_157  ))
// Xd_0__inst_mult_27_113  = CARRY(( (din_a[189] & din_b[193]) ) + ( Xd_0__inst_mult_27_158  ) + ( Xd_0__inst_mult_27_157  ))
// Xd_0__inst_mult_27_114  = SHARE((din_a[191] & din_b[192]))

	.dataa(!din_a[189]),
	.datab(!din_b[193]),
	.datac(!din_a[191]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_157 ),
	.sharein(Xd_0__inst_mult_27_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_112 ),
	.cout(Xd_0__inst_mult_27_113 ),
	.shareout(Xd_0__inst_mult_27_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_34 (
// Equation(s):
// Xd_0__inst_mult_24_108  = SUM(( (din_a[171] & din_b[169]) ) + ( Xd_0__inst_mult_24_106  ) + ( Xd_0__inst_mult_24_105  ))
// Xd_0__inst_mult_24_109  = CARRY(( (din_a[171] & din_b[169]) ) + ( Xd_0__inst_mult_24_106  ) + ( Xd_0__inst_mult_24_105  ))
// Xd_0__inst_mult_24_110  = SHARE((din_a[171] & din_b[170]))

	.dataa(!din_a[171]),
	.datab(!din_b[169]),
	.datac(!din_b[170]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_105 ),
	.sharein(Xd_0__inst_mult_24_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_108 ),
	.cout(Xd_0__inst_mult_24_109 ),
	.shareout(Xd_0__inst_mult_24_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_35 (
// Equation(s):
// Xd_0__inst_mult_24_112  = SUM(( (din_a[168] & din_b[172]) ) + ( Xd_0__inst_mult_24_158  ) + ( Xd_0__inst_mult_24_157  ))
// Xd_0__inst_mult_24_113  = CARRY(( (din_a[168] & din_b[172]) ) + ( Xd_0__inst_mult_24_158  ) + ( Xd_0__inst_mult_24_157  ))
// Xd_0__inst_mult_24_114  = SHARE((din_a[170] & din_b[171]))

	.dataa(!din_a[168]),
	.datab(!din_b[172]),
	.datac(!din_a[170]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_157 ),
	.sharein(Xd_0__inst_mult_24_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_112 ),
	.cout(Xd_0__inst_mult_24_113 ),
	.shareout(Xd_0__inst_mult_24_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_35 (
// Equation(s):
// Xd_0__inst_mult_25_112  = SUM(( (din_a[178] & din_b[176]) ) + ( Xd_0__inst_mult_25_110  ) + ( Xd_0__inst_mult_25_109  ))
// Xd_0__inst_mult_25_113  = CARRY(( (din_a[178] & din_b[176]) ) + ( Xd_0__inst_mult_25_110  ) + ( Xd_0__inst_mult_25_109  ))
// Xd_0__inst_mult_25_114  = SHARE((din_a[178] & din_b[177]))

	.dataa(!din_a[178]),
	.datab(!din_b[176]),
	.datac(!din_b[177]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_109 ),
	.sharein(Xd_0__inst_mult_25_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_112 ),
	.cout(Xd_0__inst_mult_25_113 ),
	.shareout(Xd_0__inst_mult_25_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_36 (
// Equation(s):
// Xd_0__inst_mult_25_116  = SUM(( (din_a[175] & din_b[179]) ) + ( Xd_0__inst_mult_25_158  ) + ( Xd_0__inst_mult_25_157  ))
// Xd_0__inst_mult_25_117  = CARRY(( (din_a[175] & din_b[179]) ) + ( Xd_0__inst_mult_25_158  ) + ( Xd_0__inst_mult_25_157  ))
// Xd_0__inst_mult_25_118  = SHARE((din_a[177] & din_b[178]))

	.dataa(!din_a[175]),
	.datab(!din_b[179]),
	.datac(!din_a[177]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_157 ),
	.sharein(Xd_0__inst_mult_25_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_116 ),
	.cout(Xd_0__inst_mult_25_117 ),
	.shareout(Xd_0__inst_mult_25_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_35 (
// Equation(s):
// Xd_0__inst_mult_22_112  = SUM(( (din_a[157] & din_b[155]) ) + ( Xd_0__inst_mult_22_110  ) + ( Xd_0__inst_mult_22_109  ))
// Xd_0__inst_mult_22_113  = CARRY(( (din_a[157] & din_b[155]) ) + ( Xd_0__inst_mult_22_110  ) + ( Xd_0__inst_mult_22_109  ))
// Xd_0__inst_mult_22_114  = SHARE((din_a[157] & din_b[156]))

	.dataa(!din_a[157]),
	.datab(!din_b[155]),
	.datac(!din_b[156]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_109 ),
	.sharein(Xd_0__inst_mult_22_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_112 ),
	.cout(Xd_0__inst_mult_22_113 ),
	.shareout(Xd_0__inst_mult_22_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_36 (
// Equation(s):
// Xd_0__inst_mult_22_116  = SUM(( (din_a[154] & din_b[158]) ) + ( Xd_0__inst_mult_22_158  ) + ( Xd_0__inst_mult_22_157  ))
// Xd_0__inst_mult_22_117  = CARRY(( (din_a[154] & din_b[158]) ) + ( Xd_0__inst_mult_22_158  ) + ( Xd_0__inst_mult_22_157  ))
// Xd_0__inst_mult_22_118  = SHARE((din_a[156] & din_b[157]))

	.dataa(!din_a[154]),
	.datab(!din_b[158]),
	.datac(!din_a[156]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_157 ),
	.sharein(Xd_0__inst_mult_22_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_116 ),
	.cout(Xd_0__inst_mult_22_117 ),
	.shareout(Xd_0__inst_mult_22_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_34 (
// Equation(s):
// Xd_0__inst_mult_23_108  = SUM(( (din_a[164] & din_b[162]) ) + ( Xd_0__inst_mult_23_106  ) + ( Xd_0__inst_mult_23_105  ))
// Xd_0__inst_mult_23_109  = CARRY(( (din_a[164] & din_b[162]) ) + ( Xd_0__inst_mult_23_106  ) + ( Xd_0__inst_mult_23_105  ))
// Xd_0__inst_mult_23_110  = SHARE((din_a[164] & din_b[163]))

	.dataa(!din_a[164]),
	.datab(!din_b[162]),
	.datac(!din_b[163]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_105 ),
	.sharein(Xd_0__inst_mult_23_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_108 ),
	.cout(Xd_0__inst_mult_23_109 ),
	.shareout(Xd_0__inst_mult_23_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_35 (
// Equation(s):
// Xd_0__inst_mult_23_112  = SUM(( (din_a[161] & din_b[165]) ) + ( Xd_0__inst_mult_23_158  ) + ( Xd_0__inst_mult_23_157  ))
// Xd_0__inst_mult_23_113  = CARRY(( (din_a[161] & din_b[165]) ) + ( Xd_0__inst_mult_23_158  ) + ( Xd_0__inst_mult_23_157  ))
// Xd_0__inst_mult_23_114  = SHARE((din_a[163] & din_b[164]))

	.dataa(!din_a[161]),
	.datab(!din_b[165]),
	.datac(!din_a[163]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_157 ),
	.sharein(Xd_0__inst_mult_23_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_112 ),
	.cout(Xd_0__inst_mult_23_113 ),
	.shareout(Xd_0__inst_mult_23_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_34 (
// Equation(s):
// Xd_0__inst_mult_20_108  = SUM(( (din_a[143] & din_b[141]) ) + ( Xd_0__inst_mult_20_106  ) + ( Xd_0__inst_mult_20_105  ))
// Xd_0__inst_mult_20_109  = CARRY(( (din_a[143] & din_b[141]) ) + ( Xd_0__inst_mult_20_106  ) + ( Xd_0__inst_mult_20_105  ))
// Xd_0__inst_mult_20_110  = SHARE((din_a[143] & din_b[142]))

	.dataa(!din_a[143]),
	.datab(!din_b[141]),
	.datac(!din_b[142]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_105 ),
	.sharein(Xd_0__inst_mult_20_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_108 ),
	.cout(Xd_0__inst_mult_20_109 ),
	.shareout(Xd_0__inst_mult_20_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_35 (
// Equation(s):
// Xd_0__inst_mult_20_112  = SUM(( (din_a[140] & din_b[144]) ) + ( Xd_0__inst_mult_20_158  ) + ( Xd_0__inst_mult_20_157  ))
// Xd_0__inst_mult_20_113  = CARRY(( (din_a[140] & din_b[144]) ) + ( Xd_0__inst_mult_20_158  ) + ( Xd_0__inst_mult_20_157  ))
// Xd_0__inst_mult_20_114  = SHARE((din_a[142] & din_b[143]))

	.dataa(!din_a[140]),
	.datab(!din_b[144]),
	.datac(!din_a[142]),
	.datad(!din_b[143]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_157 ),
	.sharein(Xd_0__inst_mult_20_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_112 ),
	.cout(Xd_0__inst_mult_20_113 ),
	.shareout(Xd_0__inst_mult_20_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_34 (
// Equation(s):
// Xd_0__inst_mult_21_108  = SUM(( (din_a[150] & din_b[148]) ) + ( Xd_0__inst_mult_21_106  ) + ( Xd_0__inst_mult_21_105  ))
// Xd_0__inst_mult_21_109  = CARRY(( (din_a[150] & din_b[148]) ) + ( Xd_0__inst_mult_21_106  ) + ( Xd_0__inst_mult_21_105  ))
// Xd_0__inst_mult_21_110  = SHARE((din_a[150] & din_b[149]))

	.dataa(!din_a[150]),
	.datab(!din_b[148]),
	.datac(!din_b[149]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_105 ),
	.sharein(Xd_0__inst_mult_21_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_108 ),
	.cout(Xd_0__inst_mult_21_109 ),
	.shareout(Xd_0__inst_mult_21_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_35 (
// Equation(s):
// Xd_0__inst_mult_21_112  = SUM(( (din_a[147] & din_b[151]) ) + ( Xd_0__inst_mult_21_158  ) + ( Xd_0__inst_mult_21_157  ))
// Xd_0__inst_mult_21_113  = CARRY(( (din_a[147] & din_b[151]) ) + ( Xd_0__inst_mult_21_158  ) + ( Xd_0__inst_mult_21_157  ))
// Xd_0__inst_mult_21_114  = SHARE((din_a[149] & din_b[150]))

	.dataa(!din_a[147]),
	.datab(!din_b[151]),
	.datac(!din_a[149]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_157 ),
	.sharein(Xd_0__inst_mult_21_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_112 ),
	.cout(Xd_0__inst_mult_21_113 ),
	.shareout(Xd_0__inst_mult_21_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_34 (
// Equation(s):
// Xd_0__inst_mult_18_108  = SUM(( (din_a[129] & din_b[127]) ) + ( Xd_0__inst_mult_18_106  ) + ( Xd_0__inst_mult_18_105  ))
// Xd_0__inst_mult_18_109  = CARRY(( (din_a[129] & din_b[127]) ) + ( Xd_0__inst_mult_18_106  ) + ( Xd_0__inst_mult_18_105  ))
// Xd_0__inst_mult_18_110  = SHARE((din_a[129] & din_b[128]))

	.dataa(!din_a[129]),
	.datab(!din_b[127]),
	.datac(!din_b[128]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_105 ),
	.sharein(Xd_0__inst_mult_18_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_108 ),
	.cout(Xd_0__inst_mult_18_109 ),
	.shareout(Xd_0__inst_mult_18_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_35 (
// Equation(s):
// Xd_0__inst_mult_18_112  = SUM(( (din_a[126] & din_b[130]) ) + ( Xd_0__inst_mult_18_158  ) + ( Xd_0__inst_mult_18_157  ))
// Xd_0__inst_mult_18_113  = CARRY(( (din_a[126] & din_b[130]) ) + ( Xd_0__inst_mult_18_158  ) + ( Xd_0__inst_mult_18_157  ))
// Xd_0__inst_mult_18_114  = SHARE((din_a[128] & din_b[129]))

	.dataa(!din_a[126]),
	.datab(!din_b[130]),
	.datac(!din_a[128]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_157 ),
	.sharein(Xd_0__inst_mult_18_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_112 ),
	.cout(Xd_0__inst_mult_18_113 ),
	.shareout(Xd_0__inst_mult_18_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_34 (
// Equation(s):
// Xd_0__inst_mult_19_108  = SUM(( (din_a[136] & din_b[134]) ) + ( Xd_0__inst_mult_19_106  ) + ( Xd_0__inst_mult_19_105  ))
// Xd_0__inst_mult_19_109  = CARRY(( (din_a[136] & din_b[134]) ) + ( Xd_0__inst_mult_19_106  ) + ( Xd_0__inst_mult_19_105  ))
// Xd_0__inst_mult_19_110  = SHARE((din_a[136] & din_b[135]))

	.dataa(!din_a[136]),
	.datab(!din_b[134]),
	.datac(!din_b[135]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_105 ),
	.sharein(Xd_0__inst_mult_19_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_108 ),
	.cout(Xd_0__inst_mult_19_109 ),
	.shareout(Xd_0__inst_mult_19_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_35 (
// Equation(s):
// Xd_0__inst_mult_19_112  = SUM(( (din_a[133] & din_b[137]) ) + ( Xd_0__inst_mult_19_158  ) + ( Xd_0__inst_mult_19_157  ))
// Xd_0__inst_mult_19_113  = CARRY(( (din_a[133] & din_b[137]) ) + ( Xd_0__inst_mult_19_158  ) + ( Xd_0__inst_mult_19_157  ))
// Xd_0__inst_mult_19_114  = SHARE((din_a[135] & din_b[136]))

	.dataa(!din_a[133]),
	.datab(!din_b[137]),
	.datac(!din_a[135]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_157 ),
	.sharein(Xd_0__inst_mult_19_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_112 ),
	.cout(Xd_0__inst_mult_19_113 ),
	.shareout(Xd_0__inst_mult_19_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_46 (
// Equation(s):
// Xd_0__inst_mult_30_157  = CARRY(( (din_a[212] & din_b[212]) ) + ( Xd_0__inst_mult_30_162  ) + ( Xd_0__inst_mult_30_161  ))
// Xd_0__inst_mult_30_158  = SHARE((din_a[211] & din_b[213]))

	.dataa(!din_a[212]),
	.datab(!din_b[212]),
	.datac(!din_a[211]),
	.datad(!din_b[213]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_161 ),
	.sharein(Xd_0__inst_mult_30_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_157 ),
	.shareout(Xd_0__inst_mult_30_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_46 (
// Equation(s):
// Xd_0__inst_mult_31_157  = CARRY(( (din_a[219] & din_b[219]) ) + ( Xd_0__inst_mult_31_162  ) + ( Xd_0__inst_mult_31_161  ))
// Xd_0__inst_mult_31_158  = SHARE((din_a[218] & din_b[220]))

	.dataa(!din_a[219]),
	.datab(!din_b[219]),
	.datac(!din_a[218]),
	.datad(!din_b[220]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_161 ),
	.sharein(Xd_0__inst_mult_31_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_157 ),
	.shareout(Xd_0__inst_mult_31_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_34 (
// Equation(s):
// Xd_0__inst_mult_16_108  = SUM(( (din_a[115] & din_b[113]) ) + ( Xd_0__inst_mult_16_106  ) + ( Xd_0__inst_mult_16_105  ))
// Xd_0__inst_mult_16_109  = CARRY(( (din_a[115] & din_b[113]) ) + ( Xd_0__inst_mult_16_106  ) + ( Xd_0__inst_mult_16_105  ))
// Xd_0__inst_mult_16_110  = SHARE((din_a[115] & din_b[114]))

	.dataa(!din_a[115]),
	.datab(!din_b[113]),
	.datac(!din_b[114]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_105 ),
	.sharein(Xd_0__inst_mult_16_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_108 ),
	.cout(Xd_0__inst_mult_16_109 ),
	.shareout(Xd_0__inst_mult_16_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_35 (
// Equation(s):
// Xd_0__inst_mult_16_112  = SUM(( (din_a[112] & din_b[116]) ) + ( Xd_0__inst_mult_16_158  ) + ( Xd_0__inst_mult_16_157  ))
// Xd_0__inst_mult_16_113  = CARRY(( (din_a[112] & din_b[116]) ) + ( Xd_0__inst_mult_16_158  ) + ( Xd_0__inst_mult_16_157  ))
// Xd_0__inst_mult_16_114  = SHARE((din_a[114] & din_b[115]))

	.dataa(!din_a[112]),
	.datab(!din_b[116]),
	.datac(!din_a[114]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_157 ),
	.sharein(Xd_0__inst_mult_16_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_112 ),
	.cout(Xd_0__inst_mult_16_113 ),
	.shareout(Xd_0__inst_mult_16_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_34 (
// Equation(s):
// Xd_0__inst_mult_17_108  = SUM(( (din_a[122] & din_b[120]) ) + ( Xd_0__inst_mult_17_106  ) + ( Xd_0__inst_mult_17_105  ))
// Xd_0__inst_mult_17_109  = CARRY(( (din_a[122] & din_b[120]) ) + ( Xd_0__inst_mult_17_106  ) + ( Xd_0__inst_mult_17_105  ))
// Xd_0__inst_mult_17_110  = SHARE((din_a[122] & din_b[121]))

	.dataa(!din_a[122]),
	.datab(!din_b[120]),
	.datac(!din_b[121]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_105 ),
	.sharein(Xd_0__inst_mult_17_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_108 ),
	.cout(Xd_0__inst_mult_17_109 ),
	.shareout(Xd_0__inst_mult_17_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_35 (
// Equation(s):
// Xd_0__inst_mult_17_112  = SUM(( (din_a[119] & din_b[123]) ) + ( Xd_0__inst_mult_17_158  ) + ( Xd_0__inst_mult_17_157  ))
// Xd_0__inst_mult_17_113  = CARRY(( (din_a[119] & din_b[123]) ) + ( Xd_0__inst_mult_17_158  ) + ( Xd_0__inst_mult_17_157  ))
// Xd_0__inst_mult_17_114  = SHARE((din_a[121] & din_b[122]))

	.dataa(!din_a[119]),
	.datab(!din_b[123]),
	.datac(!din_a[121]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_157 ),
	.sharein(Xd_0__inst_mult_17_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_112 ),
	.cout(Xd_0__inst_mult_17_113 ),
	.shareout(Xd_0__inst_mult_17_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_34 (
// Equation(s):
// Xd_0__inst_mult_14_108  = SUM(( (din_a[101] & din_b[99]) ) + ( Xd_0__inst_mult_14_106  ) + ( Xd_0__inst_mult_14_105  ))
// Xd_0__inst_mult_14_109  = CARRY(( (din_a[101] & din_b[99]) ) + ( Xd_0__inst_mult_14_106  ) + ( Xd_0__inst_mult_14_105  ))
// Xd_0__inst_mult_14_110  = SHARE((din_a[101] & din_b[100]))

	.dataa(!din_a[101]),
	.datab(!din_b[99]),
	.datac(!din_b[100]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_105 ),
	.sharein(Xd_0__inst_mult_14_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_108 ),
	.cout(Xd_0__inst_mult_14_109 ),
	.shareout(Xd_0__inst_mult_14_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_35 (
// Equation(s):
// Xd_0__inst_mult_14_112  = SUM(( (din_a[98] & din_b[102]) ) + ( Xd_0__inst_mult_14_158  ) + ( Xd_0__inst_mult_14_157  ))
// Xd_0__inst_mult_14_113  = CARRY(( (din_a[98] & din_b[102]) ) + ( Xd_0__inst_mult_14_158  ) + ( Xd_0__inst_mult_14_157  ))
// Xd_0__inst_mult_14_114  = SHARE((din_a[100] & din_b[101]))

	.dataa(!din_a[98]),
	.datab(!din_b[102]),
	.datac(!din_a[100]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_157 ),
	.sharein(Xd_0__inst_mult_14_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_112 ),
	.cout(Xd_0__inst_mult_14_113 ),
	.shareout(Xd_0__inst_mult_14_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_34 (
// Equation(s):
// Xd_0__inst_mult_15_108  = SUM(( (din_a[108] & din_b[106]) ) + ( Xd_0__inst_mult_15_106  ) + ( Xd_0__inst_mult_15_105  ))
// Xd_0__inst_mult_15_109  = CARRY(( (din_a[108] & din_b[106]) ) + ( Xd_0__inst_mult_15_106  ) + ( Xd_0__inst_mult_15_105  ))
// Xd_0__inst_mult_15_110  = SHARE((din_a[108] & din_b[107]))

	.dataa(!din_a[108]),
	.datab(!din_b[106]),
	.datac(!din_b[107]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_105 ),
	.sharein(Xd_0__inst_mult_15_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_108 ),
	.cout(Xd_0__inst_mult_15_109 ),
	.shareout(Xd_0__inst_mult_15_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_35 (
// Equation(s):
// Xd_0__inst_mult_15_112  = SUM(( (din_a[105] & din_b[109]) ) + ( Xd_0__inst_mult_15_158  ) + ( Xd_0__inst_mult_15_157  ))
// Xd_0__inst_mult_15_113  = CARRY(( (din_a[105] & din_b[109]) ) + ( Xd_0__inst_mult_15_158  ) + ( Xd_0__inst_mult_15_157  ))
// Xd_0__inst_mult_15_114  = SHARE((din_a[107] & din_b[108]))

	.dataa(!din_a[105]),
	.datab(!din_b[109]),
	.datac(!din_a[107]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_157 ),
	.sharein(Xd_0__inst_mult_15_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_112 ),
	.cout(Xd_0__inst_mult_15_113 ),
	.shareout(Xd_0__inst_mult_15_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_34 (
// Equation(s):
// Xd_0__inst_mult_12_108  = SUM(( (din_a[87] & din_b[85]) ) + ( Xd_0__inst_mult_12_106  ) + ( Xd_0__inst_mult_12_105  ))
// Xd_0__inst_mult_12_109  = CARRY(( (din_a[87] & din_b[85]) ) + ( Xd_0__inst_mult_12_106  ) + ( Xd_0__inst_mult_12_105  ))
// Xd_0__inst_mult_12_110  = SHARE((din_a[87] & din_b[86]))

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(!din_b[86]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_105 ),
	.sharein(Xd_0__inst_mult_12_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_108 ),
	.cout(Xd_0__inst_mult_12_109 ),
	.shareout(Xd_0__inst_mult_12_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_35 (
// Equation(s):
// Xd_0__inst_mult_12_112  = SUM(( (din_a[84] & din_b[88]) ) + ( Xd_0__inst_mult_12_158  ) + ( Xd_0__inst_mult_12_157  ))
// Xd_0__inst_mult_12_113  = CARRY(( (din_a[84] & din_b[88]) ) + ( Xd_0__inst_mult_12_158  ) + ( Xd_0__inst_mult_12_157  ))
// Xd_0__inst_mult_12_114  = SHARE((din_a[86] & din_b[87]))

	.dataa(!din_a[84]),
	.datab(!din_b[88]),
	.datac(!din_a[86]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_157 ),
	.sharein(Xd_0__inst_mult_12_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_112 ),
	.cout(Xd_0__inst_mult_12_113 ),
	.shareout(Xd_0__inst_mult_12_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_34 (
// Equation(s):
// Xd_0__inst_mult_13_108  = SUM(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_13_106  ) + ( Xd_0__inst_mult_13_105  ))
// Xd_0__inst_mult_13_109  = CARRY(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_13_106  ) + ( Xd_0__inst_mult_13_105  ))
// Xd_0__inst_mult_13_110  = SHARE((din_a[94] & din_b[93]))

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(!din_b[93]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_105 ),
	.sharein(Xd_0__inst_mult_13_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_108 ),
	.cout(Xd_0__inst_mult_13_109 ),
	.shareout(Xd_0__inst_mult_13_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_35 (
// Equation(s):
// Xd_0__inst_mult_13_112  = SUM(( (din_a[91] & din_b[95]) ) + ( Xd_0__inst_mult_13_158  ) + ( Xd_0__inst_mult_13_157  ))
// Xd_0__inst_mult_13_113  = CARRY(( (din_a[91] & din_b[95]) ) + ( Xd_0__inst_mult_13_158  ) + ( Xd_0__inst_mult_13_157  ))
// Xd_0__inst_mult_13_114  = SHARE((din_a[93] & din_b[94]))

	.dataa(!din_a[91]),
	.datab(!din_b[95]),
	.datac(!din_a[93]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_157 ),
	.sharein(Xd_0__inst_mult_13_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_112 ),
	.cout(Xd_0__inst_mult_13_113 ),
	.shareout(Xd_0__inst_mult_13_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_34 (
// Equation(s):
// Xd_0__inst_mult_10_108  = SUM(( (din_a[73] & din_b[71]) ) + ( Xd_0__inst_mult_10_106  ) + ( Xd_0__inst_mult_10_105  ))
// Xd_0__inst_mult_10_109  = CARRY(( (din_a[73] & din_b[71]) ) + ( Xd_0__inst_mult_10_106  ) + ( Xd_0__inst_mult_10_105  ))
// Xd_0__inst_mult_10_110  = SHARE((din_a[73] & din_b[72]))

	.dataa(!din_a[73]),
	.datab(!din_b[71]),
	.datac(!din_b[72]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_105 ),
	.sharein(Xd_0__inst_mult_10_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_108 ),
	.cout(Xd_0__inst_mult_10_109 ),
	.shareout(Xd_0__inst_mult_10_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_35 (
// Equation(s):
// Xd_0__inst_mult_10_112  = SUM(( (din_a[70] & din_b[74]) ) + ( Xd_0__inst_mult_10_158  ) + ( Xd_0__inst_mult_10_157  ))
// Xd_0__inst_mult_10_113  = CARRY(( (din_a[70] & din_b[74]) ) + ( Xd_0__inst_mult_10_158  ) + ( Xd_0__inst_mult_10_157  ))
// Xd_0__inst_mult_10_114  = SHARE((din_a[72] & din_b[73]))

	.dataa(!din_a[70]),
	.datab(!din_b[74]),
	.datac(!din_a[72]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_157 ),
	.sharein(Xd_0__inst_mult_10_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_112 ),
	.cout(Xd_0__inst_mult_10_113 ),
	.shareout(Xd_0__inst_mult_10_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_34 (
// Equation(s):
// Xd_0__inst_mult_11_108  = SUM(( (din_a[80] & din_b[78]) ) + ( Xd_0__inst_mult_11_106  ) + ( Xd_0__inst_mult_11_105  ))
// Xd_0__inst_mult_11_109  = CARRY(( (din_a[80] & din_b[78]) ) + ( Xd_0__inst_mult_11_106  ) + ( Xd_0__inst_mult_11_105  ))
// Xd_0__inst_mult_11_110  = SHARE((din_a[80] & din_b[79]))

	.dataa(!din_a[80]),
	.datab(!din_b[78]),
	.datac(!din_b[79]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_105 ),
	.sharein(Xd_0__inst_mult_11_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_108 ),
	.cout(Xd_0__inst_mult_11_109 ),
	.shareout(Xd_0__inst_mult_11_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_35 (
// Equation(s):
// Xd_0__inst_mult_11_112  = SUM(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_11_158  ) + ( Xd_0__inst_mult_11_157  ))
// Xd_0__inst_mult_11_113  = CARRY(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_11_158  ) + ( Xd_0__inst_mult_11_157  ))
// Xd_0__inst_mult_11_114  = SHARE((din_a[79] & din_b[80]))

	.dataa(!din_a[77]),
	.datab(!din_b[81]),
	.datac(!din_a[79]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_157 ),
	.sharein(Xd_0__inst_mult_11_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_112 ),
	.cout(Xd_0__inst_mult_11_113 ),
	.shareout(Xd_0__inst_mult_11_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_34 (
// Equation(s):
// Xd_0__inst_mult_8_108  = SUM(( (din_a[59] & din_b[57]) ) + ( Xd_0__inst_mult_8_106  ) + ( Xd_0__inst_mult_8_105  ))
// Xd_0__inst_mult_8_109  = CARRY(( (din_a[59] & din_b[57]) ) + ( Xd_0__inst_mult_8_106  ) + ( Xd_0__inst_mult_8_105  ))
// Xd_0__inst_mult_8_110  = SHARE((din_a[59] & din_b[58]))

	.dataa(!din_a[59]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_105 ),
	.sharein(Xd_0__inst_mult_8_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_108 ),
	.cout(Xd_0__inst_mult_8_109 ),
	.shareout(Xd_0__inst_mult_8_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_35 (
// Equation(s):
// Xd_0__inst_mult_8_112  = SUM(( (din_a[56] & din_b[60]) ) + ( Xd_0__inst_mult_8_158  ) + ( Xd_0__inst_mult_8_157  ))
// Xd_0__inst_mult_8_113  = CARRY(( (din_a[56] & din_b[60]) ) + ( Xd_0__inst_mult_8_158  ) + ( Xd_0__inst_mult_8_157  ))
// Xd_0__inst_mult_8_114  = SHARE((din_a[58] & din_b[59]))

	.dataa(!din_a[56]),
	.datab(!din_b[60]),
	.datac(!din_a[58]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_157 ),
	.sharein(Xd_0__inst_mult_8_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_112 ),
	.cout(Xd_0__inst_mult_8_113 ),
	.shareout(Xd_0__inst_mult_8_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_34 (
// Equation(s):
// Xd_0__inst_mult_9_108  = SUM(( (din_a[66] & din_b[64]) ) + ( Xd_0__inst_mult_9_106  ) + ( Xd_0__inst_mult_9_105  ))
// Xd_0__inst_mult_9_109  = CARRY(( (din_a[66] & din_b[64]) ) + ( Xd_0__inst_mult_9_106  ) + ( Xd_0__inst_mult_9_105  ))
// Xd_0__inst_mult_9_110  = SHARE((din_a[66] & din_b[65]))

	.dataa(!din_a[66]),
	.datab(!din_b[64]),
	.datac(!din_b[65]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_105 ),
	.sharein(Xd_0__inst_mult_9_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_108 ),
	.cout(Xd_0__inst_mult_9_109 ),
	.shareout(Xd_0__inst_mult_9_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_35 (
// Equation(s):
// Xd_0__inst_mult_9_112  = SUM(( (din_a[63] & din_b[67]) ) + ( Xd_0__inst_mult_9_158  ) + ( Xd_0__inst_mult_9_157  ))
// Xd_0__inst_mult_9_113  = CARRY(( (din_a[63] & din_b[67]) ) + ( Xd_0__inst_mult_9_158  ) + ( Xd_0__inst_mult_9_157  ))
// Xd_0__inst_mult_9_114  = SHARE((din_a[65] & din_b[66]))

	.dataa(!din_a[63]),
	.datab(!din_b[67]),
	.datac(!din_a[65]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_157 ),
	.sharein(Xd_0__inst_mult_9_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_112 ),
	.cout(Xd_0__inst_mult_9_113 ),
	.shareout(Xd_0__inst_mult_9_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_34 (
// Equation(s):
// Xd_0__inst_mult_6_108  = SUM(( (din_a[45] & din_b[43]) ) + ( Xd_0__inst_mult_6_106  ) + ( Xd_0__inst_mult_6_105  ))
// Xd_0__inst_mult_6_109  = CARRY(( (din_a[45] & din_b[43]) ) + ( Xd_0__inst_mult_6_106  ) + ( Xd_0__inst_mult_6_105  ))
// Xd_0__inst_mult_6_110  = SHARE((din_a[45] & din_b[44]))

	.dataa(!din_a[45]),
	.datab(!din_b[43]),
	.datac(!din_b[44]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_105 ),
	.sharein(Xd_0__inst_mult_6_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_108 ),
	.cout(Xd_0__inst_mult_6_109 ),
	.shareout(Xd_0__inst_mult_6_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_35 (
// Equation(s):
// Xd_0__inst_mult_6_112  = SUM(( (din_a[42] & din_b[46]) ) + ( Xd_0__inst_mult_6_158  ) + ( Xd_0__inst_mult_6_157  ))
// Xd_0__inst_mult_6_113  = CARRY(( (din_a[42] & din_b[46]) ) + ( Xd_0__inst_mult_6_158  ) + ( Xd_0__inst_mult_6_157  ))
// Xd_0__inst_mult_6_114  = SHARE((din_a[44] & din_b[45]))

	.dataa(!din_a[42]),
	.datab(!din_b[46]),
	.datac(!din_a[44]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_157 ),
	.sharein(Xd_0__inst_mult_6_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_112 ),
	.cout(Xd_0__inst_mult_6_113 ),
	.shareout(Xd_0__inst_mult_6_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_34 (
// Equation(s):
// Xd_0__inst_mult_7_108  = SUM(( (din_a[52] & din_b[50]) ) + ( Xd_0__inst_mult_7_106  ) + ( Xd_0__inst_mult_7_105  ))
// Xd_0__inst_mult_7_109  = CARRY(( (din_a[52] & din_b[50]) ) + ( Xd_0__inst_mult_7_106  ) + ( Xd_0__inst_mult_7_105  ))
// Xd_0__inst_mult_7_110  = SHARE((din_a[52] & din_b[51]))

	.dataa(!din_a[52]),
	.datab(!din_b[50]),
	.datac(!din_b[51]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_105 ),
	.sharein(Xd_0__inst_mult_7_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_108 ),
	.cout(Xd_0__inst_mult_7_109 ),
	.shareout(Xd_0__inst_mult_7_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_35 (
// Equation(s):
// Xd_0__inst_mult_7_112  = SUM(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_7_158  ) + ( Xd_0__inst_mult_7_157  ))
// Xd_0__inst_mult_7_113  = CARRY(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_7_158  ) + ( Xd_0__inst_mult_7_157  ))
// Xd_0__inst_mult_7_114  = SHARE((din_a[51] & din_b[52]))

	.dataa(!din_a[49]),
	.datab(!din_b[53]),
	.datac(!din_a[51]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_157 ),
	.sharein(Xd_0__inst_mult_7_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_112 ),
	.cout(Xd_0__inst_mult_7_113 ),
	.shareout(Xd_0__inst_mult_7_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_34 (
// Equation(s):
// Xd_0__inst_mult_4_108  = SUM(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_4_106  ) + ( Xd_0__inst_mult_4_105  ))
// Xd_0__inst_mult_4_109  = CARRY(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_4_106  ) + ( Xd_0__inst_mult_4_105  ))
// Xd_0__inst_mult_4_110  = SHARE((din_a[31] & din_b[30]))

	.dataa(!din_a[31]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_105 ),
	.sharein(Xd_0__inst_mult_4_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_108 ),
	.cout(Xd_0__inst_mult_4_109 ),
	.shareout(Xd_0__inst_mult_4_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_35 (
// Equation(s):
// Xd_0__inst_mult_4_112  = SUM(( (din_a[28] & din_b[32]) ) + ( Xd_0__inst_mult_4_158  ) + ( Xd_0__inst_mult_4_157  ))
// Xd_0__inst_mult_4_113  = CARRY(( (din_a[28] & din_b[32]) ) + ( Xd_0__inst_mult_4_158  ) + ( Xd_0__inst_mult_4_157  ))
// Xd_0__inst_mult_4_114  = SHARE((din_a[30] & din_b[31]))

	.dataa(!din_a[28]),
	.datab(!din_b[32]),
	.datac(!din_a[30]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_157 ),
	.sharein(Xd_0__inst_mult_4_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_112 ),
	.cout(Xd_0__inst_mult_4_113 ),
	.shareout(Xd_0__inst_mult_4_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_34 (
// Equation(s):
// Xd_0__inst_mult_5_108  = SUM(( (din_a[38] & din_b[36]) ) + ( Xd_0__inst_mult_5_106  ) + ( Xd_0__inst_mult_5_105  ))
// Xd_0__inst_mult_5_109  = CARRY(( (din_a[38] & din_b[36]) ) + ( Xd_0__inst_mult_5_106  ) + ( Xd_0__inst_mult_5_105  ))
// Xd_0__inst_mult_5_110  = SHARE((din_a[38] & din_b[37]))

	.dataa(!din_a[38]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_105 ),
	.sharein(Xd_0__inst_mult_5_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_108 ),
	.cout(Xd_0__inst_mult_5_109 ),
	.shareout(Xd_0__inst_mult_5_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_35 (
// Equation(s):
// Xd_0__inst_mult_5_112  = SUM(( (din_a[35] & din_b[39]) ) + ( Xd_0__inst_mult_5_158  ) + ( Xd_0__inst_mult_5_157  ))
// Xd_0__inst_mult_5_113  = CARRY(( (din_a[35] & din_b[39]) ) + ( Xd_0__inst_mult_5_158  ) + ( Xd_0__inst_mult_5_157  ))
// Xd_0__inst_mult_5_114  = SHARE((din_a[37] & din_b[38]))

	.dataa(!din_a[35]),
	.datab(!din_b[39]),
	.datac(!din_a[37]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_157 ),
	.sharein(Xd_0__inst_mult_5_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_112 ),
	.cout(Xd_0__inst_mult_5_113 ),
	.shareout(Xd_0__inst_mult_5_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_34 (
// Equation(s):
// Xd_0__inst_mult_2_108  = SUM(( (din_a[17] & din_b[15]) ) + ( Xd_0__inst_mult_2_106  ) + ( Xd_0__inst_mult_2_105  ))
// Xd_0__inst_mult_2_109  = CARRY(( (din_a[17] & din_b[15]) ) + ( Xd_0__inst_mult_2_106  ) + ( Xd_0__inst_mult_2_105  ))
// Xd_0__inst_mult_2_110  = SHARE((din_a[17] & din_b[16]))

	.dataa(!din_a[17]),
	.datab(!din_b[15]),
	.datac(!din_b[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_105 ),
	.sharein(Xd_0__inst_mult_2_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_108 ),
	.cout(Xd_0__inst_mult_2_109 ),
	.shareout(Xd_0__inst_mult_2_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_35 (
// Equation(s):
// Xd_0__inst_mult_2_112  = SUM(( (din_a[14] & din_b[18]) ) + ( Xd_0__inst_mult_2_158  ) + ( Xd_0__inst_mult_2_157  ))
// Xd_0__inst_mult_2_113  = CARRY(( (din_a[14] & din_b[18]) ) + ( Xd_0__inst_mult_2_158  ) + ( Xd_0__inst_mult_2_157  ))
// Xd_0__inst_mult_2_114  = SHARE((din_a[16] & din_b[17]))

	.dataa(!din_a[14]),
	.datab(!din_b[18]),
	.datac(!din_a[16]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_157 ),
	.sharein(Xd_0__inst_mult_2_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_112 ),
	.cout(Xd_0__inst_mult_2_113 ),
	.shareout(Xd_0__inst_mult_2_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_34 (
// Equation(s):
// Xd_0__inst_mult_3_108  = SUM(( (din_a[24] & din_b[22]) ) + ( Xd_0__inst_mult_3_106  ) + ( Xd_0__inst_mult_3_105  ))
// Xd_0__inst_mult_3_109  = CARRY(( (din_a[24] & din_b[22]) ) + ( Xd_0__inst_mult_3_106  ) + ( Xd_0__inst_mult_3_105  ))
// Xd_0__inst_mult_3_110  = SHARE((din_a[24] & din_b[23]))

	.dataa(!din_a[24]),
	.datab(!din_b[22]),
	.datac(!din_b[23]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_105 ),
	.sharein(Xd_0__inst_mult_3_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_108 ),
	.cout(Xd_0__inst_mult_3_109 ),
	.shareout(Xd_0__inst_mult_3_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_35 (
// Equation(s):
// Xd_0__inst_mult_3_112  = SUM(( (din_a[21] & din_b[25]) ) + ( Xd_0__inst_mult_3_158  ) + ( Xd_0__inst_mult_3_157  ))
// Xd_0__inst_mult_3_113  = CARRY(( (din_a[21] & din_b[25]) ) + ( Xd_0__inst_mult_3_158  ) + ( Xd_0__inst_mult_3_157  ))
// Xd_0__inst_mult_3_114  = SHARE((din_a[23] & din_b[24]))

	.dataa(!din_a[21]),
	.datab(!din_b[25]),
	.datac(!din_a[23]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_157 ),
	.sharein(Xd_0__inst_mult_3_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_112 ),
	.cout(Xd_0__inst_mult_3_113 ),
	.shareout(Xd_0__inst_mult_3_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_34 (
// Equation(s):
// Xd_0__inst_mult_0_108  = SUM(( (din_a[3] & din_b[1]) ) + ( Xd_0__inst_mult_0_106  ) + ( Xd_0__inst_mult_0_105  ))
// Xd_0__inst_mult_0_109  = CARRY(( (din_a[3] & din_b[1]) ) + ( Xd_0__inst_mult_0_106  ) + ( Xd_0__inst_mult_0_105  ))
// Xd_0__inst_mult_0_110  = SHARE((din_a[3] & din_b[2]))

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(!din_b[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_105 ),
	.sharein(Xd_0__inst_mult_0_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_108 ),
	.cout(Xd_0__inst_mult_0_109 ),
	.shareout(Xd_0__inst_mult_0_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_35 (
// Equation(s):
// Xd_0__inst_mult_0_112  = SUM(( (din_a[0] & din_b[4]) ) + ( Xd_0__inst_mult_0_158  ) + ( Xd_0__inst_mult_0_157  ))
// Xd_0__inst_mult_0_113  = CARRY(( (din_a[0] & din_b[4]) ) + ( Xd_0__inst_mult_0_158  ) + ( Xd_0__inst_mult_0_157  ))
// Xd_0__inst_mult_0_114  = SHARE((din_a[2] & din_b[3]))

	.dataa(!din_a[0]),
	.datab(!din_b[4]),
	.datac(!din_a[2]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_157 ),
	.sharein(Xd_0__inst_mult_0_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_112 ),
	.cout(Xd_0__inst_mult_0_113 ),
	.shareout(Xd_0__inst_mult_0_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_34 (
// Equation(s):
// Xd_0__inst_mult_1_108  = SUM(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_106  ) + ( Xd_0__inst_mult_1_105  ))
// Xd_0__inst_mult_1_109  = CARRY(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_106  ) + ( Xd_0__inst_mult_1_105  ))
// Xd_0__inst_mult_1_110  = SHARE((din_a[10] & din_b[9]))

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(!din_b[9]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_105 ),
	.sharein(Xd_0__inst_mult_1_106 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_108 ),
	.cout(Xd_0__inst_mult_1_109 ),
	.shareout(Xd_0__inst_mult_1_110 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_35 (
// Equation(s):
// Xd_0__inst_mult_1_112  = SUM(( (din_a[7] & din_b[11]) ) + ( Xd_0__inst_mult_1_158  ) + ( Xd_0__inst_mult_1_157  ))
// Xd_0__inst_mult_1_113  = CARRY(( (din_a[7] & din_b[11]) ) + ( Xd_0__inst_mult_1_158  ) + ( Xd_0__inst_mult_1_157  ))
// Xd_0__inst_mult_1_114  = SHARE((din_a[9] & din_b[10]))

	.dataa(!din_a[7]),
	.datab(!din_b[11]),
	.datac(!din_a[9]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_157 ),
	.sharein(Xd_0__inst_mult_1_158 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_112 ),
	.cout(Xd_0__inst_mult_1_113 ),
	.shareout(Xd_0__inst_mult_1_114 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_36 (
// Equation(s):
// Xd_0__inst_mult_28_116  = SUM(( (!din_a[201] & (((din_a[200] & din_b[197])))) # (din_a[201] & (!din_b[196] $ (((!din_a[200]) # (!din_b[197]))))) ) + ( Xd_0__inst_mult_28_110  ) + ( Xd_0__inst_mult_28_109  ))
// Xd_0__inst_mult_28_117  = CARRY(( (!din_a[201] & (((din_a[200] & din_b[197])))) # (din_a[201] & (!din_b[196] $ (((!din_a[200]) # (!din_b[197]))))) ) + ( Xd_0__inst_mult_28_110  ) + ( Xd_0__inst_mult_28_109  ))
// Xd_0__inst_mult_28_118  = SHARE((din_a[201] & (din_b[196] & (din_a[200] & din_b[197]))))

	.dataa(!din_a[201]),
	.datab(!din_b[196]),
	.datac(!din_a[200]),
	.datad(!din_b[197]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_109 ),
	.sharein(Xd_0__inst_mult_28_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_116 ),
	.cout(Xd_0__inst_mult_28_117 ),
	.shareout(Xd_0__inst_mult_28_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_37 (
// Equation(s):
// Xd_0__inst_mult_28_120  = SUM(( (!din_a[197] & (((din_a[196] & din_b[201])))) # (din_a[197] & (!din_b[200] $ (((!din_a[196]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_114  ) + ( Xd_0__inst_mult_28_113  ))
// Xd_0__inst_mult_28_121  = CARRY(( (!din_a[197] & (((din_a[196] & din_b[201])))) # (din_a[197] & (!din_b[200] $ (((!din_a[196]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_114  ) + ( Xd_0__inst_mult_28_113  ))
// Xd_0__inst_mult_28_122  = SHARE((din_a[197] & (din_b[200] & (din_a[196] & din_b[201]))))

	.dataa(!din_a[197]),
	.datab(!din_b[200]),
	.datac(!din_a[196]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_113 ),
	.sharein(Xd_0__inst_mult_28_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_120 ),
	.cout(Xd_0__inst_mult_28_121 ),
	.shareout(Xd_0__inst_mult_28_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_36 (
// Equation(s):
// Xd_0__inst_mult_29_116  = SUM(( (!din_a[208] & (((din_a[207] & din_b[204])))) # (din_a[208] & (!din_b[203] $ (((!din_a[207]) # (!din_b[204]))))) ) + ( Xd_0__inst_mult_29_110  ) + ( Xd_0__inst_mult_29_109  ))
// Xd_0__inst_mult_29_117  = CARRY(( (!din_a[208] & (((din_a[207] & din_b[204])))) # (din_a[208] & (!din_b[203] $ (((!din_a[207]) # (!din_b[204]))))) ) + ( Xd_0__inst_mult_29_110  ) + ( Xd_0__inst_mult_29_109  ))
// Xd_0__inst_mult_29_118  = SHARE((din_a[208] & (din_b[203] & (din_a[207] & din_b[204]))))

	.dataa(!din_a[208]),
	.datab(!din_b[203]),
	.datac(!din_a[207]),
	.datad(!din_b[204]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_109 ),
	.sharein(Xd_0__inst_mult_29_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_116 ),
	.cout(Xd_0__inst_mult_29_117 ),
	.shareout(Xd_0__inst_mult_29_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_37 (
// Equation(s):
// Xd_0__inst_mult_29_120  = SUM(( (!din_a[204] & (((din_a[203] & din_b[208])))) # (din_a[204] & (!din_b[207] $ (((!din_a[203]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_114  ) + ( Xd_0__inst_mult_29_113  ))
// Xd_0__inst_mult_29_121  = CARRY(( (!din_a[204] & (((din_a[203] & din_b[208])))) # (din_a[204] & (!din_b[207] $ (((!din_a[203]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_114  ) + ( Xd_0__inst_mult_29_113  ))
// Xd_0__inst_mult_29_122  = SHARE((din_a[204] & (din_b[207] & (din_a[203] & din_b[208]))))

	.dataa(!din_a[204]),
	.datab(!din_b[207]),
	.datac(!din_a[203]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_113 ),
	.sharein(Xd_0__inst_mult_29_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_120 ),
	.cout(Xd_0__inst_mult_29_121 ),
	.shareout(Xd_0__inst_mult_29_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_36 (
// Equation(s):
// Xd_0__inst_mult_26_116  = SUM(( (!din_a[187] & (((din_a[186] & din_b[183])))) # (din_a[187] & (!din_b[182] $ (((!din_a[186]) # (!din_b[183]))))) ) + ( Xd_0__inst_mult_26_110  ) + ( Xd_0__inst_mult_26_109  ))
// Xd_0__inst_mult_26_117  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[183])))) # (din_a[187] & (!din_b[182] $ (((!din_a[186]) # (!din_b[183]))))) ) + ( Xd_0__inst_mult_26_110  ) + ( Xd_0__inst_mult_26_109  ))
// Xd_0__inst_mult_26_118  = SHARE((din_a[187] & (din_b[182] & (din_a[186] & din_b[183]))))

	.dataa(!din_a[187]),
	.datab(!din_b[182]),
	.datac(!din_a[186]),
	.datad(!din_b[183]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_109 ),
	.sharein(Xd_0__inst_mult_26_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_116 ),
	.cout(Xd_0__inst_mult_26_117 ),
	.shareout(Xd_0__inst_mult_26_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_37 (
// Equation(s):
// Xd_0__inst_mult_26_120  = SUM(( (!din_a[183] & (((din_a[182] & din_b[187])))) # (din_a[183] & (!din_b[186] $ (((!din_a[182]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_114  ) + ( Xd_0__inst_mult_26_113  ))
// Xd_0__inst_mult_26_121  = CARRY(( (!din_a[183] & (((din_a[182] & din_b[187])))) # (din_a[183] & (!din_b[186] $ (((!din_a[182]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_114  ) + ( Xd_0__inst_mult_26_113  ))
// Xd_0__inst_mult_26_122  = SHARE((din_a[183] & (din_b[186] & (din_a[182] & din_b[187]))))

	.dataa(!din_a[183]),
	.datab(!din_b[186]),
	.datac(!din_a[182]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_113 ),
	.sharein(Xd_0__inst_mult_26_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_120 ),
	.cout(Xd_0__inst_mult_26_121 ),
	.shareout(Xd_0__inst_mult_26_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_36 (
// Equation(s):
// Xd_0__inst_mult_27_116  = SUM(( (!din_a[194] & (((din_a[193] & din_b[190])))) # (din_a[194] & (!din_b[189] $ (((!din_a[193]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_27_110  ) + ( Xd_0__inst_mult_27_109  ))
// Xd_0__inst_mult_27_117  = CARRY(( (!din_a[194] & (((din_a[193] & din_b[190])))) # (din_a[194] & (!din_b[189] $ (((!din_a[193]) # (!din_b[190]))))) ) + ( Xd_0__inst_mult_27_110  ) + ( Xd_0__inst_mult_27_109  ))
// Xd_0__inst_mult_27_118  = SHARE((din_a[194] & (din_b[189] & (din_a[193] & din_b[190]))))

	.dataa(!din_a[194]),
	.datab(!din_b[189]),
	.datac(!din_a[193]),
	.datad(!din_b[190]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_109 ),
	.sharein(Xd_0__inst_mult_27_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_116 ),
	.cout(Xd_0__inst_mult_27_117 ),
	.shareout(Xd_0__inst_mult_27_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_37 (
// Equation(s):
// Xd_0__inst_mult_27_120  = SUM(( (!din_a[190] & (((din_a[189] & din_b[194])))) # (din_a[190] & (!din_b[193] $ (((!din_a[189]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_114  ) + ( Xd_0__inst_mult_27_113  ))
// Xd_0__inst_mult_27_121  = CARRY(( (!din_a[190] & (((din_a[189] & din_b[194])))) # (din_a[190] & (!din_b[193] $ (((!din_a[189]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_114  ) + ( Xd_0__inst_mult_27_113  ))
// Xd_0__inst_mult_27_122  = SHARE((din_a[190] & (din_b[193] & (din_a[189] & din_b[194]))))

	.dataa(!din_a[190]),
	.datab(!din_b[193]),
	.datac(!din_a[189]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_113 ),
	.sharein(Xd_0__inst_mult_27_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_120 ),
	.cout(Xd_0__inst_mult_27_121 ),
	.shareout(Xd_0__inst_mult_27_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_36 (
// Equation(s):
// Xd_0__inst_mult_24_116  = SUM(( (!din_a[173] & (((din_a[172] & din_b[169])))) # (din_a[173] & (!din_b[168] $ (((!din_a[172]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_24_110  ) + ( Xd_0__inst_mult_24_109  ))
// Xd_0__inst_mult_24_117  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[169])))) # (din_a[173] & (!din_b[168] $ (((!din_a[172]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_24_110  ) + ( Xd_0__inst_mult_24_109  ))
// Xd_0__inst_mult_24_118  = SHARE((din_a[173] & (din_b[168] & (din_a[172] & din_b[169]))))

	.dataa(!din_a[173]),
	.datab(!din_b[168]),
	.datac(!din_a[172]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_109 ),
	.sharein(Xd_0__inst_mult_24_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_116 ),
	.cout(Xd_0__inst_mult_24_117 ),
	.shareout(Xd_0__inst_mult_24_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_37 (
// Equation(s):
// Xd_0__inst_mult_24_120  = SUM(( (!din_a[169] & (((din_a[168] & din_b[173])))) # (din_a[169] & (!din_b[172] $ (((!din_a[168]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_114  ) + ( Xd_0__inst_mult_24_113  ))
// Xd_0__inst_mult_24_121  = CARRY(( (!din_a[169] & (((din_a[168] & din_b[173])))) # (din_a[169] & (!din_b[172] $ (((!din_a[168]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_114  ) + ( Xd_0__inst_mult_24_113  ))
// Xd_0__inst_mult_24_122  = SHARE((din_a[169] & (din_b[172] & (din_a[168] & din_b[173]))))

	.dataa(!din_a[169]),
	.datab(!din_b[172]),
	.datac(!din_a[168]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_113 ),
	.sharein(Xd_0__inst_mult_24_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_120 ),
	.cout(Xd_0__inst_mult_24_121 ),
	.shareout(Xd_0__inst_mult_24_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_37 (
// Equation(s):
// Xd_0__inst_mult_25_120  = SUM(( (!din_a[180] & (((din_a[179] & din_b[176])))) # (din_a[180] & (!din_b[175] $ (((!din_a[179]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_25_114  ) + ( Xd_0__inst_mult_25_113  ))
// Xd_0__inst_mult_25_121  = CARRY(( (!din_a[180] & (((din_a[179] & din_b[176])))) # (din_a[180] & (!din_b[175] $ (((!din_a[179]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_25_114  ) + ( Xd_0__inst_mult_25_113  ))
// Xd_0__inst_mult_25_122  = SHARE((din_a[180] & (din_b[175] & (din_a[179] & din_b[176]))))

	.dataa(!din_a[180]),
	.datab(!din_b[175]),
	.datac(!din_a[179]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_113 ),
	.sharein(Xd_0__inst_mult_25_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_120 ),
	.cout(Xd_0__inst_mult_25_121 ),
	.shareout(Xd_0__inst_mult_25_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_38 (
// Equation(s):
// Xd_0__inst_mult_25_124  = SUM(( (!din_a[176] & (((din_a[175] & din_b[180])))) # (din_a[176] & (!din_b[179] $ (((!din_a[175]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_118  ) + ( Xd_0__inst_mult_25_117  ))
// Xd_0__inst_mult_25_125  = CARRY(( (!din_a[176] & (((din_a[175] & din_b[180])))) # (din_a[176] & (!din_b[179] $ (((!din_a[175]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_118  ) + ( Xd_0__inst_mult_25_117  ))
// Xd_0__inst_mult_25_126  = SHARE((din_a[176] & (din_b[179] & (din_a[175] & din_b[180]))))

	.dataa(!din_a[176]),
	.datab(!din_b[179]),
	.datac(!din_a[175]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_117 ),
	.sharein(Xd_0__inst_mult_25_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_124 ),
	.cout(Xd_0__inst_mult_25_125 ),
	.shareout(Xd_0__inst_mult_25_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_37 (
// Equation(s):
// Xd_0__inst_mult_22_120  = SUM(( (!din_a[159] & (((din_a[158] & din_b[155])))) # (din_a[159] & (!din_b[154] $ (((!din_a[158]) # (!din_b[155]))))) ) + ( Xd_0__inst_mult_22_114  ) + ( Xd_0__inst_mult_22_113  ))
// Xd_0__inst_mult_22_121  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[155])))) # (din_a[159] & (!din_b[154] $ (((!din_a[158]) # (!din_b[155]))))) ) + ( Xd_0__inst_mult_22_114  ) + ( Xd_0__inst_mult_22_113  ))
// Xd_0__inst_mult_22_122  = SHARE((din_a[159] & (din_b[154] & (din_a[158] & din_b[155]))))

	.dataa(!din_a[159]),
	.datab(!din_b[154]),
	.datac(!din_a[158]),
	.datad(!din_b[155]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_113 ),
	.sharein(Xd_0__inst_mult_22_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_120 ),
	.cout(Xd_0__inst_mult_22_121 ),
	.shareout(Xd_0__inst_mult_22_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_38 (
// Equation(s):
// Xd_0__inst_mult_22_124  = SUM(( (!din_a[155] & (((din_a[154] & din_b[159])))) # (din_a[155] & (!din_b[158] $ (((!din_a[154]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_118  ) + ( Xd_0__inst_mult_22_117  ))
// Xd_0__inst_mult_22_125  = CARRY(( (!din_a[155] & (((din_a[154] & din_b[159])))) # (din_a[155] & (!din_b[158] $ (((!din_a[154]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_118  ) + ( Xd_0__inst_mult_22_117  ))
// Xd_0__inst_mult_22_126  = SHARE((din_a[155] & (din_b[158] & (din_a[154] & din_b[159]))))

	.dataa(!din_a[155]),
	.datab(!din_b[158]),
	.datac(!din_a[154]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_117 ),
	.sharein(Xd_0__inst_mult_22_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_124 ),
	.cout(Xd_0__inst_mult_22_125 ),
	.shareout(Xd_0__inst_mult_22_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_36 (
// Equation(s):
// Xd_0__inst_mult_23_116  = SUM(( (!din_a[166] & (((din_a[165] & din_b[162])))) # (din_a[166] & (!din_b[161] $ (((!din_a[165]) # (!din_b[162]))))) ) + ( Xd_0__inst_mult_23_110  ) + ( Xd_0__inst_mult_23_109  ))
// Xd_0__inst_mult_23_117  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[162])))) # (din_a[166] & (!din_b[161] $ (((!din_a[165]) # (!din_b[162]))))) ) + ( Xd_0__inst_mult_23_110  ) + ( Xd_0__inst_mult_23_109  ))
// Xd_0__inst_mult_23_118  = SHARE((din_a[166] & (din_b[161] & (din_a[165] & din_b[162]))))

	.dataa(!din_a[166]),
	.datab(!din_b[161]),
	.datac(!din_a[165]),
	.datad(!din_b[162]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_109 ),
	.sharein(Xd_0__inst_mult_23_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_116 ),
	.cout(Xd_0__inst_mult_23_117 ),
	.shareout(Xd_0__inst_mult_23_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_37 (
// Equation(s):
// Xd_0__inst_mult_23_120  = SUM(( (!din_a[162] & (((din_a[161] & din_b[166])))) # (din_a[162] & (!din_b[165] $ (((!din_a[161]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_114  ) + ( Xd_0__inst_mult_23_113  ))
// Xd_0__inst_mult_23_121  = CARRY(( (!din_a[162] & (((din_a[161] & din_b[166])))) # (din_a[162] & (!din_b[165] $ (((!din_a[161]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_114  ) + ( Xd_0__inst_mult_23_113  ))
// Xd_0__inst_mult_23_122  = SHARE((din_a[162] & (din_b[165] & (din_a[161] & din_b[166]))))

	.dataa(!din_a[162]),
	.datab(!din_b[165]),
	.datac(!din_a[161]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_113 ),
	.sharein(Xd_0__inst_mult_23_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_120 ),
	.cout(Xd_0__inst_mult_23_121 ),
	.shareout(Xd_0__inst_mult_23_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_36 (
// Equation(s):
// Xd_0__inst_mult_20_116  = SUM(( (!din_a[145] & (((din_a[144] & din_b[141])))) # (din_a[145] & (!din_b[140] $ (((!din_a[144]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_20_110  ) + ( Xd_0__inst_mult_20_109  ))
// Xd_0__inst_mult_20_117  = CARRY(( (!din_a[145] & (((din_a[144] & din_b[141])))) # (din_a[145] & (!din_b[140] $ (((!din_a[144]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_20_110  ) + ( Xd_0__inst_mult_20_109  ))
// Xd_0__inst_mult_20_118  = SHARE((din_a[145] & (din_b[140] & (din_a[144] & din_b[141]))))

	.dataa(!din_a[145]),
	.datab(!din_b[140]),
	.datac(!din_a[144]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_109 ),
	.sharein(Xd_0__inst_mult_20_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_116 ),
	.cout(Xd_0__inst_mult_20_117 ),
	.shareout(Xd_0__inst_mult_20_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_37 (
// Equation(s):
// Xd_0__inst_mult_20_120  = SUM(( (!din_a[141] & (((din_a[140] & din_b[145])))) # (din_a[141] & (!din_b[144] $ (((!din_a[140]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_114  ) + ( Xd_0__inst_mult_20_113  ))
// Xd_0__inst_mult_20_121  = CARRY(( (!din_a[141] & (((din_a[140] & din_b[145])))) # (din_a[141] & (!din_b[144] $ (((!din_a[140]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_114  ) + ( Xd_0__inst_mult_20_113  ))
// Xd_0__inst_mult_20_122  = SHARE((din_a[141] & (din_b[144] & (din_a[140] & din_b[145]))))

	.dataa(!din_a[141]),
	.datab(!din_b[144]),
	.datac(!din_a[140]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_113 ),
	.sharein(Xd_0__inst_mult_20_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_120 ),
	.cout(Xd_0__inst_mult_20_121 ),
	.shareout(Xd_0__inst_mult_20_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_36 (
// Equation(s):
// Xd_0__inst_mult_21_116  = SUM(( (!din_a[152] & (((din_a[151] & din_b[148])))) # (din_a[152] & (!din_b[147] $ (((!din_a[151]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_21_110  ) + ( Xd_0__inst_mult_21_109  ))
// Xd_0__inst_mult_21_117  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[148])))) # (din_a[152] & (!din_b[147] $ (((!din_a[151]) # (!din_b[148]))))) ) + ( Xd_0__inst_mult_21_110  ) + ( Xd_0__inst_mult_21_109  ))
// Xd_0__inst_mult_21_118  = SHARE((din_a[152] & (din_b[147] & (din_a[151] & din_b[148]))))

	.dataa(!din_a[152]),
	.datab(!din_b[147]),
	.datac(!din_a[151]),
	.datad(!din_b[148]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_109 ),
	.sharein(Xd_0__inst_mult_21_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_116 ),
	.cout(Xd_0__inst_mult_21_117 ),
	.shareout(Xd_0__inst_mult_21_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_37 (
// Equation(s):
// Xd_0__inst_mult_21_120  = SUM(( (!din_a[148] & (((din_a[147] & din_b[152])))) # (din_a[148] & (!din_b[151] $ (((!din_a[147]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_114  ) + ( Xd_0__inst_mult_21_113  ))
// Xd_0__inst_mult_21_121  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[152])))) # (din_a[148] & (!din_b[151] $ (((!din_a[147]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_114  ) + ( Xd_0__inst_mult_21_113  ))
// Xd_0__inst_mult_21_122  = SHARE((din_a[148] & (din_b[151] & (din_a[147] & din_b[152]))))

	.dataa(!din_a[148]),
	.datab(!din_b[151]),
	.datac(!din_a[147]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_113 ),
	.sharein(Xd_0__inst_mult_21_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_120 ),
	.cout(Xd_0__inst_mult_21_121 ),
	.shareout(Xd_0__inst_mult_21_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_36 (
// Equation(s):
// Xd_0__inst_mult_18_116  = SUM(( (!din_a[131] & (((din_a[130] & din_b[127])))) # (din_a[131] & (!din_b[126] $ (((!din_a[130]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_18_110  ) + ( Xd_0__inst_mult_18_109  ))
// Xd_0__inst_mult_18_117  = CARRY(( (!din_a[131] & (((din_a[130] & din_b[127])))) # (din_a[131] & (!din_b[126] $ (((!din_a[130]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_18_110  ) + ( Xd_0__inst_mult_18_109  ))
// Xd_0__inst_mult_18_118  = SHARE((din_a[131] & (din_b[126] & (din_a[130] & din_b[127]))))

	.dataa(!din_a[131]),
	.datab(!din_b[126]),
	.datac(!din_a[130]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_109 ),
	.sharein(Xd_0__inst_mult_18_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_116 ),
	.cout(Xd_0__inst_mult_18_117 ),
	.shareout(Xd_0__inst_mult_18_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_37 (
// Equation(s):
// Xd_0__inst_mult_18_120  = SUM(( (!din_a[127] & (((din_a[126] & din_b[131])))) # (din_a[127] & (!din_b[130] $ (((!din_a[126]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_114  ) + ( Xd_0__inst_mult_18_113  ))
// Xd_0__inst_mult_18_121  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[131])))) # (din_a[127] & (!din_b[130] $ (((!din_a[126]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_114  ) + ( Xd_0__inst_mult_18_113  ))
// Xd_0__inst_mult_18_122  = SHARE((din_a[127] & (din_b[130] & (din_a[126] & din_b[131]))))

	.dataa(!din_a[127]),
	.datab(!din_b[130]),
	.datac(!din_a[126]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_113 ),
	.sharein(Xd_0__inst_mult_18_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_120 ),
	.cout(Xd_0__inst_mult_18_121 ),
	.shareout(Xd_0__inst_mult_18_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_36 (
// Equation(s):
// Xd_0__inst_mult_19_116  = SUM(( (!din_a[138] & (((din_a[137] & din_b[134])))) # (din_a[138] & (!din_b[133] $ (((!din_a[137]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_19_110  ) + ( Xd_0__inst_mult_19_109  ))
// Xd_0__inst_mult_19_117  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[134])))) # (din_a[138] & (!din_b[133] $ (((!din_a[137]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_19_110  ) + ( Xd_0__inst_mult_19_109  ))
// Xd_0__inst_mult_19_118  = SHARE((din_a[138] & (din_b[133] & (din_a[137] & din_b[134]))))

	.dataa(!din_a[138]),
	.datab(!din_b[133]),
	.datac(!din_a[137]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_109 ),
	.sharein(Xd_0__inst_mult_19_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_116 ),
	.cout(Xd_0__inst_mult_19_117 ),
	.shareout(Xd_0__inst_mult_19_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_37 (
// Equation(s):
// Xd_0__inst_mult_19_120  = SUM(( (!din_a[134] & (((din_a[133] & din_b[138])))) # (din_a[134] & (!din_b[137] $ (((!din_a[133]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_114  ) + ( Xd_0__inst_mult_19_113  ))
// Xd_0__inst_mult_19_121  = CARRY(( (!din_a[134] & (((din_a[133] & din_b[138])))) # (din_a[134] & (!din_b[137] $ (((!din_a[133]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_114  ) + ( Xd_0__inst_mult_19_113  ))
// Xd_0__inst_mult_19_122  = SHARE((din_a[134] & (din_b[137] & (din_a[133] & din_b[138]))))

	.dataa(!din_a[134]),
	.datab(!din_b[137]),
	.datac(!din_a[133]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_113 ),
	.sharein(Xd_0__inst_mult_19_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_120 ),
	.cout(Xd_0__inst_mult_19_121 ),
	.shareout(Xd_0__inst_mult_19_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_36 (
// Equation(s):
// Xd_0__inst_mult_16_116  = SUM(( (!din_a[117] & (((din_a[116] & din_b[113])))) # (din_a[117] & (!din_b[112] $ (((!din_a[116]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_16_110  ) + ( Xd_0__inst_mult_16_109  ))
// Xd_0__inst_mult_16_117  = CARRY(( (!din_a[117] & (((din_a[116] & din_b[113])))) # (din_a[117] & (!din_b[112] $ (((!din_a[116]) # (!din_b[113]))))) ) + ( Xd_0__inst_mult_16_110  ) + ( Xd_0__inst_mult_16_109  ))
// Xd_0__inst_mult_16_118  = SHARE((din_a[117] & (din_b[112] & (din_a[116] & din_b[113]))))

	.dataa(!din_a[117]),
	.datab(!din_b[112]),
	.datac(!din_a[116]),
	.datad(!din_b[113]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_109 ),
	.sharein(Xd_0__inst_mult_16_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_116 ),
	.cout(Xd_0__inst_mult_16_117 ),
	.shareout(Xd_0__inst_mult_16_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_37 (
// Equation(s):
// Xd_0__inst_mult_16_120  = SUM(( (!din_a[113] & (((din_a[112] & din_b[117])))) # (din_a[113] & (!din_b[116] $ (((!din_a[112]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_114  ) + ( Xd_0__inst_mult_16_113  ))
// Xd_0__inst_mult_16_121  = CARRY(( (!din_a[113] & (((din_a[112] & din_b[117])))) # (din_a[113] & (!din_b[116] $ (((!din_a[112]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_114  ) + ( Xd_0__inst_mult_16_113  ))
// Xd_0__inst_mult_16_122  = SHARE((din_a[113] & (din_b[116] & (din_a[112] & din_b[117]))))

	.dataa(!din_a[113]),
	.datab(!din_b[116]),
	.datac(!din_a[112]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_113 ),
	.sharein(Xd_0__inst_mult_16_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_120 ),
	.cout(Xd_0__inst_mult_16_121 ),
	.shareout(Xd_0__inst_mult_16_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_36 (
// Equation(s):
// Xd_0__inst_mult_17_116  = SUM(( (!din_a[124] & (((din_a[123] & din_b[120])))) # (din_a[124] & (!din_b[119] $ (((!din_a[123]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_17_110  ) + ( Xd_0__inst_mult_17_109  ))
// Xd_0__inst_mult_17_117  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[120])))) # (din_a[124] & (!din_b[119] $ (((!din_a[123]) # (!din_b[120]))))) ) + ( Xd_0__inst_mult_17_110  ) + ( Xd_0__inst_mult_17_109  ))
// Xd_0__inst_mult_17_118  = SHARE((din_a[124] & (din_b[119] & (din_a[123] & din_b[120]))))

	.dataa(!din_a[124]),
	.datab(!din_b[119]),
	.datac(!din_a[123]),
	.datad(!din_b[120]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_109 ),
	.sharein(Xd_0__inst_mult_17_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_116 ),
	.cout(Xd_0__inst_mult_17_117 ),
	.shareout(Xd_0__inst_mult_17_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_37 (
// Equation(s):
// Xd_0__inst_mult_17_120  = SUM(( (!din_a[120] & (((din_a[119] & din_b[124])))) # (din_a[120] & (!din_b[123] $ (((!din_a[119]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_114  ) + ( Xd_0__inst_mult_17_113  ))
// Xd_0__inst_mult_17_121  = CARRY(( (!din_a[120] & (((din_a[119] & din_b[124])))) # (din_a[120] & (!din_b[123] $ (((!din_a[119]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_114  ) + ( Xd_0__inst_mult_17_113  ))
// Xd_0__inst_mult_17_122  = SHARE((din_a[120] & (din_b[123] & (din_a[119] & din_b[124]))))

	.dataa(!din_a[120]),
	.datab(!din_b[123]),
	.datac(!din_a[119]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_113 ),
	.sharein(Xd_0__inst_mult_17_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_120 ),
	.cout(Xd_0__inst_mult_17_121 ),
	.shareout(Xd_0__inst_mult_17_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_36 (
// Equation(s):
// Xd_0__inst_mult_14_116  = SUM(( (!din_a[103] & (((din_a[102] & din_b[99])))) # (din_a[103] & (!din_b[98] $ (((!din_a[102]) # (!din_b[99]))))) ) + ( Xd_0__inst_mult_14_110  ) + ( Xd_0__inst_mult_14_109  ))
// Xd_0__inst_mult_14_117  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[99])))) # (din_a[103] & (!din_b[98] $ (((!din_a[102]) # (!din_b[99]))))) ) + ( Xd_0__inst_mult_14_110  ) + ( Xd_0__inst_mult_14_109  ))
// Xd_0__inst_mult_14_118  = SHARE((din_a[103] & (din_b[98] & (din_a[102] & din_b[99]))))

	.dataa(!din_a[103]),
	.datab(!din_b[98]),
	.datac(!din_a[102]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_109 ),
	.sharein(Xd_0__inst_mult_14_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_116 ),
	.cout(Xd_0__inst_mult_14_117 ),
	.shareout(Xd_0__inst_mult_14_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_37 (
// Equation(s):
// Xd_0__inst_mult_14_120  = SUM(( (!din_a[99] & (((din_a[98] & din_b[103])))) # (din_a[99] & (!din_b[102] $ (((!din_a[98]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_114  ) + ( Xd_0__inst_mult_14_113  ))
// Xd_0__inst_mult_14_121  = CARRY(( (!din_a[99] & (((din_a[98] & din_b[103])))) # (din_a[99] & (!din_b[102] $ (((!din_a[98]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_114  ) + ( Xd_0__inst_mult_14_113  ))
// Xd_0__inst_mult_14_122  = SHARE((din_a[99] & (din_b[102] & (din_a[98] & din_b[103]))))

	.dataa(!din_a[99]),
	.datab(!din_b[102]),
	.datac(!din_a[98]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_113 ),
	.sharein(Xd_0__inst_mult_14_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_120 ),
	.cout(Xd_0__inst_mult_14_121 ),
	.shareout(Xd_0__inst_mult_14_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_36 (
// Equation(s):
// Xd_0__inst_mult_15_116  = SUM(( (!din_a[110] & (((din_a[109] & din_b[106])))) # (din_a[110] & (!din_b[105] $ (((!din_a[109]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_15_110  ) + ( Xd_0__inst_mult_15_109  ))
// Xd_0__inst_mult_15_117  = CARRY(( (!din_a[110] & (((din_a[109] & din_b[106])))) # (din_a[110] & (!din_b[105] $ (((!din_a[109]) # (!din_b[106]))))) ) + ( Xd_0__inst_mult_15_110  ) + ( Xd_0__inst_mult_15_109  ))
// Xd_0__inst_mult_15_118  = SHARE((din_a[110] & (din_b[105] & (din_a[109] & din_b[106]))))

	.dataa(!din_a[110]),
	.datab(!din_b[105]),
	.datac(!din_a[109]),
	.datad(!din_b[106]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_109 ),
	.sharein(Xd_0__inst_mult_15_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_116 ),
	.cout(Xd_0__inst_mult_15_117 ),
	.shareout(Xd_0__inst_mult_15_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_37 (
// Equation(s):
// Xd_0__inst_mult_15_120  = SUM(( (!din_a[106] & (((din_a[105] & din_b[110])))) # (din_a[106] & (!din_b[109] $ (((!din_a[105]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_114  ) + ( Xd_0__inst_mult_15_113  ))
// Xd_0__inst_mult_15_121  = CARRY(( (!din_a[106] & (((din_a[105] & din_b[110])))) # (din_a[106] & (!din_b[109] $ (((!din_a[105]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_114  ) + ( Xd_0__inst_mult_15_113  ))
// Xd_0__inst_mult_15_122  = SHARE((din_a[106] & (din_b[109] & (din_a[105] & din_b[110]))))

	.dataa(!din_a[106]),
	.datab(!din_b[109]),
	.datac(!din_a[105]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_113 ),
	.sharein(Xd_0__inst_mult_15_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_120 ),
	.cout(Xd_0__inst_mult_15_121 ),
	.shareout(Xd_0__inst_mult_15_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_36 (
// Equation(s):
// Xd_0__inst_mult_12_116  = SUM(( (!din_a[89] & (((din_a[88] & din_b[85])))) # (din_a[89] & (!din_b[84] $ (((!din_a[88]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_12_110  ) + ( Xd_0__inst_mult_12_109  ))
// Xd_0__inst_mult_12_117  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[85])))) # (din_a[89] & (!din_b[84] $ (((!din_a[88]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_12_110  ) + ( Xd_0__inst_mult_12_109  ))
// Xd_0__inst_mult_12_118  = SHARE((din_a[89] & (din_b[84] & (din_a[88] & din_b[85]))))

	.dataa(!din_a[89]),
	.datab(!din_b[84]),
	.datac(!din_a[88]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_109 ),
	.sharein(Xd_0__inst_mult_12_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_116 ),
	.cout(Xd_0__inst_mult_12_117 ),
	.shareout(Xd_0__inst_mult_12_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_37 (
// Equation(s):
// Xd_0__inst_mult_12_120  = SUM(( (!din_a[85] & (((din_a[84] & din_b[89])))) # (din_a[85] & (!din_b[88] $ (((!din_a[84]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_114  ) + ( Xd_0__inst_mult_12_113  ))
// Xd_0__inst_mult_12_121  = CARRY(( (!din_a[85] & (((din_a[84] & din_b[89])))) # (din_a[85] & (!din_b[88] $ (((!din_a[84]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_114  ) + ( Xd_0__inst_mult_12_113  ))
// Xd_0__inst_mult_12_122  = SHARE((din_a[85] & (din_b[88] & (din_a[84] & din_b[89]))))

	.dataa(!din_a[85]),
	.datab(!din_b[88]),
	.datac(!din_a[84]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_113 ),
	.sharein(Xd_0__inst_mult_12_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_120 ),
	.cout(Xd_0__inst_mult_12_121 ),
	.shareout(Xd_0__inst_mult_12_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_36 (
// Equation(s):
// Xd_0__inst_mult_13_116  = SUM(( (!din_a[96] & (((din_a[95] & din_b[92])))) # (din_a[96] & (!din_b[91] $ (((!din_a[95]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_13_110  ) + ( Xd_0__inst_mult_13_109  ))
// Xd_0__inst_mult_13_117  = CARRY(( (!din_a[96] & (((din_a[95] & din_b[92])))) # (din_a[96] & (!din_b[91] $ (((!din_a[95]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_13_110  ) + ( Xd_0__inst_mult_13_109  ))
// Xd_0__inst_mult_13_118  = SHARE((din_a[96] & (din_b[91] & (din_a[95] & din_b[92]))))

	.dataa(!din_a[96]),
	.datab(!din_b[91]),
	.datac(!din_a[95]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_109 ),
	.sharein(Xd_0__inst_mult_13_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_116 ),
	.cout(Xd_0__inst_mult_13_117 ),
	.shareout(Xd_0__inst_mult_13_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_37 (
// Equation(s):
// Xd_0__inst_mult_13_120  = SUM(( (!din_a[92] & (((din_a[91] & din_b[96])))) # (din_a[92] & (!din_b[95] $ (((!din_a[91]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_114  ) + ( Xd_0__inst_mult_13_113  ))
// Xd_0__inst_mult_13_121  = CARRY(( (!din_a[92] & (((din_a[91] & din_b[96])))) # (din_a[92] & (!din_b[95] $ (((!din_a[91]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_114  ) + ( Xd_0__inst_mult_13_113  ))
// Xd_0__inst_mult_13_122  = SHARE((din_a[92] & (din_b[95] & (din_a[91] & din_b[96]))))

	.dataa(!din_a[92]),
	.datab(!din_b[95]),
	.datac(!din_a[91]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_113 ),
	.sharein(Xd_0__inst_mult_13_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_120 ),
	.cout(Xd_0__inst_mult_13_121 ),
	.shareout(Xd_0__inst_mult_13_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_36 (
// Equation(s):
// Xd_0__inst_mult_10_116  = SUM(( (!din_a[75] & (((din_a[74] & din_b[71])))) # (din_a[75] & (!din_b[70] $ (((!din_a[74]) # (!din_b[71]))))) ) + ( Xd_0__inst_mult_10_110  ) + ( Xd_0__inst_mult_10_109  ))
// Xd_0__inst_mult_10_117  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[71])))) # (din_a[75] & (!din_b[70] $ (((!din_a[74]) # (!din_b[71]))))) ) + ( Xd_0__inst_mult_10_110  ) + ( Xd_0__inst_mult_10_109  ))
// Xd_0__inst_mult_10_118  = SHARE((din_a[75] & (din_b[70] & (din_a[74] & din_b[71]))))

	.dataa(!din_a[75]),
	.datab(!din_b[70]),
	.datac(!din_a[74]),
	.datad(!din_b[71]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_109 ),
	.sharein(Xd_0__inst_mult_10_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_116 ),
	.cout(Xd_0__inst_mult_10_117 ),
	.shareout(Xd_0__inst_mult_10_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_37 (
// Equation(s):
// Xd_0__inst_mult_10_120  = SUM(( (!din_a[71] & (((din_a[70] & din_b[75])))) # (din_a[71] & (!din_b[74] $ (((!din_a[70]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_114  ) + ( Xd_0__inst_mult_10_113  ))
// Xd_0__inst_mult_10_121  = CARRY(( (!din_a[71] & (((din_a[70] & din_b[75])))) # (din_a[71] & (!din_b[74] $ (((!din_a[70]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_114  ) + ( Xd_0__inst_mult_10_113  ))
// Xd_0__inst_mult_10_122  = SHARE((din_a[71] & (din_b[74] & (din_a[70] & din_b[75]))))

	.dataa(!din_a[71]),
	.datab(!din_b[74]),
	.datac(!din_a[70]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_113 ),
	.sharein(Xd_0__inst_mult_10_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_120 ),
	.cout(Xd_0__inst_mult_10_121 ),
	.shareout(Xd_0__inst_mult_10_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_36 (
// Equation(s):
// Xd_0__inst_mult_11_116  = SUM(( (!din_a[82] & (((din_a[81] & din_b[78])))) # (din_a[82] & (!din_b[77] $ (((!din_a[81]) # (!din_b[78]))))) ) + ( Xd_0__inst_mult_11_110  ) + ( Xd_0__inst_mult_11_109  ))
// Xd_0__inst_mult_11_117  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[78])))) # (din_a[82] & (!din_b[77] $ (((!din_a[81]) # (!din_b[78]))))) ) + ( Xd_0__inst_mult_11_110  ) + ( Xd_0__inst_mult_11_109  ))
// Xd_0__inst_mult_11_118  = SHARE((din_a[82] & (din_b[77] & (din_a[81] & din_b[78]))))

	.dataa(!din_a[82]),
	.datab(!din_b[77]),
	.datac(!din_a[81]),
	.datad(!din_b[78]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_109 ),
	.sharein(Xd_0__inst_mult_11_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_116 ),
	.cout(Xd_0__inst_mult_11_117 ),
	.shareout(Xd_0__inst_mult_11_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_37 (
// Equation(s):
// Xd_0__inst_mult_11_120  = SUM(( (!din_a[78] & (((din_a[77] & din_b[82])))) # (din_a[78] & (!din_b[81] $ (((!din_a[77]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_114  ) + ( Xd_0__inst_mult_11_113  ))
// Xd_0__inst_mult_11_121  = CARRY(( (!din_a[78] & (((din_a[77] & din_b[82])))) # (din_a[78] & (!din_b[81] $ (((!din_a[77]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_114  ) + ( Xd_0__inst_mult_11_113  ))
// Xd_0__inst_mult_11_122  = SHARE((din_a[78] & (din_b[81] & (din_a[77] & din_b[82]))))

	.dataa(!din_a[78]),
	.datab(!din_b[81]),
	.datac(!din_a[77]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_113 ),
	.sharein(Xd_0__inst_mult_11_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_120 ),
	.cout(Xd_0__inst_mult_11_121 ),
	.shareout(Xd_0__inst_mult_11_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_36 (
// Equation(s):
// Xd_0__inst_mult_8_116  = SUM(( (!din_a[61] & (((din_a[60] & din_b[57])))) # (din_a[61] & (!din_b[56] $ (((!din_a[60]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_8_110  ) + ( Xd_0__inst_mult_8_109  ))
// Xd_0__inst_mult_8_117  = CARRY(( (!din_a[61] & (((din_a[60] & din_b[57])))) # (din_a[61] & (!din_b[56] $ (((!din_a[60]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_8_110  ) + ( Xd_0__inst_mult_8_109  ))
// Xd_0__inst_mult_8_118  = SHARE((din_a[61] & (din_b[56] & (din_a[60] & din_b[57]))))

	.dataa(!din_a[61]),
	.datab(!din_b[56]),
	.datac(!din_a[60]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_109 ),
	.sharein(Xd_0__inst_mult_8_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_116 ),
	.cout(Xd_0__inst_mult_8_117 ),
	.shareout(Xd_0__inst_mult_8_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_37 (
// Equation(s):
// Xd_0__inst_mult_8_120  = SUM(( (!din_a[57] & (((din_a[56] & din_b[61])))) # (din_a[57] & (!din_b[60] $ (((!din_a[56]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_114  ) + ( Xd_0__inst_mult_8_113  ))
// Xd_0__inst_mult_8_121  = CARRY(( (!din_a[57] & (((din_a[56] & din_b[61])))) # (din_a[57] & (!din_b[60] $ (((!din_a[56]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_114  ) + ( Xd_0__inst_mult_8_113  ))
// Xd_0__inst_mult_8_122  = SHARE((din_a[57] & (din_b[60] & (din_a[56] & din_b[61]))))

	.dataa(!din_a[57]),
	.datab(!din_b[60]),
	.datac(!din_a[56]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_113 ),
	.sharein(Xd_0__inst_mult_8_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_120 ),
	.cout(Xd_0__inst_mult_8_121 ),
	.shareout(Xd_0__inst_mult_8_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_36 (
// Equation(s):
// Xd_0__inst_mult_9_116  = SUM(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_9_110  ) + ( Xd_0__inst_mult_9_109  ))
// Xd_0__inst_mult_9_117  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_9_110  ) + ( Xd_0__inst_mult_9_109  ))
// Xd_0__inst_mult_9_118  = SHARE((din_a[68] & (din_b[63] & (din_a[67] & din_b[64]))))

	.dataa(!din_a[68]),
	.datab(!din_b[63]),
	.datac(!din_a[67]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_109 ),
	.sharein(Xd_0__inst_mult_9_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_116 ),
	.cout(Xd_0__inst_mult_9_117 ),
	.shareout(Xd_0__inst_mult_9_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_37 (
// Equation(s):
// Xd_0__inst_mult_9_120  = SUM(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_114  ) + ( Xd_0__inst_mult_9_113  ))
// Xd_0__inst_mult_9_121  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_114  ) + ( Xd_0__inst_mult_9_113  ))
// Xd_0__inst_mult_9_122  = SHARE((din_a[64] & (din_b[67] & (din_a[63] & din_b[68]))))

	.dataa(!din_a[64]),
	.datab(!din_b[67]),
	.datac(!din_a[63]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_113 ),
	.sharein(Xd_0__inst_mult_9_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_120 ),
	.cout(Xd_0__inst_mult_9_121 ),
	.shareout(Xd_0__inst_mult_9_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_36 (
// Equation(s):
// Xd_0__inst_mult_6_116  = SUM(( (!din_a[47] & (((din_a[46] & din_b[43])))) # (din_a[47] & (!din_b[42] $ (((!din_a[46]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_6_110  ) + ( Xd_0__inst_mult_6_109  ))
// Xd_0__inst_mult_6_117  = CARRY(( (!din_a[47] & (((din_a[46] & din_b[43])))) # (din_a[47] & (!din_b[42] $ (((!din_a[46]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_6_110  ) + ( Xd_0__inst_mult_6_109  ))
// Xd_0__inst_mult_6_118  = SHARE((din_a[47] & (din_b[42] & (din_a[46] & din_b[43]))))

	.dataa(!din_a[47]),
	.datab(!din_b[42]),
	.datac(!din_a[46]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_109 ),
	.sharein(Xd_0__inst_mult_6_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_116 ),
	.cout(Xd_0__inst_mult_6_117 ),
	.shareout(Xd_0__inst_mult_6_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_37 (
// Equation(s):
// Xd_0__inst_mult_6_120  = SUM(( (!din_a[43] & (((din_a[42] & din_b[47])))) # (din_a[43] & (!din_b[46] $ (((!din_a[42]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_114  ) + ( Xd_0__inst_mult_6_113  ))
// Xd_0__inst_mult_6_121  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[47])))) # (din_a[43] & (!din_b[46] $ (((!din_a[42]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_114  ) + ( Xd_0__inst_mult_6_113  ))
// Xd_0__inst_mult_6_122  = SHARE((din_a[43] & (din_b[46] & (din_a[42] & din_b[47]))))

	.dataa(!din_a[43]),
	.datab(!din_b[46]),
	.datac(!din_a[42]),
	.datad(!din_b[47]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_113 ),
	.sharein(Xd_0__inst_mult_6_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_120 ),
	.cout(Xd_0__inst_mult_6_121 ),
	.shareout(Xd_0__inst_mult_6_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_36 (
// Equation(s):
// Xd_0__inst_mult_7_116  = SUM(( (!din_a[54] & (((din_a[53] & din_b[50])))) # (din_a[54] & (!din_b[49] $ (((!din_a[53]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_7_110  ) + ( Xd_0__inst_mult_7_109  ))
// Xd_0__inst_mult_7_117  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[50])))) # (din_a[54] & (!din_b[49] $ (((!din_a[53]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_7_110  ) + ( Xd_0__inst_mult_7_109  ))
// Xd_0__inst_mult_7_118  = SHARE((din_a[54] & (din_b[49] & (din_a[53] & din_b[50]))))

	.dataa(!din_a[54]),
	.datab(!din_b[49]),
	.datac(!din_a[53]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_109 ),
	.sharein(Xd_0__inst_mult_7_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_116 ),
	.cout(Xd_0__inst_mult_7_117 ),
	.shareout(Xd_0__inst_mult_7_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_37 (
// Equation(s):
// Xd_0__inst_mult_7_120  = SUM(( (!din_a[50] & (((din_a[49] & din_b[54])))) # (din_a[50] & (!din_b[53] $ (((!din_a[49]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_114  ) + ( Xd_0__inst_mult_7_113  ))
// Xd_0__inst_mult_7_121  = CARRY(( (!din_a[50] & (((din_a[49] & din_b[54])))) # (din_a[50] & (!din_b[53] $ (((!din_a[49]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_114  ) + ( Xd_0__inst_mult_7_113  ))
// Xd_0__inst_mult_7_122  = SHARE((din_a[50] & (din_b[53] & (din_a[49] & din_b[54]))))

	.dataa(!din_a[50]),
	.datab(!din_b[53]),
	.datac(!din_a[49]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_113 ),
	.sharein(Xd_0__inst_mult_7_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_120 ),
	.cout(Xd_0__inst_mult_7_121 ),
	.shareout(Xd_0__inst_mult_7_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_36 (
// Equation(s):
// Xd_0__inst_mult_4_116  = SUM(( (!din_a[33] & (((din_a[32] & din_b[29])))) # (din_a[33] & (!din_b[28] $ (((!din_a[32]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_4_110  ) + ( Xd_0__inst_mult_4_109  ))
// Xd_0__inst_mult_4_117  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[29])))) # (din_a[33] & (!din_b[28] $ (((!din_a[32]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_4_110  ) + ( Xd_0__inst_mult_4_109  ))
// Xd_0__inst_mult_4_118  = SHARE((din_a[33] & (din_b[28] & (din_a[32] & din_b[29]))))

	.dataa(!din_a[33]),
	.datab(!din_b[28]),
	.datac(!din_a[32]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_109 ),
	.sharein(Xd_0__inst_mult_4_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_116 ),
	.cout(Xd_0__inst_mult_4_117 ),
	.shareout(Xd_0__inst_mult_4_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_37 (
// Equation(s):
// Xd_0__inst_mult_4_120  = SUM(( (!din_a[29] & (((din_a[28] & din_b[33])))) # (din_a[29] & (!din_b[32] $ (((!din_a[28]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_114  ) + ( Xd_0__inst_mult_4_113  ))
// Xd_0__inst_mult_4_121  = CARRY(( (!din_a[29] & (((din_a[28] & din_b[33])))) # (din_a[29] & (!din_b[32] $ (((!din_a[28]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_114  ) + ( Xd_0__inst_mult_4_113  ))
// Xd_0__inst_mult_4_122  = SHARE((din_a[29] & (din_b[32] & (din_a[28] & din_b[33]))))

	.dataa(!din_a[29]),
	.datab(!din_b[32]),
	.datac(!din_a[28]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_113 ),
	.sharein(Xd_0__inst_mult_4_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_120 ),
	.cout(Xd_0__inst_mult_4_121 ),
	.shareout(Xd_0__inst_mult_4_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_36 (
// Equation(s):
// Xd_0__inst_mult_5_116  = SUM(( (!din_a[40] & (((din_a[39] & din_b[36])))) # (din_a[40] & (!din_b[35] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_5_110  ) + ( Xd_0__inst_mult_5_109  ))
// Xd_0__inst_mult_5_117  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[36])))) # (din_a[40] & (!din_b[35] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_5_110  ) + ( Xd_0__inst_mult_5_109  ))
// Xd_0__inst_mult_5_118  = SHARE((din_a[40] & (din_b[35] & (din_a[39] & din_b[36]))))

	.dataa(!din_a[40]),
	.datab(!din_b[35]),
	.datac(!din_a[39]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_109 ),
	.sharein(Xd_0__inst_mult_5_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_116 ),
	.cout(Xd_0__inst_mult_5_117 ),
	.shareout(Xd_0__inst_mult_5_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_37 (
// Equation(s):
// Xd_0__inst_mult_5_120  = SUM(( (!din_a[36] & (((din_a[35] & din_b[40])))) # (din_a[36] & (!din_b[39] $ (((!din_a[35]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_114  ) + ( Xd_0__inst_mult_5_113  ))
// Xd_0__inst_mult_5_121  = CARRY(( (!din_a[36] & (((din_a[35] & din_b[40])))) # (din_a[36] & (!din_b[39] $ (((!din_a[35]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_114  ) + ( Xd_0__inst_mult_5_113  ))
// Xd_0__inst_mult_5_122  = SHARE((din_a[36] & (din_b[39] & (din_a[35] & din_b[40]))))

	.dataa(!din_a[36]),
	.datab(!din_b[39]),
	.datac(!din_a[35]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_113 ),
	.sharein(Xd_0__inst_mult_5_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_120 ),
	.cout(Xd_0__inst_mult_5_121 ),
	.shareout(Xd_0__inst_mult_5_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_36 (
// Equation(s):
// Xd_0__inst_mult_2_116  = SUM(( (!din_a[19] & (((din_a[18] & din_b[15])))) # (din_a[19] & (!din_b[14] $ (((!din_a[18]) # (!din_b[15]))))) ) + ( Xd_0__inst_mult_2_110  ) + ( Xd_0__inst_mult_2_109  ))
// Xd_0__inst_mult_2_117  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[15])))) # (din_a[19] & (!din_b[14] $ (((!din_a[18]) # (!din_b[15]))))) ) + ( Xd_0__inst_mult_2_110  ) + ( Xd_0__inst_mult_2_109  ))
// Xd_0__inst_mult_2_118  = SHARE((din_a[19] & (din_b[14] & (din_a[18] & din_b[15]))))

	.dataa(!din_a[19]),
	.datab(!din_b[14]),
	.datac(!din_a[18]),
	.datad(!din_b[15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_109 ),
	.sharein(Xd_0__inst_mult_2_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_116 ),
	.cout(Xd_0__inst_mult_2_117 ),
	.shareout(Xd_0__inst_mult_2_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_37 (
// Equation(s):
// Xd_0__inst_mult_2_120  = SUM(( (!din_a[15] & (((din_a[14] & din_b[19])))) # (din_a[15] & (!din_b[18] $ (((!din_a[14]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_114  ) + ( Xd_0__inst_mult_2_113  ))
// Xd_0__inst_mult_2_121  = CARRY(( (!din_a[15] & (((din_a[14] & din_b[19])))) # (din_a[15] & (!din_b[18] $ (((!din_a[14]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_114  ) + ( Xd_0__inst_mult_2_113  ))
// Xd_0__inst_mult_2_122  = SHARE((din_a[15] & (din_b[18] & (din_a[14] & din_b[19]))))

	.dataa(!din_a[15]),
	.datab(!din_b[18]),
	.datac(!din_a[14]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_113 ),
	.sharein(Xd_0__inst_mult_2_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_120 ),
	.cout(Xd_0__inst_mult_2_121 ),
	.shareout(Xd_0__inst_mult_2_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_36 (
// Equation(s):
// Xd_0__inst_mult_3_116  = SUM(( (!din_a[26] & (((din_a[25] & din_b[22])))) # (din_a[26] & (!din_b[21] $ (((!din_a[25]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_3_110  ) + ( Xd_0__inst_mult_3_109  ))
// Xd_0__inst_mult_3_117  = CARRY(( (!din_a[26] & (((din_a[25] & din_b[22])))) # (din_a[26] & (!din_b[21] $ (((!din_a[25]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_3_110  ) + ( Xd_0__inst_mult_3_109  ))
// Xd_0__inst_mult_3_118  = SHARE((din_a[26] & (din_b[21] & (din_a[25] & din_b[22]))))

	.dataa(!din_a[26]),
	.datab(!din_b[21]),
	.datac(!din_a[25]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_109 ),
	.sharein(Xd_0__inst_mult_3_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_116 ),
	.cout(Xd_0__inst_mult_3_117 ),
	.shareout(Xd_0__inst_mult_3_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_37 (
// Equation(s):
// Xd_0__inst_mult_3_120  = SUM(( (!din_a[22] & (((din_a[21] & din_b[26])))) # (din_a[22] & (!din_b[25] $ (((!din_a[21]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_114  ) + ( Xd_0__inst_mult_3_113  ))
// Xd_0__inst_mult_3_121  = CARRY(( (!din_a[22] & (((din_a[21] & din_b[26])))) # (din_a[22] & (!din_b[25] $ (((!din_a[21]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_114  ) + ( Xd_0__inst_mult_3_113  ))
// Xd_0__inst_mult_3_122  = SHARE((din_a[22] & (din_b[25] & (din_a[21] & din_b[26]))))

	.dataa(!din_a[22]),
	.datab(!din_b[25]),
	.datac(!din_a[21]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_113 ),
	.sharein(Xd_0__inst_mult_3_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_120 ),
	.cout(Xd_0__inst_mult_3_121 ),
	.shareout(Xd_0__inst_mult_3_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_36 (
// Equation(s):
// Xd_0__inst_mult_0_116  = SUM(( (!din_a[5] & (((din_a[4] & din_b[1])))) # (din_a[5] & (!din_b[0] $ (((!din_a[4]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_110  ) + ( Xd_0__inst_mult_0_109  ))
// Xd_0__inst_mult_0_117  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[1])))) # (din_a[5] & (!din_b[0] $ (((!din_a[4]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_110  ) + ( Xd_0__inst_mult_0_109  ))
// Xd_0__inst_mult_0_118  = SHARE((din_a[5] & (din_b[0] & (din_a[4] & din_b[1]))))

	.dataa(!din_a[5]),
	.datab(!din_b[0]),
	.datac(!din_a[4]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_109 ),
	.sharein(Xd_0__inst_mult_0_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_116 ),
	.cout(Xd_0__inst_mult_0_117 ),
	.shareout(Xd_0__inst_mult_0_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_37 (
// Equation(s):
// Xd_0__inst_mult_0_120  = SUM(( (!din_a[1] & (((din_a[0] & din_b[5])))) # (din_a[1] & (!din_b[4] $ (((!din_a[0]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_114  ) + ( Xd_0__inst_mult_0_113  ))
// Xd_0__inst_mult_0_121  = CARRY(( (!din_a[1] & (((din_a[0] & din_b[5])))) # (din_a[1] & (!din_b[4] $ (((!din_a[0]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_114  ) + ( Xd_0__inst_mult_0_113  ))
// Xd_0__inst_mult_0_122  = SHARE((din_a[1] & (din_b[4] & (din_a[0] & din_b[5]))))

	.dataa(!din_a[1]),
	.datab(!din_b[4]),
	.datac(!din_a[0]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_113 ),
	.sharein(Xd_0__inst_mult_0_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_120 ),
	.cout(Xd_0__inst_mult_0_121 ),
	.shareout(Xd_0__inst_mult_0_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_36 (
// Equation(s):
// Xd_0__inst_mult_1_116  = SUM(( (!din_a[12] & (((din_a[11] & din_b[8])))) # (din_a[12] & (!din_b[7] $ (((!din_a[11]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_110  ) + ( Xd_0__inst_mult_1_109  ))
// Xd_0__inst_mult_1_117  = CARRY(( (!din_a[12] & (((din_a[11] & din_b[8])))) # (din_a[12] & (!din_b[7] $ (((!din_a[11]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_110  ) + ( Xd_0__inst_mult_1_109  ))
// Xd_0__inst_mult_1_118  = SHARE((din_a[12] & (din_b[7] & (din_a[11] & din_b[8]))))

	.dataa(!din_a[12]),
	.datab(!din_b[7]),
	.datac(!din_a[11]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_109 ),
	.sharein(Xd_0__inst_mult_1_110 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_116 ),
	.cout(Xd_0__inst_mult_1_117 ),
	.shareout(Xd_0__inst_mult_1_118 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_37 (
// Equation(s):
// Xd_0__inst_mult_1_120  = SUM(( (!din_a[8] & (((din_a[7] & din_b[12])))) # (din_a[8] & (!din_b[11] $ (((!din_a[7]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_114  ) + ( Xd_0__inst_mult_1_113  ))
// Xd_0__inst_mult_1_121  = CARRY(( (!din_a[8] & (((din_a[7] & din_b[12])))) # (din_a[8] & (!din_b[11] $ (((!din_a[7]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_114  ) + ( Xd_0__inst_mult_1_113  ))
// Xd_0__inst_mult_1_122  = SHARE((din_a[8] & (din_b[11] & (din_a[7] & din_b[12]))))

	.dataa(!din_a[8]),
	.datab(!din_b[11]),
	.datac(!din_a[7]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_113 ),
	.sharein(Xd_0__inst_mult_1_114 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_120 ),
	.cout(Xd_0__inst_mult_1_121 ),
	.shareout(Xd_0__inst_mult_1_122 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_38 (
// Equation(s):
// Xd_0__inst_mult_28_124  = SUM(( (!din_a[201] & (((din_a[200] & din_b[198])))) # (din_a[201] & (!din_b[197] $ (((!din_a[200]) # (!din_b[198]))))) ) + ( Xd_0__inst_mult_28_118  ) + ( Xd_0__inst_mult_28_117  ))
// Xd_0__inst_mult_28_125  = CARRY(( (!din_a[201] & (((din_a[200] & din_b[198])))) # (din_a[201] & (!din_b[197] $ (((!din_a[200]) # (!din_b[198]))))) ) + ( Xd_0__inst_mult_28_118  ) + ( Xd_0__inst_mult_28_117  ))
// Xd_0__inst_mult_28_126  = SHARE((din_a[201] & (din_b[197] & (din_a[200] & din_b[198]))))

	.dataa(!din_a[201]),
	.datab(!din_b[197]),
	.datac(!din_a[200]),
	.datad(!din_b[198]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_117 ),
	.sharein(Xd_0__inst_mult_28_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_124 ),
	.cout(Xd_0__inst_mult_28_125 ),
	.shareout(Xd_0__inst_mult_28_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_39 (
// Equation(s):
// Xd_0__inst_mult_28_128  = SUM(( (!din_a[198] & (((din_a[197] & din_b[201])))) # (din_a[198] & (!din_b[200] $ (((!din_a[197]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_122  ) + ( Xd_0__inst_mult_28_121  ))
// Xd_0__inst_mult_28_129  = CARRY(( (!din_a[198] & (((din_a[197] & din_b[201])))) # (din_a[198] & (!din_b[200] $ (((!din_a[197]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_122  ) + ( Xd_0__inst_mult_28_121  ))
// Xd_0__inst_mult_28_130  = SHARE((din_a[198] & (din_b[200] & (din_a[197] & din_b[201]))))

	.dataa(!din_a[198]),
	.datab(!din_b[200]),
	.datac(!din_a[197]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_121 ),
	.sharein(Xd_0__inst_mult_28_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_128 ),
	.cout(Xd_0__inst_mult_28_129 ),
	.shareout(Xd_0__inst_mult_28_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_38 (
// Equation(s):
// Xd_0__inst_mult_29_124  = SUM(( (!din_a[208] & (((din_a[207] & din_b[205])))) # (din_a[208] & (!din_b[204] $ (((!din_a[207]) # (!din_b[205]))))) ) + ( Xd_0__inst_mult_29_118  ) + ( Xd_0__inst_mult_29_117  ))
// Xd_0__inst_mult_29_125  = CARRY(( (!din_a[208] & (((din_a[207] & din_b[205])))) # (din_a[208] & (!din_b[204] $ (((!din_a[207]) # (!din_b[205]))))) ) + ( Xd_0__inst_mult_29_118  ) + ( Xd_0__inst_mult_29_117  ))
// Xd_0__inst_mult_29_126  = SHARE((din_a[208] & (din_b[204] & (din_a[207] & din_b[205]))))

	.dataa(!din_a[208]),
	.datab(!din_b[204]),
	.datac(!din_a[207]),
	.datad(!din_b[205]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_117 ),
	.sharein(Xd_0__inst_mult_29_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_124 ),
	.cout(Xd_0__inst_mult_29_125 ),
	.shareout(Xd_0__inst_mult_29_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_39 (
// Equation(s):
// Xd_0__inst_mult_29_128  = SUM(( (!din_a[205] & (((din_a[204] & din_b[208])))) # (din_a[205] & (!din_b[207] $ (((!din_a[204]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_122  ) + ( Xd_0__inst_mult_29_121  ))
// Xd_0__inst_mult_29_129  = CARRY(( (!din_a[205] & (((din_a[204] & din_b[208])))) # (din_a[205] & (!din_b[207] $ (((!din_a[204]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_122  ) + ( Xd_0__inst_mult_29_121  ))
// Xd_0__inst_mult_29_130  = SHARE((din_a[205] & (din_b[207] & (din_a[204] & din_b[208]))))

	.dataa(!din_a[205]),
	.datab(!din_b[207]),
	.datac(!din_a[204]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_121 ),
	.sharein(Xd_0__inst_mult_29_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_128 ),
	.cout(Xd_0__inst_mult_29_129 ),
	.shareout(Xd_0__inst_mult_29_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_38 (
// Equation(s):
// Xd_0__inst_mult_26_124  = SUM(( (!din_a[187] & (((din_a[186] & din_b[184])))) # (din_a[187] & (!din_b[183] $ (((!din_a[186]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_26_118  ) + ( Xd_0__inst_mult_26_117  ))
// Xd_0__inst_mult_26_125  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[184])))) # (din_a[187] & (!din_b[183] $ (((!din_a[186]) # (!din_b[184]))))) ) + ( Xd_0__inst_mult_26_118  ) + ( Xd_0__inst_mult_26_117  ))
// Xd_0__inst_mult_26_126  = SHARE((din_a[187] & (din_b[183] & (din_a[186] & din_b[184]))))

	.dataa(!din_a[187]),
	.datab(!din_b[183]),
	.datac(!din_a[186]),
	.datad(!din_b[184]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_117 ),
	.sharein(Xd_0__inst_mult_26_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_124 ),
	.cout(Xd_0__inst_mult_26_125 ),
	.shareout(Xd_0__inst_mult_26_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_39 (
// Equation(s):
// Xd_0__inst_mult_26_128  = SUM(( (!din_a[184] & (((din_a[183] & din_b[187])))) # (din_a[184] & (!din_b[186] $ (((!din_a[183]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_122  ) + ( Xd_0__inst_mult_26_121  ))
// Xd_0__inst_mult_26_129  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[187])))) # (din_a[184] & (!din_b[186] $ (((!din_a[183]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_122  ) + ( Xd_0__inst_mult_26_121  ))
// Xd_0__inst_mult_26_130  = SHARE((din_a[184] & (din_b[186] & (din_a[183] & din_b[187]))))

	.dataa(!din_a[184]),
	.datab(!din_b[186]),
	.datac(!din_a[183]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_121 ),
	.sharein(Xd_0__inst_mult_26_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_128 ),
	.cout(Xd_0__inst_mult_26_129 ),
	.shareout(Xd_0__inst_mult_26_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_38 (
// Equation(s):
// Xd_0__inst_mult_27_124  = SUM(( (!din_a[194] & (((din_a[193] & din_b[191])))) # (din_a[194] & (!din_b[190] $ (((!din_a[193]) # (!din_b[191]))))) ) + ( Xd_0__inst_mult_27_118  ) + ( Xd_0__inst_mult_27_117  ))
// Xd_0__inst_mult_27_125  = CARRY(( (!din_a[194] & (((din_a[193] & din_b[191])))) # (din_a[194] & (!din_b[190] $ (((!din_a[193]) # (!din_b[191]))))) ) + ( Xd_0__inst_mult_27_118  ) + ( Xd_0__inst_mult_27_117  ))
// Xd_0__inst_mult_27_126  = SHARE((din_a[194] & (din_b[190] & (din_a[193] & din_b[191]))))

	.dataa(!din_a[194]),
	.datab(!din_b[190]),
	.datac(!din_a[193]),
	.datad(!din_b[191]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_117 ),
	.sharein(Xd_0__inst_mult_27_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_124 ),
	.cout(Xd_0__inst_mult_27_125 ),
	.shareout(Xd_0__inst_mult_27_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_39 (
// Equation(s):
// Xd_0__inst_mult_27_128  = SUM(( (!din_a[191] & (((din_a[190] & din_b[194])))) # (din_a[191] & (!din_b[193] $ (((!din_a[190]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_122  ) + ( Xd_0__inst_mult_27_121  ))
// Xd_0__inst_mult_27_129  = CARRY(( (!din_a[191] & (((din_a[190] & din_b[194])))) # (din_a[191] & (!din_b[193] $ (((!din_a[190]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_122  ) + ( Xd_0__inst_mult_27_121  ))
// Xd_0__inst_mult_27_130  = SHARE((din_a[191] & (din_b[193] & (din_a[190] & din_b[194]))))

	.dataa(!din_a[191]),
	.datab(!din_b[193]),
	.datac(!din_a[190]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_121 ),
	.sharein(Xd_0__inst_mult_27_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_128 ),
	.cout(Xd_0__inst_mult_27_129 ),
	.shareout(Xd_0__inst_mult_27_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_38 (
// Equation(s):
// Xd_0__inst_mult_24_124  = SUM(( (!din_a[173] & (((din_a[172] & din_b[170])))) # (din_a[173] & (!din_b[169] $ (((!din_a[172]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_24_118  ) + ( Xd_0__inst_mult_24_117  ))
// Xd_0__inst_mult_24_125  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[170])))) # (din_a[173] & (!din_b[169] $ (((!din_a[172]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_24_118  ) + ( Xd_0__inst_mult_24_117  ))
// Xd_0__inst_mult_24_126  = SHARE((din_a[173] & (din_b[169] & (din_a[172] & din_b[170]))))

	.dataa(!din_a[173]),
	.datab(!din_b[169]),
	.datac(!din_a[172]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_117 ),
	.sharein(Xd_0__inst_mult_24_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_124 ),
	.cout(Xd_0__inst_mult_24_125 ),
	.shareout(Xd_0__inst_mult_24_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_39 (
// Equation(s):
// Xd_0__inst_mult_24_128  = SUM(( (!din_a[170] & (((din_a[169] & din_b[173])))) # (din_a[170] & (!din_b[172] $ (((!din_a[169]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_122  ) + ( Xd_0__inst_mult_24_121  ))
// Xd_0__inst_mult_24_129  = CARRY(( (!din_a[170] & (((din_a[169] & din_b[173])))) # (din_a[170] & (!din_b[172] $ (((!din_a[169]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_122  ) + ( Xd_0__inst_mult_24_121  ))
// Xd_0__inst_mult_24_130  = SHARE((din_a[170] & (din_b[172] & (din_a[169] & din_b[173]))))

	.dataa(!din_a[170]),
	.datab(!din_b[172]),
	.datac(!din_a[169]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_121 ),
	.sharein(Xd_0__inst_mult_24_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_128 ),
	.cout(Xd_0__inst_mult_24_129 ),
	.shareout(Xd_0__inst_mult_24_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_39 (
// Equation(s):
// Xd_0__inst_mult_25_128  = SUM(( (!din_a[180] & (((din_a[179] & din_b[177])))) # (din_a[180] & (!din_b[176] $ (((!din_a[179]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_25_122  ) + ( Xd_0__inst_mult_25_121  ))
// Xd_0__inst_mult_25_129  = CARRY(( (!din_a[180] & (((din_a[179] & din_b[177])))) # (din_a[180] & (!din_b[176] $ (((!din_a[179]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_25_122  ) + ( Xd_0__inst_mult_25_121  ))
// Xd_0__inst_mult_25_130  = SHARE((din_a[180] & (din_b[176] & (din_a[179] & din_b[177]))))

	.dataa(!din_a[180]),
	.datab(!din_b[176]),
	.datac(!din_a[179]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_121 ),
	.sharein(Xd_0__inst_mult_25_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_128 ),
	.cout(Xd_0__inst_mult_25_129 ),
	.shareout(Xd_0__inst_mult_25_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_40 (
// Equation(s):
// Xd_0__inst_mult_25_132  = SUM(( (!din_a[177] & (((din_a[176] & din_b[180])))) # (din_a[177] & (!din_b[179] $ (((!din_a[176]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_126  ) + ( Xd_0__inst_mult_25_125  ))
// Xd_0__inst_mult_25_133  = CARRY(( (!din_a[177] & (((din_a[176] & din_b[180])))) # (din_a[177] & (!din_b[179] $ (((!din_a[176]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_126  ) + ( Xd_0__inst_mult_25_125  ))
// Xd_0__inst_mult_25_134  = SHARE((din_a[177] & (din_b[179] & (din_a[176] & din_b[180]))))

	.dataa(!din_a[177]),
	.datab(!din_b[179]),
	.datac(!din_a[176]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_125 ),
	.sharein(Xd_0__inst_mult_25_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_132 ),
	.cout(Xd_0__inst_mult_25_133 ),
	.shareout(Xd_0__inst_mult_25_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_39 (
// Equation(s):
// Xd_0__inst_mult_22_128  = SUM(( (!din_a[159] & (((din_a[158] & din_b[156])))) # (din_a[159] & (!din_b[155] $ (((!din_a[158]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_22_122  ) + ( Xd_0__inst_mult_22_121  ))
// Xd_0__inst_mult_22_129  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[156])))) # (din_a[159] & (!din_b[155] $ (((!din_a[158]) # (!din_b[156]))))) ) + ( Xd_0__inst_mult_22_122  ) + ( Xd_0__inst_mult_22_121  ))
// Xd_0__inst_mult_22_130  = SHARE((din_a[159] & (din_b[155] & (din_a[158] & din_b[156]))))

	.dataa(!din_a[159]),
	.datab(!din_b[155]),
	.datac(!din_a[158]),
	.datad(!din_b[156]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_121 ),
	.sharein(Xd_0__inst_mult_22_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_128 ),
	.cout(Xd_0__inst_mult_22_129 ),
	.shareout(Xd_0__inst_mult_22_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_40 (
// Equation(s):
// Xd_0__inst_mult_22_132  = SUM(( (!din_a[156] & (((din_a[155] & din_b[159])))) # (din_a[156] & (!din_b[158] $ (((!din_a[155]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_126  ) + ( Xd_0__inst_mult_22_125  ))
// Xd_0__inst_mult_22_133  = CARRY(( (!din_a[156] & (((din_a[155] & din_b[159])))) # (din_a[156] & (!din_b[158] $ (((!din_a[155]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_126  ) + ( Xd_0__inst_mult_22_125  ))
// Xd_0__inst_mult_22_134  = SHARE((din_a[156] & (din_b[158] & (din_a[155] & din_b[159]))))

	.dataa(!din_a[156]),
	.datab(!din_b[158]),
	.datac(!din_a[155]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_125 ),
	.sharein(Xd_0__inst_mult_22_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_132 ),
	.cout(Xd_0__inst_mult_22_133 ),
	.shareout(Xd_0__inst_mult_22_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_38 (
// Equation(s):
// Xd_0__inst_mult_23_124  = SUM(( (!din_a[166] & (((din_a[165] & din_b[163])))) # (din_a[166] & (!din_b[162] $ (((!din_a[165]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_23_118  ) + ( Xd_0__inst_mult_23_117  ))
// Xd_0__inst_mult_23_125  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[163])))) # (din_a[166] & (!din_b[162] $ (((!din_a[165]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_23_118  ) + ( Xd_0__inst_mult_23_117  ))
// Xd_0__inst_mult_23_126  = SHARE((din_a[166] & (din_b[162] & (din_a[165] & din_b[163]))))

	.dataa(!din_a[166]),
	.datab(!din_b[162]),
	.datac(!din_a[165]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_117 ),
	.sharein(Xd_0__inst_mult_23_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_124 ),
	.cout(Xd_0__inst_mult_23_125 ),
	.shareout(Xd_0__inst_mult_23_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_39 (
// Equation(s):
// Xd_0__inst_mult_23_128  = SUM(( (!din_a[163] & (((din_a[162] & din_b[166])))) # (din_a[163] & (!din_b[165] $ (((!din_a[162]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_122  ) + ( Xd_0__inst_mult_23_121  ))
// Xd_0__inst_mult_23_129  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[166])))) # (din_a[163] & (!din_b[165] $ (((!din_a[162]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_122  ) + ( Xd_0__inst_mult_23_121  ))
// Xd_0__inst_mult_23_130  = SHARE((din_a[163] & (din_b[165] & (din_a[162] & din_b[166]))))

	.dataa(!din_a[163]),
	.datab(!din_b[165]),
	.datac(!din_a[162]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_121 ),
	.sharein(Xd_0__inst_mult_23_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_128 ),
	.cout(Xd_0__inst_mult_23_129 ),
	.shareout(Xd_0__inst_mult_23_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_38 (
// Equation(s):
// Xd_0__inst_mult_20_124  = SUM(( (!din_a[145] & (((din_a[144] & din_b[142])))) # (din_a[145] & (!din_b[141] $ (((!din_a[144]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_20_118  ) + ( Xd_0__inst_mult_20_117  ))
// Xd_0__inst_mult_20_125  = CARRY(( (!din_a[145] & (((din_a[144] & din_b[142])))) # (din_a[145] & (!din_b[141] $ (((!din_a[144]) # (!din_b[142]))))) ) + ( Xd_0__inst_mult_20_118  ) + ( Xd_0__inst_mult_20_117  ))
// Xd_0__inst_mult_20_126  = SHARE((din_a[145] & (din_b[141] & (din_a[144] & din_b[142]))))

	.dataa(!din_a[145]),
	.datab(!din_b[141]),
	.datac(!din_a[144]),
	.datad(!din_b[142]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_117 ),
	.sharein(Xd_0__inst_mult_20_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_124 ),
	.cout(Xd_0__inst_mult_20_125 ),
	.shareout(Xd_0__inst_mult_20_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_39 (
// Equation(s):
// Xd_0__inst_mult_20_128  = SUM(( (!din_a[142] & (((din_a[141] & din_b[145])))) # (din_a[142] & (!din_b[144] $ (((!din_a[141]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_122  ) + ( Xd_0__inst_mult_20_121  ))
// Xd_0__inst_mult_20_129  = CARRY(( (!din_a[142] & (((din_a[141] & din_b[145])))) # (din_a[142] & (!din_b[144] $ (((!din_a[141]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_122  ) + ( Xd_0__inst_mult_20_121  ))
// Xd_0__inst_mult_20_130  = SHARE((din_a[142] & (din_b[144] & (din_a[141] & din_b[145]))))

	.dataa(!din_a[142]),
	.datab(!din_b[144]),
	.datac(!din_a[141]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_121 ),
	.sharein(Xd_0__inst_mult_20_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_128 ),
	.cout(Xd_0__inst_mult_20_129 ),
	.shareout(Xd_0__inst_mult_20_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_38 (
// Equation(s):
// Xd_0__inst_mult_21_124  = SUM(( (!din_a[152] & (((din_a[151] & din_b[149])))) # (din_a[152] & (!din_b[148] $ (((!din_a[151]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_21_118  ) + ( Xd_0__inst_mult_21_117  ))
// Xd_0__inst_mult_21_125  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[149])))) # (din_a[152] & (!din_b[148] $ (((!din_a[151]) # (!din_b[149]))))) ) + ( Xd_0__inst_mult_21_118  ) + ( Xd_0__inst_mult_21_117  ))
// Xd_0__inst_mult_21_126  = SHARE((din_a[152] & (din_b[148] & (din_a[151] & din_b[149]))))

	.dataa(!din_a[152]),
	.datab(!din_b[148]),
	.datac(!din_a[151]),
	.datad(!din_b[149]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_117 ),
	.sharein(Xd_0__inst_mult_21_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_124 ),
	.cout(Xd_0__inst_mult_21_125 ),
	.shareout(Xd_0__inst_mult_21_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_39 (
// Equation(s):
// Xd_0__inst_mult_21_128  = SUM(( (!din_a[149] & (((din_a[148] & din_b[152])))) # (din_a[149] & (!din_b[151] $ (((!din_a[148]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_122  ) + ( Xd_0__inst_mult_21_121  ))
// Xd_0__inst_mult_21_129  = CARRY(( (!din_a[149] & (((din_a[148] & din_b[152])))) # (din_a[149] & (!din_b[151] $ (((!din_a[148]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_122  ) + ( Xd_0__inst_mult_21_121  ))
// Xd_0__inst_mult_21_130  = SHARE((din_a[149] & (din_b[151] & (din_a[148] & din_b[152]))))

	.dataa(!din_a[149]),
	.datab(!din_b[151]),
	.datac(!din_a[148]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_121 ),
	.sharein(Xd_0__inst_mult_21_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_128 ),
	.cout(Xd_0__inst_mult_21_129 ),
	.shareout(Xd_0__inst_mult_21_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_38 (
// Equation(s):
// Xd_0__inst_mult_18_124  = SUM(( (!din_a[131] & (((din_a[130] & din_b[128])))) # (din_a[131] & (!din_b[127] $ (((!din_a[130]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_18_118  ) + ( Xd_0__inst_mult_18_117  ))
// Xd_0__inst_mult_18_125  = CARRY(( (!din_a[131] & (((din_a[130] & din_b[128])))) # (din_a[131] & (!din_b[127] $ (((!din_a[130]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_18_118  ) + ( Xd_0__inst_mult_18_117  ))
// Xd_0__inst_mult_18_126  = SHARE((din_a[131] & (din_b[127] & (din_a[130] & din_b[128]))))

	.dataa(!din_a[131]),
	.datab(!din_b[127]),
	.datac(!din_a[130]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_117 ),
	.sharein(Xd_0__inst_mult_18_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_124 ),
	.cout(Xd_0__inst_mult_18_125 ),
	.shareout(Xd_0__inst_mult_18_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_39 (
// Equation(s):
// Xd_0__inst_mult_18_128  = SUM(( (!din_a[128] & (((din_a[127] & din_b[131])))) # (din_a[128] & (!din_b[130] $ (((!din_a[127]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_122  ) + ( Xd_0__inst_mult_18_121  ))
// Xd_0__inst_mult_18_129  = CARRY(( (!din_a[128] & (((din_a[127] & din_b[131])))) # (din_a[128] & (!din_b[130] $ (((!din_a[127]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_122  ) + ( Xd_0__inst_mult_18_121  ))
// Xd_0__inst_mult_18_130  = SHARE((din_a[128] & (din_b[130] & (din_a[127] & din_b[131]))))

	.dataa(!din_a[128]),
	.datab(!din_b[130]),
	.datac(!din_a[127]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_121 ),
	.sharein(Xd_0__inst_mult_18_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_128 ),
	.cout(Xd_0__inst_mult_18_129 ),
	.shareout(Xd_0__inst_mult_18_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_38 (
// Equation(s):
// Xd_0__inst_mult_19_124  = SUM(( (!din_a[138] & (((din_a[137] & din_b[135])))) # (din_a[138] & (!din_b[134] $ (((!din_a[137]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_19_118  ) + ( Xd_0__inst_mult_19_117  ))
// Xd_0__inst_mult_19_125  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[135])))) # (din_a[138] & (!din_b[134] $ (((!din_a[137]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_19_118  ) + ( Xd_0__inst_mult_19_117  ))
// Xd_0__inst_mult_19_126  = SHARE((din_a[138] & (din_b[134] & (din_a[137] & din_b[135]))))

	.dataa(!din_a[138]),
	.datab(!din_b[134]),
	.datac(!din_a[137]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_117 ),
	.sharein(Xd_0__inst_mult_19_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_124 ),
	.cout(Xd_0__inst_mult_19_125 ),
	.shareout(Xd_0__inst_mult_19_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_39 (
// Equation(s):
// Xd_0__inst_mult_19_128  = SUM(( (!din_a[135] & (((din_a[134] & din_b[138])))) # (din_a[135] & (!din_b[137] $ (((!din_a[134]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_122  ) + ( Xd_0__inst_mult_19_121  ))
// Xd_0__inst_mult_19_129  = CARRY(( (!din_a[135] & (((din_a[134] & din_b[138])))) # (din_a[135] & (!din_b[137] $ (((!din_a[134]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_122  ) + ( Xd_0__inst_mult_19_121  ))
// Xd_0__inst_mult_19_130  = SHARE((din_a[135] & (din_b[137] & (din_a[134] & din_b[138]))))

	.dataa(!din_a[135]),
	.datab(!din_b[137]),
	.datac(!din_a[134]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_121 ),
	.sharein(Xd_0__inst_mult_19_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_128 ),
	.cout(Xd_0__inst_mult_19_129 ),
	.shareout(Xd_0__inst_mult_19_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_38 (
// Equation(s):
// Xd_0__inst_mult_16_124  = SUM(( (!din_a[117] & (((din_a[116] & din_b[114])))) # (din_a[117] & (!din_b[113] $ (((!din_a[116]) # (!din_b[114]))))) ) + ( Xd_0__inst_mult_16_118  ) + ( Xd_0__inst_mult_16_117  ))
// Xd_0__inst_mult_16_125  = CARRY(( (!din_a[117] & (((din_a[116] & din_b[114])))) # (din_a[117] & (!din_b[113] $ (((!din_a[116]) # (!din_b[114]))))) ) + ( Xd_0__inst_mult_16_118  ) + ( Xd_0__inst_mult_16_117  ))
// Xd_0__inst_mult_16_126  = SHARE((din_a[117] & (din_b[113] & (din_a[116] & din_b[114]))))

	.dataa(!din_a[117]),
	.datab(!din_b[113]),
	.datac(!din_a[116]),
	.datad(!din_b[114]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_117 ),
	.sharein(Xd_0__inst_mult_16_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_124 ),
	.cout(Xd_0__inst_mult_16_125 ),
	.shareout(Xd_0__inst_mult_16_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_39 (
// Equation(s):
// Xd_0__inst_mult_16_128  = SUM(( (!din_a[114] & (((din_a[113] & din_b[117])))) # (din_a[114] & (!din_b[116] $ (((!din_a[113]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_122  ) + ( Xd_0__inst_mult_16_121  ))
// Xd_0__inst_mult_16_129  = CARRY(( (!din_a[114] & (((din_a[113] & din_b[117])))) # (din_a[114] & (!din_b[116] $ (((!din_a[113]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_122  ) + ( Xd_0__inst_mult_16_121  ))
// Xd_0__inst_mult_16_130  = SHARE((din_a[114] & (din_b[116] & (din_a[113] & din_b[117]))))

	.dataa(!din_a[114]),
	.datab(!din_b[116]),
	.datac(!din_a[113]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_121 ),
	.sharein(Xd_0__inst_mult_16_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_128 ),
	.cout(Xd_0__inst_mult_16_129 ),
	.shareout(Xd_0__inst_mult_16_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_38 (
// Equation(s):
// Xd_0__inst_mult_17_124  = SUM(( (!din_a[124] & (((din_a[123] & din_b[121])))) # (din_a[124] & (!din_b[120] $ (((!din_a[123]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_17_118  ) + ( Xd_0__inst_mult_17_117  ))
// Xd_0__inst_mult_17_125  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[121])))) # (din_a[124] & (!din_b[120] $ (((!din_a[123]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_17_118  ) + ( Xd_0__inst_mult_17_117  ))
// Xd_0__inst_mult_17_126  = SHARE((din_a[124] & (din_b[120] & (din_a[123] & din_b[121]))))

	.dataa(!din_a[124]),
	.datab(!din_b[120]),
	.datac(!din_a[123]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_117 ),
	.sharein(Xd_0__inst_mult_17_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_124 ),
	.cout(Xd_0__inst_mult_17_125 ),
	.shareout(Xd_0__inst_mult_17_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_39 (
// Equation(s):
// Xd_0__inst_mult_17_128  = SUM(( (!din_a[121] & (((din_a[120] & din_b[124])))) # (din_a[121] & (!din_b[123] $ (((!din_a[120]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_122  ) + ( Xd_0__inst_mult_17_121  ))
// Xd_0__inst_mult_17_129  = CARRY(( (!din_a[121] & (((din_a[120] & din_b[124])))) # (din_a[121] & (!din_b[123] $ (((!din_a[120]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_122  ) + ( Xd_0__inst_mult_17_121  ))
// Xd_0__inst_mult_17_130  = SHARE((din_a[121] & (din_b[123] & (din_a[120] & din_b[124]))))

	.dataa(!din_a[121]),
	.datab(!din_b[123]),
	.datac(!din_a[120]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_121 ),
	.sharein(Xd_0__inst_mult_17_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_128 ),
	.cout(Xd_0__inst_mult_17_129 ),
	.shareout(Xd_0__inst_mult_17_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_38 (
// Equation(s):
// Xd_0__inst_mult_14_124  = SUM(( (!din_a[103] & (((din_a[102] & din_b[100])))) # (din_a[103] & (!din_b[99] $ (((!din_a[102]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_14_118  ) + ( Xd_0__inst_mult_14_117  ))
// Xd_0__inst_mult_14_125  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[100])))) # (din_a[103] & (!din_b[99] $ (((!din_a[102]) # (!din_b[100]))))) ) + ( Xd_0__inst_mult_14_118  ) + ( Xd_0__inst_mult_14_117  ))
// Xd_0__inst_mult_14_126  = SHARE((din_a[103] & (din_b[99] & (din_a[102] & din_b[100]))))

	.dataa(!din_a[103]),
	.datab(!din_b[99]),
	.datac(!din_a[102]),
	.datad(!din_b[100]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_117 ),
	.sharein(Xd_0__inst_mult_14_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_124 ),
	.cout(Xd_0__inst_mult_14_125 ),
	.shareout(Xd_0__inst_mult_14_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_39 (
// Equation(s):
// Xd_0__inst_mult_14_128  = SUM(( (!din_a[100] & (((din_a[99] & din_b[103])))) # (din_a[100] & (!din_b[102] $ (((!din_a[99]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_122  ) + ( Xd_0__inst_mult_14_121  ))
// Xd_0__inst_mult_14_129  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[103])))) # (din_a[100] & (!din_b[102] $ (((!din_a[99]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_122  ) + ( Xd_0__inst_mult_14_121  ))
// Xd_0__inst_mult_14_130  = SHARE((din_a[100] & (din_b[102] & (din_a[99] & din_b[103]))))

	.dataa(!din_a[100]),
	.datab(!din_b[102]),
	.datac(!din_a[99]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_121 ),
	.sharein(Xd_0__inst_mult_14_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_128 ),
	.cout(Xd_0__inst_mult_14_129 ),
	.shareout(Xd_0__inst_mult_14_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_38 (
// Equation(s):
// Xd_0__inst_mult_15_124  = SUM(( (!din_a[110] & (((din_a[109] & din_b[107])))) # (din_a[110] & (!din_b[106] $ (((!din_a[109]) # (!din_b[107]))))) ) + ( Xd_0__inst_mult_15_118  ) + ( Xd_0__inst_mult_15_117  ))
// Xd_0__inst_mult_15_125  = CARRY(( (!din_a[110] & (((din_a[109] & din_b[107])))) # (din_a[110] & (!din_b[106] $ (((!din_a[109]) # (!din_b[107]))))) ) + ( Xd_0__inst_mult_15_118  ) + ( Xd_0__inst_mult_15_117  ))
// Xd_0__inst_mult_15_126  = SHARE((din_a[110] & (din_b[106] & (din_a[109] & din_b[107]))))

	.dataa(!din_a[110]),
	.datab(!din_b[106]),
	.datac(!din_a[109]),
	.datad(!din_b[107]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_117 ),
	.sharein(Xd_0__inst_mult_15_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_124 ),
	.cout(Xd_0__inst_mult_15_125 ),
	.shareout(Xd_0__inst_mult_15_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_39 (
// Equation(s):
// Xd_0__inst_mult_15_128  = SUM(( (!din_a[107] & (((din_a[106] & din_b[110])))) # (din_a[107] & (!din_b[109] $ (((!din_a[106]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_122  ) + ( Xd_0__inst_mult_15_121  ))
// Xd_0__inst_mult_15_129  = CARRY(( (!din_a[107] & (((din_a[106] & din_b[110])))) # (din_a[107] & (!din_b[109] $ (((!din_a[106]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_122  ) + ( Xd_0__inst_mult_15_121  ))
// Xd_0__inst_mult_15_130  = SHARE((din_a[107] & (din_b[109] & (din_a[106] & din_b[110]))))

	.dataa(!din_a[107]),
	.datab(!din_b[109]),
	.datac(!din_a[106]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_121 ),
	.sharein(Xd_0__inst_mult_15_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_128 ),
	.cout(Xd_0__inst_mult_15_129 ),
	.shareout(Xd_0__inst_mult_15_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_38 (
// Equation(s):
// Xd_0__inst_mult_12_124  = SUM(( (!din_a[89] & (((din_a[88] & din_b[86])))) # (din_a[89] & (!din_b[85] $ (((!din_a[88]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_12_118  ) + ( Xd_0__inst_mult_12_117  ))
// Xd_0__inst_mult_12_125  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[86])))) # (din_a[89] & (!din_b[85] $ (((!din_a[88]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_12_118  ) + ( Xd_0__inst_mult_12_117  ))
// Xd_0__inst_mult_12_126  = SHARE((din_a[89] & (din_b[85] & (din_a[88] & din_b[86]))))

	.dataa(!din_a[89]),
	.datab(!din_b[85]),
	.datac(!din_a[88]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_117 ),
	.sharein(Xd_0__inst_mult_12_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_124 ),
	.cout(Xd_0__inst_mult_12_125 ),
	.shareout(Xd_0__inst_mult_12_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_39 (
// Equation(s):
// Xd_0__inst_mult_12_128  = SUM(( (!din_a[86] & (((din_a[85] & din_b[89])))) # (din_a[86] & (!din_b[88] $ (((!din_a[85]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_122  ) + ( Xd_0__inst_mult_12_121  ))
// Xd_0__inst_mult_12_129  = CARRY(( (!din_a[86] & (((din_a[85] & din_b[89])))) # (din_a[86] & (!din_b[88] $ (((!din_a[85]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_122  ) + ( Xd_0__inst_mult_12_121  ))
// Xd_0__inst_mult_12_130  = SHARE((din_a[86] & (din_b[88] & (din_a[85] & din_b[89]))))

	.dataa(!din_a[86]),
	.datab(!din_b[88]),
	.datac(!din_a[85]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_121 ),
	.sharein(Xd_0__inst_mult_12_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_128 ),
	.cout(Xd_0__inst_mult_12_129 ),
	.shareout(Xd_0__inst_mult_12_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_38 (
// Equation(s):
// Xd_0__inst_mult_13_124  = SUM(( (!din_a[96] & (((din_a[95] & din_b[93])))) # (din_a[96] & (!din_b[92] $ (((!din_a[95]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_13_118  ) + ( Xd_0__inst_mult_13_117  ))
// Xd_0__inst_mult_13_125  = CARRY(( (!din_a[96] & (((din_a[95] & din_b[93])))) # (din_a[96] & (!din_b[92] $ (((!din_a[95]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_13_118  ) + ( Xd_0__inst_mult_13_117  ))
// Xd_0__inst_mult_13_126  = SHARE((din_a[96] & (din_b[92] & (din_a[95] & din_b[93]))))

	.dataa(!din_a[96]),
	.datab(!din_b[92]),
	.datac(!din_a[95]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_117 ),
	.sharein(Xd_0__inst_mult_13_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_124 ),
	.cout(Xd_0__inst_mult_13_125 ),
	.shareout(Xd_0__inst_mult_13_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_39 (
// Equation(s):
// Xd_0__inst_mult_13_128  = SUM(( (!din_a[93] & (((din_a[92] & din_b[96])))) # (din_a[93] & (!din_b[95] $ (((!din_a[92]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_122  ) + ( Xd_0__inst_mult_13_121  ))
// Xd_0__inst_mult_13_129  = CARRY(( (!din_a[93] & (((din_a[92] & din_b[96])))) # (din_a[93] & (!din_b[95] $ (((!din_a[92]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_122  ) + ( Xd_0__inst_mult_13_121  ))
// Xd_0__inst_mult_13_130  = SHARE((din_a[93] & (din_b[95] & (din_a[92] & din_b[96]))))

	.dataa(!din_a[93]),
	.datab(!din_b[95]),
	.datac(!din_a[92]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_121 ),
	.sharein(Xd_0__inst_mult_13_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_128 ),
	.cout(Xd_0__inst_mult_13_129 ),
	.shareout(Xd_0__inst_mult_13_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_38 (
// Equation(s):
// Xd_0__inst_mult_10_124  = SUM(( (!din_a[75] & (((din_a[74] & din_b[72])))) # (din_a[75] & (!din_b[71] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_10_118  ) + ( Xd_0__inst_mult_10_117  ))
// Xd_0__inst_mult_10_125  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[72])))) # (din_a[75] & (!din_b[71] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_10_118  ) + ( Xd_0__inst_mult_10_117  ))
// Xd_0__inst_mult_10_126  = SHARE((din_a[75] & (din_b[71] & (din_a[74] & din_b[72]))))

	.dataa(!din_a[75]),
	.datab(!din_b[71]),
	.datac(!din_a[74]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_117 ),
	.sharein(Xd_0__inst_mult_10_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_124 ),
	.cout(Xd_0__inst_mult_10_125 ),
	.shareout(Xd_0__inst_mult_10_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_39 (
// Equation(s):
// Xd_0__inst_mult_10_128  = SUM(( (!din_a[72] & (((din_a[71] & din_b[75])))) # (din_a[72] & (!din_b[74] $ (((!din_a[71]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_122  ) + ( Xd_0__inst_mult_10_121  ))
// Xd_0__inst_mult_10_129  = CARRY(( (!din_a[72] & (((din_a[71] & din_b[75])))) # (din_a[72] & (!din_b[74] $ (((!din_a[71]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_122  ) + ( Xd_0__inst_mult_10_121  ))
// Xd_0__inst_mult_10_130  = SHARE((din_a[72] & (din_b[74] & (din_a[71] & din_b[75]))))

	.dataa(!din_a[72]),
	.datab(!din_b[74]),
	.datac(!din_a[71]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_121 ),
	.sharein(Xd_0__inst_mult_10_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_128 ),
	.cout(Xd_0__inst_mult_10_129 ),
	.shareout(Xd_0__inst_mult_10_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_38 (
// Equation(s):
// Xd_0__inst_mult_11_124  = SUM(( (!din_a[82] & (((din_a[81] & din_b[79])))) # (din_a[82] & (!din_b[78] $ (((!din_a[81]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_11_118  ) + ( Xd_0__inst_mult_11_117  ))
// Xd_0__inst_mult_11_125  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[79])))) # (din_a[82] & (!din_b[78] $ (((!din_a[81]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_11_118  ) + ( Xd_0__inst_mult_11_117  ))
// Xd_0__inst_mult_11_126  = SHARE((din_a[82] & (din_b[78] & (din_a[81] & din_b[79]))))

	.dataa(!din_a[82]),
	.datab(!din_b[78]),
	.datac(!din_a[81]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_117 ),
	.sharein(Xd_0__inst_mult_11_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_124 ),
	.cout(Xd_0__inst_mult_11_125 ),
	.shareout(Xd_0__inst_mult_11_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_39 (
// Equation(s):
// Xd_0__inst_mult_11_128  = SUM(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_122  ) + ( Xd_0__inst_mult_11_121  ))
// Xd_0__inst_mult_11_129  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_122  ) + ( Xd_0__inst_mult_11_121  ))
// Xd_0__inst_mult_11_130  = SHARE((din_a[79] & (din_b[81] & (din_a[78] & din_b[82]))))

	.dataa(!din_a[79]),
	.datab(!din_b[81]),
	.datac(!din_a[78]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_121 ),
	.sharein(Xd_0__inst_mult_11_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_128 ),
	.cout(Xd_0__inst_mult_11_129 ),
	.shareout(Xd_0__inst_mult_11_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_38 (
// Equation(s):
// Xd_0__inst_mult_8_124  = SUM(( (!din_a[61] & (((din_a[60] & din_b[58])))) # (din_a[61] & (!din_b[57] $ (((!din_a[60]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_8_118  ) + ( Xd_0__inst_mult_8_117  ))
// Xd_0__inst_mult_8_125  = CARRY(( (!din_a[61] & (((din_a[60] & din_b[58])))) # (din_a[61] & (!din_b[57] $ (((!din_a[60]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_8_118  ) + ( Xd_0__inst_mult_8_117  ))
// Xd_0__inst_mult_8_126  = SHARE((din_a[61] & (din_b[57] & (din_a[60] & din_b[58]))))

	.dataa(!din_a[61]),
	.datab(!din_b[57]),
	.datac(!din_a[60]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_117 ),
	.sharein(Xd_0__inst_mult_8_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_124 ),
	.cout(Xd_0__inst_mult_8_125 ),
	.shareout(Xd_0__inst_mult_8_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_39 (
// Equation(s):
// Xd_0__inst_mult_8_128  = SUM(( (!din_a[58] & (((din_a[57] & din_b[61])))) # (din_a[58] & (!din_b[60] $ (((!din_a[57]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_122  ) + ( Xd_0__inst_mult_8_121  ))
// Xd_0__inst_mult_8_129  = CARRY(( (!din_a[58] & (((din_a[57] & din_b[61])))) # (din_a[58] & (!din_b[60] $ (((!din_a[57]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_122  ) + ( Xd_0__inst_mult_8_121  ))
// Xd_0__inst_mult_8_130  = SHARE((din_a[58] & (din_b[60] & (din_a[57] & din_b[61]))))

	.dataa(!din_a[58]),
	.datab(!din_b[60]),
	.datac(!din_a[57]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_121 ),
	.sharein(Xd_0__inst_mult_8_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_128 ),
	.cout(Xd_0__inst_mult_8_129 ),
	.shareout(Xd_0__inst_mult_8_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_38 (
// Equation(s):
// Xd_0__inst_mult_9_124  = SUM(( (!din_a[68] & (((din_a[67] & din_b[65])))) # (din_a[68] & (!din_b[64] $ (((!din_a[67]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_9_118  ) + ( Xd_0__inst_mult_9_117  ))
// Xd_0__inst_mult_9_125  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[65])))) # (din_a[68] & (!din_b[64] $ (((!din_a[67]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_9_118  ) + ( Xd_0__inst_mult_9_117  ))
// Xd_0__inst_mult_9_126  = SHARE((din_a[68] & (din_b[64] & (din_a[67] & din_b[65]))))

	.dataa(!din_a[68]),
	.datab(!din_b[64]),
	.datac(!din_a[67]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_117 ),
	.sharein(Xd_0__inst_mult_9_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_124 ),
	.cout(Xd_0__inst_mult_9_125 ),
	.shareout(Xd_0__inst_mult_9_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_39 (
// Equation(s):
// Xd_0__inst_mult_9_128  = SUM(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_122  ) + ( Xd_0__inst_mult_9_121  ))
// Xd_0__inst_mult_9_129  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_122  ) + ( Xd_0__inst_mult_9_121  ))
// Xd_0__inst_mult_9_130  = SHARE((din_a[65] & (din_b[67] & (din_a[64] & din_b[68]))))

	.dataa(!din_a[65]),
	.datab(!din_b[67]),
	.datac(!din_a[64]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_121 ),
	.sharein(Xd_0__inst_mult_9_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_128 ),
	.cout(Xd_0__inst_mult_9_129 ),
	.shareout(Xd_0__inst_mult_9_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_38 (
// Equation(s):
// Xd_0__inst_mult_6_124  = SUM(( (!din_a[47] & (((din_a[46] & din_b[44])))) # (din_a[47] & (!din_b[43] $ (((!din_a[46]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_6_118  ) + ( Xd_0__inst_mult_6_117  ))
// Xd_0__inst_mult_6_125  = CARRY(( (!din_a[47] & (((din_a[46] & din_b[44])))) # (din_a[47] & (!din_b[43] $ (((!din_a[46]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_6_118  ) + ( Xd_0__inst_mult_6_117  ))
// Xd_0__inst_mult_6_126  = SHARE((din_a[47] & (din_b[43] & (din_a[46] & din_b[44]))))

	.dataa(!din_a[47]),
	.datab(!din_b[43]),
	.datac(!din_a[46]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_117 ),
	.sharein(Xd_0__inst_mult_6_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_124 ),
	.cout(Xd_0__inst_mult_6_125 ),
	.shareout(Xd_0__inst_mult_6_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_39 (
// Equation(s):
// Xd_0__inst_mult_6_128  = SUM(( (!din_a[44] & (((din_a[43] & din_b[47])))) # (din_a[44] & (!din_b[46] $ (((!din_a[43]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_122  ) + ( Xd_0__inst_mult_6_121  ))
// Xd_0__inst_mult_6_129  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[47])))) # (din_a[44] & (!din_b[46] $ (((!din_a[43]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_122  ) + ( Xd_0__inst_mult_6_121  ))
// Xd_0__inst_mult_6_130  = SHARE((din_a[44] & (din_b[46] & (din_a[43] & din_b[47]))))

	.dataa(!din_a[44]),
	.datab(!din_b[46]),
	.datac(!din_a[43]),
	.datad(!din_b[47]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_121 ),
	.sharein(Xd_0__inst_mult_6_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_128 ),
	.cout(Xd_0__inst_mult_6_129 ),
	.shareout(Xd_0__inst_mult_6_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_38 (
// Equation(s):
// Xd_0__inst_mult_7_124  = SUM(( (!din_a[54] & (((din_a[53] & din_b[51])))) # (din_a[54] & (!din_b[50] $ (((!din_a[53]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_7_118  ) + ( Xd_0__inst_mult_7_117  ))
// Xd_0__inst_mult_7_125  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[51])))) # (din_a[54] & (!din_b[50] $ (((!din_a[53]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_7_118  ) + ( Xd_0__inst_mult_7_117  ))
// Xd_0__inst_mult_7_126  = SHARE((din_a[54] & (din_b[50] & (din_a[53] & din_b[51]))))

	.dataa(!din_a[54]),
	.datab(!din_b[50]),
	.datac(!din_a[53]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_117 ),
	.sharein(Xd_0__inst_mult_7_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_124 ),
	.cout(Xd_0__inst_mult_7_125 ),
	.shareout(Xd_0__inst_mult_7_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_39 (
// Equation(s):
// Xd_0__inst_mult_7_128  = SUM(( (!din_a[51] & (((din_a[50] & din_b[54])))) # (din_a[51] & (!din_b[53] $ (((!din_a[50]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_122  ) + ( Xd_0__inst_mult_7_121  ))
// Xd_0__inst_mult_7_129  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[54])))) # (din_a[51] & (!din_b[53] $ (((!din_a[50]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_122  ) + ( Xd_0__inst_mult_7_121  ))
// Xd_0__inst_mult_7_130  = SHARE((din_a[51] & (din_b[53] & (din_a[50] & din_b[54]))))

	.dataa(!din_a[51]),
	.datab(!din_b[53]),
	.datac(!din_a[50]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_121 ),
	.sharein(Xd_0__inst_mult_7_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_128 ),
	.cout(Xd_0__inst_mult_7_129 ),
	.shareout(Xd_0__inst_mult_7_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_38 (
// Equation(s):
// Xd_0__inst_mult_4_124  = SUM(( (!din_a[33] & (((din_a[32] & din_b[30])))) # (din_a[33] & (!din_b[29] $ (((!din_a[32]) # (!din_b[30]))))) ) + ( Xd_0__inst_mult_4_118  ) + ( Xd_0__inst_mult_4_117  ))
// Xd_0__inst_mult_4_125  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[30])))) # (din_a[33] & (!din_b[29] $ (((!din_a[32]) # (!din_b[30]))))) ) + ( Xd_0__inst_mult_4_118  ) + ( Xd_0__inst_mult_4_117  ))
// Xd_0__inst_mult_4_126  = SHARE((din_a[33] & (din_b[29] & (din_a[32] & din_b[30]))))

	.dataa(!din_a[33]),
	.datab(!din_b[29]),
	.datac(!din_a[32]),
	.datad(!din_b[30]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_117 ),
	.sharein(Xd_0__inst_mult_4_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_124 ),
	.cout(Xd_0__inst_mult_4_125 ),
	.shareout(Xd_0__inst_mult_4_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_39 (
// Equation(s):
// Xd_0__inst_mult_4_128  = SUM(( (!din_a[30] & (((din_a[29] & din_b[33])))) # (din_a[30] & (!din_b[32] $ (((!din_a[29]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_122  ) + ( Xd_0__inst_mult_4_121  ))
// Xd_0__inst_mult_4_129  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[33])))) # (din_a[30] & (!din_b[32] $ (((!din_a[29]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_122  ) + ( Xd_0__inst_mult_4_121  ))
// Xd_0__inst_mult_4_130  = SHARE((din_a[30] & (din_b[32] & (din_a[29] & din_b[33]))))

	.dataa(!din_a[30]),
	.datab(!din_b[32]),
	.datac(!din_a[29]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_121 ),
	.sharein(Xd_0__inst_mult_4_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_128 ),
	.cout(Xd_0__inst_mult_4_129 ),
	.shareout(Xd_0__inst_mult_4_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_38 (
// Equation(s):
// Xd_0__inst_mult_5_124  = SUM(( (!din_a[40] & (((din_a[39] & din_b[37])))) # (din_a[40] & (!din_b[36] $ (((!din_a[39]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_5_118  ) + ( Xd_0__inst_mult_5_117  ))
// Xd_0__inst_mult_5_125  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[37])))) # (din_a[40] & (!din_b[36] $ (((!din_a[39]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_5_118  ) + ( Xd_0__inst_mult_5_117  ))
// Xd_0__inst_mult_5_126  = SHARE((din_a[40] & (din_b[36] & (din_a[39] & din_b[37]))))

	.dataa(!din_a[40]),
	.datab(!din_b[36]),
	.datac(!din_a[39]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_117 ),
	.sharein(Xd_0__inst_mult_5_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_124 ),
	.cout(Xd_0__inst_mult_5_125 ),
	.shareout(Xd_0__inst_mult_5_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_39 (
// Equation(s):
// Xd_0__inst_mult_5_128  = SUM(( (!din_a[37] & (((din_a[36] & din_b[40])))) # (din_a[37] & (!din_b[39] $ (((!din_a[36]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_122  ) + ( Xd_0__inst_mult_5_121  ))
// Xd_0__inst_mult_5_129  = CARRY(( (!din_a[37] & (((din_a[36] & din_b[40])))) # (din_a[37] & (!din_b[39] $ (((!din_a[36]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_122  ) + ( Xd_0__inst_mult_5_121  ))
// Xd_0__inst_mult_5_130  = SHARE((din_a[37] & (din_b[39] & (din_a[36] & din_b[40]))))

	.dataa(!din_a[37]),
	.datab(!din_b[39]),
	.datac(!din_a[36]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_121 ),
	.sharein(Xd_0__inst_mult_5_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_128 ),
	.cout(Xd_0__inst_mult_5_129 ),
	.shareout(Xd_0__inst_mult_5_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_38 (
// Equation(s):
// Xd_0__inst_mult_2_124  = SUM(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_2_118  ) + ( Xd_0__inst_mult_2_117  ))
// Xd_0__inst_mult_2_125  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_2_118  ) + ( Xd_0__inst_mult_2_117  ))
// Xd_0__inst_mult_2_126  = SHARE((din_a[19] & (din_b[15] & (din_a[18] & din_b[16]))))

	.dataa(!din_a[19]),
	.datab(!din_b[15]),
	.datac(!din_a[18]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_117 ),
	.sharein(Xd_0__inst_mult_2_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_124 ),
	.cout(Xd_0__inst_mult_2_125 ),
	.shareout(Xd_0__inst_mult_2_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_39 (
// Equation(s):
// Xd_0__inst_mult_2_128  = SUM(( (!din_a[16] & (((din_a[15] & din_b[19])))) # (din_a[16] & (!din_b[18] $ (((!din_a[15]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_122  ) + ( Xd_0__inst_mult_2_121  ))
// Xd_0__inst_mult_2_129  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[19])))) # (din_a[16] & (!din_b[18] $ (((!din_a[15]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_122  ) + ( Xd_0__inst_mult_2_121  ))
// Xd_0__inst_mult_2_130  = SHARE((din_a[16] & (din_b[18] & (din_a[15] & din_b[19]))))

	.dataa(!din_a[16]),
	.datab(!din_b[18]),
	.datac(!din_a[15]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_121 ),
	.sharein(Xd_0__inst_mult_2_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_128 ),
	.cout(Xd_0__inst_mult_2_129 ),
	.shareout(Xd_0__inst_mult_2_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_38 (
// Equation(s):
// Xd_0__inst_mult_3_124  = SUM(( (!din_a[26] & (((din_a[25] & din_b[23])))) # (din_a[26] & (!din_b[22] $ (((!din_a[25]) # (!din_b[23]))))) ) + ( Xd_0__inst_mult_3_118  ) + ( Xd_0__inst_mult_3_117  ))
// Xd_0__inst_mult_3_125  = CARRY(( (!din_a[26] & (((din_a[25] & din_b[23])))) # (din_a[26] & (!din_b[22] $ (((!din_a[25]) # (!din_b[23]))))) ) + ( Xd_0__inst_mult_3_118  ) + ( Xd_0__inst_mult_3_117  ))
// Xd_0__inst_mult_3_126  = SHARE((din_a[26] & (din_b[22] & (din_a[25] & din_b[23]))))

	.dataa(!din_a[26]),
	.datab(!din_b[22]),
	.datac(!din_a[25]),
	.datad(!din_b[23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_117 ),
	.sharein(Xd_0__inst_mult_3_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_124 ),
	.cout(Xd_0__inst_mult_3_125 ),
	.shareout(Xd_0__inst_mult_3_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_39 (
// Equation(s):
// Xd_0__inst_mult_3_128  = SUM(( (!din_a[23] & (((din_a[22] & din_b[26])))) # (din_a[23] & (!din_b[25] $ (((!din_a[22]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_122  ) + ( Xd_0__inst_mult_3_121  ))
// Xd_0__inst_mult_3_129  = CARRY(( (!din_a[23] & (((din_a[22] & din_b[26])))) # (din_a[23] & (!din_b[25] $ (((!din_a[22]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_122  ) + ( Xd_0__inst_mult_3_121  ))
// Xd_0__inst_mult_3_130  = SHARE((din_a[23] & (din_b[25] & (din_a[22] & din_b[26]))))

	.dataa(!din_a[23]),
	.datab(!din_b[25]),
	.datac(!din_a[22]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_121 ),
	.sharein(Xd_0__inst_mult_3_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_128 ),
	.cout(Xd_0__inst_mult_3_129 ),
	.shareout(Xd_0__inst_mult_3_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_38 (
// Equation(s):
// Xd_0__inst_mult_0_124  = SUM(( (!din_a[5] & (((din_a[4] & din_b[2])))) # (din_a[5] & (!din_b[1] $ (((!din_a[4]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_118  ) + ( Xd_0__inst_mult_0_117  ))
// Xd_0__inst_mult_0_125  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[2])))) # (din_a[5] & (!din_b[1] $ (((!din_a[4]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_118  ) + ( Xd_0__inst_mult_0_117  ))
// Xd_0__inst_mult_0_126  = SHARE((din_a[5] & (din_b[1] & (din_a[4] & din_b[2]))))

	.dataa(!din_a[5]),
	.datab(!din_b[1]),
	.datac(!din_a[4]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_117 ),
	.sharein(Xd_0__inst_mult_0_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_124 ),
	.cout(Xd_0__inst_mult_0_125 ),
	.shareout(Xd_0__inst_mult_0_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_39 (
// Equation(s):
// Xd_0__inst_mult_0_128  = SUM(( (!din_a[2] & (((din_a[1] & din_b[5])))) # (din_a[2] & (!din_b[4] $ (((!din_a[1]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_122  ) + ( Xd_0__inst_mult_0_121  ))
// Xd_0__inst_mult_0_129  = CARRY(( (!din_a[2] & (((din_a[1] & din_b[5])))) # (din_a[2] & (!din_b[4] $ (((!din_a[1]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_122  ) + ( Xd_0__inst_mult_0_121  ))
// Xd_0__inst_mult_0_130  = SHARE((din_a[2] & (din_b[4] & (din_a[1] & din_b[5]))))

	.dataa(!din_a[2]),
	.datab(!din_b[4]),
	.datac(!din_a[1]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_121 ),
	.sharein(Xd_0__inst_mult_0_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_128 ),
	.cout(Xd_0__inst_mult_0_129 ),
	.shareout(Xd_0__inst_mult_0_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_38 (
// Equation(s):
// Xd_0__inst_mult_1_124  = SUM(( (!din_a[12] & (((din_a[11] & din_b[9])))) # (din_a[12] & (!din_b[8] $ (((!din_a[11]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_118  ) + ( Xd_0__inst_mult_1_117  ))
// Xd_0__inst_mult_1_125  = CARRY(( (!din_a[12] & (((din_a[11] & din_b[9])))) # (din_a[12] & (!din_b[8] $ (((!din_a[11]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_118  ) + ( Xd_0__inst_mult_1_117  ))
// Xd_0__inst_mult_1_126  = SHARE((din_a[12] & (din_b[8] & (din_a[11] & din_b[9]))))

	.dataa(!din_a[12]),
	.datab(!din_b[8]),
	.datac(!din_a[11]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_117 ),
	.sharein(Xd_0__inst_mult_1_118 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_124 ),
	.cout(Xd_0__inst_mult_1_125 ),
	.shareout(Xd_0__inst_mult_1_126 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_39 (
// Equation(s):
// Xd_0__inst_mult_1_128  = SUM(( (!din_a[9] & (((din_a[8] & din_b[12])))) # (din_a[9] & (!din_b[11] $ (((!din_a[8]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_122  ) + ( Xd_0__inst_mult_1_121  ))
// Xd_0__inst_mult_1_129  = CARRY(( (!din_a[9] & (((din_a[8] & din_b[12])))) # (din_a[9] & (!din_b[11] $ (((!din_a[8]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_122  ) + ( Xd_0__inst_mult_1_121  ))
// Xd_0__inst_mult_1_130  = SHARE((din_a[9] & (din_b[11] & (din_a[8] & din_b[12]))))

	.dataa(!din_a[9]),
	.datab(!din_b[11]),
	.datac(!din_a[8]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_121 ),
	.sharein(Xd_0__inst_mult_1_122 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_128 ),
	.cout(Xd_0__inst_mult_1_129 ),
	.shareout(Xd_0__inst_mult_1_130 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_40 (
// Equation(s):
// Xd_0__inst_mult_28_132  = SUM(( (!din_a[201] & (((din_a[200] & din_b[199])))) # (din_a[201] & (!din_b[198] $ (((!din_a[200]) # (!din_b[199]))))) ) + ( Xd_0__inst_mult_28_126  ) + ( Xd_0__inst_mult_28_125  ))
// Xd_0__inst_mult_28_133  = CARRY(( (!din_a[201] & (((din_a[200] & din_b[199])))) # (din_a[201] & (!din_b[198] $ (((!din_a[200]) # (!din_b[199]))))) ) + ( Xd_0__inst_mult_28_126  ) + ( Xd_0__inst_mult_28_125  ))
// Xd_0__inst_mult_28_134  = SHARE((din_a[201] & (din_b[198] & (din_a[200] & din_b[199]))))

	.dataa(!din_a[201]),
	.datab(!din_b[198]),
	.datac(!din_a[200]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_125 ),
	.sharein(Xd_0__inst_mult_28_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_132 ),
	.cout(Xd_0__inst_mult_28_133 ),
	.shareout(Xd_0__inst_mult_28_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_41 (
// Equation(s):
// Xd_0__inst_mult_28_136  = SUM(( (!din_a[199] & (((din_a[198] & din_b[201])))) # (din_a[199] & (!din_b[200] $ (((!din_a[198]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_130  ) + ( Xd_0__inst_mult_28_129  ))
// Xd_0__inst_mult_28_137  = CARRY(( (!din_a[199] & (((din_a[198] & din_b[201])))) # (din_a[199] & (!din_b[200] $ (((!din_a[198]) # (!din_b[201]))))) ) + ( Xd_0__inst_mult_28_130  ) + ( Xd_0__inst_mult_28_129  ))
// Xd_0__inst_mult_28_138  = SHARE((din_a[199] & (din_b[200] & (din_a[198] & din_b[201]))))

	.dataa(!din_a[199]),
	.datab(!din_b[200]),
	.datac(!din_a[198]),
	.datad(!din_b[201]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_129 ),
	.sharein(Xd_0__inst_mult_28_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_136 ),
	.cout(Xd_0__inst_mult_28_137 ),
	.shareout(Xd_0__inst_mult_28_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_40 (
// Equation(s):
// Xd_0__inst_mult_29_132  = SUM(( (!din_a[208] & (((din_a[207] & din_b[206])))) # (din_a[208] & (!din_b[205] $ (((!din_a[207]) # (!din_b[206]))))) ) + ( Xd_0__inst_mult_29_126  ) + ( Xd_0__inst_mult_29_125  ))
// Xd_0__inst_mult_29_133  = CARRY(( (!din_a[208] & (((din_a[207] & din_b[206])))) # (din_a[208] & (!din_b[205] $ (((!din_a[207]) # (!din_b[206]))))) ) + ( Xd_0__inst_mult_29_126  ) + ( Xd_0__inst_mult_29_125  ))
// Xd_0__inst_mult_29_134  = SHARE((din_a[208] & (din_b[205] & (din_a[207] & din_b[206]))))

	.dataa(!din_a[208]),
	.datab(!din_b[205]),
	.datac(!din_a[207]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_125 ),
	.sharein(Xd_0__inst_mult_29_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_132 ),
	.cout(Xd_0__inst_mult_29_133 ),
	.shareout(Xd_0__inst_mult_29_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_41 (
// Equation(s):
// Xd_0__inst_mult_29_136  = SUM(( (!din_a[206] & (((din_a[205] & din_b[208])))) # (din_a[206] & (!din_b[207] $ (((!din_a[205]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_130  ) + ( Xd_0__inst_mult_29_129  ))
// Xd_0__inst_mult_29_137  = CARRY(( (!din_a[206] & (((din_a[205] & din_b[208])))) # (din_a[206] & (!din_b[207] $ (((!din_a[205]) # (!din_b[208]))))) ) + ( Xd_0__inst_mult_29_130  ) + ( Xd_0__inst_mult_29_129  ))
// Xd_0__inst_mult_29_138  = SHARE((din_a[206] & (din_b[207] & (din_a[205] & din_b[208]))))

	.dataa(!din_a[206]),
	.datab(!din_b[207]),
	.datac(!din_a[205]),
	.datad(!din_b[208]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_129 ),
	.sharein(Xd_0__inst_mult_29_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_136 ),
	.cout(Xd_0__inst_mult_29_137 ),
	.shareout(Xd_0__inst_mult_29_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_40 (
// Equation(s):
// Xd_0__inst_mult_26_132  = SUM(( (!din_a[187] & (((din_a[186] & din_b[185])))) # (din_a[187] & (!din_b[184] $ (((!din_a[186]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_26_126  ) + ( Xd_0__inst_mult_26_125  ))
// Xd_0__inst_mult_26_133  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[185])))) # (din_a[187] & (!din_b[184] $ (((!din_a[186]) # (!din_b[185]))))) ) + ( Xd_0__inst_mult_26_126  ) + ( Xd_0__inst_mult_26_125  ))
// Xd_0__inst_mult_26_134  = SHARE((din_a[187] & (din_b[184] & (din_a[186] & din_b[185]))))

	.dataa(!din_a[187]),
	.datab(!din_b[184]),
	.datac(!din_a[186]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_125 ),
	.sharein(Xd_0__inst_mult_26_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_132 ),
	.cout(Xd_0__inst_mult_26_133 ),
	.shareout(Xd_0__inst_mult_26_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_41 (
// Equation(s):
// Xd_0__inst_mult_26_136  = SUM(( (!din_a[185] & (((din_a[184] & din_b[187])))) # (din_a[185] & (!din_b[186] $ (((!din_a[184]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_130  ) + ( Xd_0__inst_mult_26_129  ))
// Xd_0__inst_mult_26_137  = CARRY(( (!din_a[185] & (((din_a[184] & din_b[187])))) # (din_a[185] & (!din_b[186] $ (((!din_a[184]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_26_130  ) + ( Xd_0__inst_mult_26_129  ))
// Xd_0__inst_mult_26_138  = SHARE((din_a[185] & (din_b[186] & (din_a[184] & din_b[187]))))

	.dataa(!din_a[185]),
	.datab(!din_b[186]),
	.datac(!din_a[184]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_129 ),
	.sharein(Xd_0__inst_mult_26_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_136 ),
	.cout(Xd_0__inst_mult_26_137 ),
	.shareout(Xd_0__inst_mult_26_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_40 (
// Equation(s):
// Xd_0__inst_mult_27_132  = SUM(( (!din_a[194] & (((din_a[193] & din_b[192])))) # (din_a[194] & (!din_b[191] $ (((!din_a[193]) # (!din_b[192]))))) ) + ( Xd_0__inst_mult_27_126  ) + ( Xd_0__inst_mult_27_125  ))
// Xd_0__inst_mult_27_133  = CARRY(( (!din_a[194] & (((din_a[193] & din_b[192])))) # (din_a[194] & (!din_b[191] $ (((!din_a[193]) # (!din_b[192]))))) ) + ( Xd_0__inst_mult_27_126  ) + ( Xd_0__inst_mult_27_125  ))
// Xd_0__inst_mult_27_134  = SHARE((din_a[194] & (din_b[191] & (din_a[193] & din_b[192]))))

	.dataa(!din_a[194]),
	.datab(!din_b[191]),
	.datac(!din_a[193]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_125 ),
	.sharein(Xd_0__inst_mult_27_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_132 ),
	.cout(Xd_0__inst_mult_27_133 ),
	.shareout(Xd_0__inst_mult_27_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_41 (
// Equation(s):
// Xd_0__inst_mult_27_136  = SUM(( (!din_a[192] & (((din_a[191] & din_b[194])))) # (din_a[192] & (!din_b[193] $ (((!din_a[191]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_130  ) + ( Xd_0__inst_mult_27_129  ))
// Xd_0__inst_mult_27_137  = CARRY(( (!din_a[192] & (((din_a[191] & din_b[194])))) # (din_a[192] & (!din_b[193] $ (((!din_a[191]) # (!din_b[194]))))) ) + ( Xd_0__inst_mult_27_130  ) + ( Xd_0__inst_mult_27_129  ))
// Xd_0__inst_mult_27_138  = SHARE((din_a[192] & (din_b[193] & (din_a[191] & din_b[194]))))

	.dataa(!din_a[192]),
	.datab(!din_b[193]),
	.datac(!din_a[191]),
	.datad(!din_b[194]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_129 ),
	.sharein(Xd_0__inst_mult_27_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_136 ),
	.cout(Xd_0__inst_mult_27_137 ),
	.shareout(Xd_0__inst_mult_27_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_40 (
// Equation(s):
// Xd_0__inst_mult_24_132  = SUM(( (!din_a[173] & (((din_a[172] & din_b[171])))) # (din_a[173] & (!din_b[170] $ (((!din_a[172]) # (!din_b[171]))))) ) + ( Xd_0__inst_mult_24_126  ) + ( Xd_0__inst_mult_24_125  ))
// Xd_0__inst_mult_24_133  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[171])))) # (din_a[173] & (!din_b[170] $ (((!din_a[172]) # (!din_b[171]))))) ) + ( Xd_0__inst_mult_24_126  ) + ( Xd_0__inst_mult_24_125  ))
// Xd_0__inst_mult_24_134  = SHARE((din_a[173] & (din_b[170] & (din_a[172] & din_b[171]))))

	.dataa(!din_a[173]),
	.datab(!din_b[170]),
	.datac(!din_a[172]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_125 ),
	.sharein(Xd_0__inst_mult_24_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_132 ),
	.cout(Xd_0__inst_mult_24_133 ),
	.shareout(Xd_0__inst_mult_24_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_41 (
// Equation(s):
// Xd_0__inst_mult_24_136  = SUM(( (!din_a[171] & (((din_a[170] & din_b[173])))) # (din_a[171] & (!din_b[172] $ (((!din_a[170]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_130  ) + ( Xd_0__inst_mult_24_129  ))
// Xd_0__inst_mult_24_137  = CARRY(( (!din_a[171] & (((din_a[170] & din_b[173])))) # (din_a[171] & (!din_b[172] $ (((!din_a[170]) # (!din_b[173]))))) ) + ( Xd_0__inst_mult_24_130  ) + ( Xd_0__inst_mult_24_129  ))
// Xd_0__inst_mult_24_138  = SHARE((din_a[171] & (din_b[172] & (din_a[170] & din_b[173]))))

	.dataa(!din_a[171]),
	.datab(!din_b[172]),
	.datac(!din_a[170]),
	.datad(!din_b[173]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_129 ),
	.sharein(Xd_0__inst_mult_24_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_136 ),
	.cout(Xd_0__inst_mult_24_137 ),
	.shareout(Xd_0__inst_mult_24_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_41 (
// Equation(s):
// Xd_0__inst_mult_25_136  = SUM(( (!din_a[180] & (((din_a[179] & din_b[178])))) # (din_a[180] & (!din_b[177] $ (((!din_a[179]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_25_130  ) + ( Xd_0__inst_mult_25_129  ))
// Xd_0__inst_mult_25_137  = CARRY(( (!din_a[180] & (((din_a[179] & din_b[178])))) # (din_a[180] & (!din_b[177] $ (((!din_a[179]) # (!din_b[178]))))) ) + ( Xd_0__inst_mult_25_130  ) + ( Xd_0__inst_mult_25_129  ))
// Xd_0__inst_mult_25_138  = SHARE((din_a[180] & (din_b[177] & (din_a[179] & din_b[178]))))

	.dataa(!din_a[180]),
	.datab(!din_b[177]),
	.datac(!din_a[179]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_129 ),
	.sharein(Xd_0__inst_mult_25_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_136 ),
	.cout(Xd_0__inst_mult_25_137 ),
	.shareout(Xd_0__inst_mult_25_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_42 (
// Equation(s):
// Xd_0__inst_mult_25_140  = SUM(( (!din_a[178] & (((din_a[177] & din_b[180])))) # (din_a[178] & (!din_b[179] $ (((!din_a[177]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_134  ) + ( Xd_0__inst_mult_25_133  ))
// Xd_0__inst_mult_25_141  = CARRY(( (!din_a[178] & (((din_a[177] & din_b[180])))) # (din_a[178] & (!din_b[179] $ (((!din_a[177]) # (!din_b[180]))))) ) + ( Xd_0__inst_mult_25_134  ) + ( Xd_0__inst_mult_25_133  ))
// Xd_0__inst_mult_25_142  = SHARE((din_a[178] & (din_b[179] & (din_a[177] & din_b[180]))))

	.dataa(!din_a[178]),
	.datab(!din_b[179]),
	.datac(!din_a[177]),
	.datad(!din_b[180]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_133 ),
	.sharein(Xd_0__inst_mult_25_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_140 ),
	.cout(Xd_0__inst_mult_25_141 ),
	.shareout(Xd_0__inst_mult_25_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_41 (
// Equation(s):
// Xd_0__inst_mult_22_136  = SUM(( (!din_a[159] & (((din_a[158] & din_b[157])))) # (din_a[159] & (!din_b[156] $ (((!din_a[158]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_22_130  ) + ( Xd_0__inst_mult_22_129  ))
// Xd_0__inst_mult_22_137  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[157])))) # (din_a[159] & (!din_b[156] $ (((!din_a[158]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_22_130  ) + ( Xd_0__inst_mult_22_129  ))
// Xd_0__inst_mult_22_138  = SHARE((din_a[159] & (din_b[156] & (din_a[158] & din_b[157]))))

	.dataa(!din_a[159]),
	.datab(!din_b[156]),
	.datac(!din_a[158]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_129 ),
	.sharein(Xd_0__inst_mult_22_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_136 ),
	.cout(Xd_0__inst_mult_22_137 ),
	.shareout(Xd_0__inst_mult_22_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_42 (
// Equation(s):
// Xd_0__inst_mult_22_140  = SUM(( (!din_a[157] & (((din_a[156] & din_b[159])))) # (din_a[157] & (!din_b[158] $ (((!din_a[156]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_134  ) + ( Xd_0__inst_mult_22_133  ))
// Xd_0__inst_mult_22_141  = CARRY(( (!din_a[157] & (((din_a[156] & din_b[159])))) # (din_a[157] & (!din_b[158] $ (((!din_a[156]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_22_134  ) + ( Xd_0__inst_mult_22_133  ))
// Xd_0__inst_mult_22_142  = SHARE((din_a[157] & (din_b[158] & (din_a[156] & din_b[159]))))

	.dataa(!din_a[157]),
	.datab(!din_b[158]),
	.datac(!din_a[156]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_133 ),
	.sharein(Xd_0__inst_mult_22_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_140 ),
	.cout(Xd_0__inst_mult_22_141 ),
	.shareout(Xd_0__inst_mult_22_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_40 (
// Equation(s):
// Xd_0__inst_mult_23_132  = SUM(( (!din_a[166] & (((din_a[165] & din_b[164])))) # (din_a[166] & (!din_b[163] $ (((!din_a[165]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_23_126  ) + ( Xd_0__inst_mult_23_125  ))
// Xd_0__inst_mult_23_133  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[164])))) # (din_a[166] & (!din_b[163] $ (((!din_a[165]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_23_126  ) + ( Xd_0__inst_mult_23_125  ))
// Xd_0__inst_mult_23_134  = SHARE((din_a[166] & (din_b[163] & (din_a[165] & din_b[164]))))

	.dataa(!din_a[166]),
	.datab(!din_b[163]),
	.datac(!din_a[165]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_125 ),
	.sharein(Xd_0__inst_mult_23_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_132 ),
	.cout(Xd_0__inst_mult_23_133 ),
	.shareout(Xd_0__inst_mult_23_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_41 (
// Equation(s):
// Xd_0__inst_mult_23_136  = SUM(( (!din_a[164] & (((din_a[163] & din_b[166])))) # (din_a[164] & (!din_b[165] $ (((!din_a[163]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_130  ) + ( Xd_0__inst_mult_23_129  ))
// Xd_0__inst_mult_23_137  = CARRY(( (!din_a[164] & (((din_a[163] & din_b[166])))) # (din_a[164] & (!din_b[165] $ (((!din_a[163]) # (!din_b[166]))))) ) + ( Xd_0__inst_mult_23_130  ) + ( Xd_0__inst_mult_23_129  ))
// Xd_0__inst_mult_23_138  = SHARE((din_a[164] & (din_b[165] & (din_a[163] & din_b[166]))))

	.dataa(!din_a[164]),
	.datab(!din_b[165]),
	.datac(!din_a[163]),
	.datad(!din_b[166]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_129 ),
	.sharein(Xd_0__inst_mult_23_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_136 ),
	.cout(Xd_0__inst_mult_23_137 ),
	.shareout(Xd_0__inst_mult_23_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_40 (
// Equation(s):
// Xd_0__inst_mult_20_132  = SUM(( (!din_a[145] & (((din_a[144] & din_b[143])))) # (din_a[145] & (!din_b[142] $ (((!din_a[144]) # (!din_b[143]))))) ) + ( Xd_0__inst_mult_20_126  ) + ( Xd_0__inst_mult_20_125  ))
// Xd_0__inst_mult_20_133  = CARRY(( (!din_a[145] & (((din_a[144] & din_b[143])))) # (din_a[145] & (!din_b[142] $ (((!din_a[144]) # (!din_b[143]))))) ) + ( Xd_0__inst_mult_20_126  ) + ( Xd_0__inst_mult_20_125  ))
// Xd_0__inst_mult_20_134  = SHARE((din_a[145] & (din_b[142] & (din_a[144] & din_b[143]))))

	.dataa(!din_a[145]),
	.datab(!din_b[142]),
	.datac(!din_a[144]),
	.datad(!din_b[143]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_125 ),
	.sharein(Xd_0__inst_mult_20_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_132 ),
	.cout(Xd_0__inst_mult_20_133 ),
	.shareout(Xd_0__inst_mult_20_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_41 (
// Equation(s):
// Xd_0__inst_mult_20_136  = SUM(( (!din_a[143] & (((din_a[142] & din_b[145])))) # (din_a[143] & (!din_b[144] $ (((!din_a[142]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_130  ) + ( Xd_0__inst_mult_20_129  ))
// Xd_0__inst_mult_20_137  = CARRY(( (!din_a[143] & (((din_a[142] & din_b[145])))) # (din_a[143] & (!din_b[144] $ (((!din_a[142]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_20_130  ) + ( Xd_0__inst_mult_20_129  ))
// Xd_0__inst_mult_20_138  = SHARE((din_a[143] & (din_b[144] & (din_a[142] & din_b[145]))))

	.dataa(!din_a[143]),
	.datab(!din_b[144]),
	.datac(!din_a[142]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_129 ),
	.sharein(Xd_0__inst_mult_20_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_136 ),
	.cout(Xd_0__inst_mult_20_137 ),
	.shareout(Xd_0__inst_mult_20_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_40 (
// Equation(s):
// Xd_0__inst_mult_21_132  = SUM(( (!din_a[152] & (((din_a[151] & din_b[150])))) # (din_a[152] & (!din_b[149] $ (((!din_a[151]) # (!din_b[150]))))) ) + ( Xd_0__inst_mult_21_126  ) + ( Xd_0__inst_mult_21_125  ))
// Xd_0__inst_mult_21_133  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[150])))) # (din_a[152] & (!din_b[149] $ (((!din_a[151]) # (!din_b[150]))))) ) + ( Xd_0__inst_mult_21_126  ) + ( Xd_0__inst_mult_21_125  ))
// Xd_0__inst_mult_21_134  = SHARE((din_a[152] & (din_b[149] & (din_a[151] & din_b[150]))))

	.dataa(!din_a[152]),
	.datab(!din_b[149]),
	.datac(!din_a[151]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_125 ),
	.sharein(Xd_0__inst_mult_21_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_132 ),
	.cout(Xd_0__inst_mult_21_133 ),
	.shareout(Xd_0__inst_mult_21_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_41 (
// Equation(s):
// Xd_0__inst_mult_21_136  = SUM(( (!din_a[150] & (((din_a[149] & din_b[152])))) # (din_a[150] & (!din_b[151] $ (((!din_a[149]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_130  ) + ( Xd_0__inst_mult_21_129  ))
// Xd_0__inst_mult_21_137  = CARRY(( (!din_a[150] & (((din_a[149] & din_b[152])))) # (din_a[150] & (!din_b[151] $ (((!din_a[149]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_21_130  ) + ( Xd_0__inst_mult_21_129  ))
// Xd_0__inst_mult_21_138  = SHARE((din_a[150] & (din_b[151] & (din_a[149] & din_b[152]))))

	.dataa(!din_a[150]),
	.datab(!din_b[151]),
	.datac(!din_a[149]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_129 ),
	.sharein(Xd_0__inst_mult_21_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_136 ),
	.cout(Xd_0__inst_mult_21_137 ),
	.shareout(Xd_0__inst_mult_21_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_40 (
// Equation(s):
// Xd_0__inst_mult_18_132  = SUM(( (!din_a[131] & (((din_a[130] & din_b[129])))) # (din_a[131] & (!din_b[128] $ (((!din_a[130]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_18_126  ) + ( Xd_0__inst_mult_18_125  ))
// Xd_0__inst_mult_18_133  = CARRY(( (!din_a[131] & (((din_a[130] & din_b[129])))) # (din_a[131] & (!din_b[128] $ (((!din_a[130]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_18_126  ) + ( Xd_0__inst_mult_18_125  ))
// Xd_0__inst_mult_18_134  = SHARE((din_a[131] & (din_b[128] & (din_a[130] & din_b[129]))))

	.dataa(!din_a[131]),
	.datab(!din_b[128]),
	.datac(!din_a[130]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_125 ),
	.sharein(Xd_0__inst_mult_18_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_132 ),
	.cout(Xd_0__inst_mult_18_133 ),
	.shareout(Xd_0__inst_mult_18_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_41 (
// Equation(s):
// Xd_0__inst_mult_18_136  = SUM(( (!din_a[129] & (((din_a[128] & din_b[131])))) # (din_a[129] & (!din_b[130] $ (((!din_a[128]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_130  ) + ( Xd_0__inst_mult_18_129  ))
// Xd_0__inst_mult_18_137  = CARRY(( (!din_a[129] & (((din_a[128] & din_b[131])))) # (din_a[129] & (!din_b[130] $ (((!din_a[128]) # (!din_b[131]))))) ) + ( Xd_0__inst_mult_18_130  ) + ( Xd_0__inst_mult_18_129  ))
// Xd_0__inst_mult_18_138  = SHARE((din_a[129] & (din_b[130] & (din_a[128] & din_b[131]))))

	.dataa(!din_a[129]),
	.datab(!din_b[130]),
	.datac(!din_a[128]),
	.datad(!din_b[131]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_129 ),
	.sharein(Xd_0__inst_mult_18_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_136 ),
	.cout(Xd_0__inst_mult_18_137 ),
	.shareout(Xd_0__inst_mult_18_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_40 (
// Equation(s):
// Xd_0__inst_mult_19_132  = SUM(( (!din_a[138] & (((din_a[137] & din_b[136])))) # (din_a[138] & (!din_b[135] $ (((!din_a[137]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_19_126  ) + ( Xd_0__inst_mult_19_125  ))
// Xd_0__inst_mult_19_133  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[136])))) # (din_a[138] & (!din_b[135] $ (((!din_a[137]) # (!din_b[136]))))) ) + ( Xd_0__inst_mult_19_126  ) + ( Xd_0__inst_mult_19_125  ))
// Xd_0__inst_mult_19_134  = SHARE((din_a[138] & (din_b[135] & (din_a[137] & din_b[136]))))

	.dataa(!din_a[138]),
	.datab(!din_b[135]),
	.datac(!din_a[137]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_125 ),
	.sharein(Xd_0__inst_mult_19_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_132 ),
	.cout(Xd_0__inst_mult_19_133 ),
	.shareout(Xd_0__inst_mult_19_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_41 (
// Equation(s):
// Xd_0__inst_mult_19_136  = SUM(( (!din_a[136] & (((din_a[135] & din_b[138])))) # (din_a[136] & (!din_b[137] $ (((!din_a[135]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_130  ) + ( Xd_0__inst_mult_19_129  ))
// Xd_0__inst_mult_19_137  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[138])))) # (din_a[136] & (!din_b[137] $ (((!din_a[135]) # (!din_b[138]))))) ) + ( Xd_0__inst_mult_19_130  ) + ( Xd_0__inst_mult_19_129  ))
// Xd_0__inst_mult_19_138  = SHARE((din_a[136] & (din_b[137] & (din_a[135] & din_b[138]))))

	.dataa(!din_a[136]),
	.datab(!din_b[137]),
	.datac(!din_a[135]),
	.datad(!din_b[138]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_129 ),
	.sharein(Xd_0__inst_mult_19_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_136 ),
	.cout(Xd_0__inst_mult_19_137 ),
	.shareout(Xd_0__inst_mult_19_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_40 (
// Equation(s):
// Xd_0__inst_mult_16_132  = SUM(( (!din_a[117] & (((din_a[116] & din_b[115])))) # (din_a[117] & (!din_b[114] $ (((!din_a[116]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_16_126  ) + ( Xd_0__inst_mult_16_125  ))
// Xd_0__inst_mult_16_133  = CARRY(( (!din_a[117] & (((din_a[116] & din_b[115])))) # (din_a[117] & (!din_b[114] $ (((!din_a[116]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_16_126  ) + ( Xd_0__inst_mult_16_125  ))
// Xd_0__inst_mult_16_134  = SHARE((din_a[117] & (din_b[114] & (din_a[116] & din_b[115]))))

	.dataa(!din_a[117]),
	.datab(!din_b[114]),
	.datac(!din_a[116]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_125 ),
	.sharein(Xd_0__inst_mult_16_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_132 ),
	.cout(Xd_0__inst_mult_16_133 ),
	.shareout(Xd_0__inst_mult_16_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_41 (
// Equation(s):
// Xd_0__inst_mult_16_136  = SUM(( (!din_a[115] & (((din_a[114] & din_b[117])))) # (din_a[115] & (!din_b[116] $ (((!din_a[114]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_130  ) + ( Xd_0__inst_mult_16_129  ))
// Xd_0__inst_mult_16_137  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[117])))) # (din_a[115] & (!din_b[116] $ (((!din_a[114]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_16_130  ) + ( Xd_0__inst_mult_16_129  ))
// Xd_0__inst_mult_16_138  = SHARE((din_a[115] & (din_b[116] & (din_a[114] & din_b[117]))))

	.dataa(!din_a[115]),
	.datab(!din_b[116]),
	.datac(!din_a[114]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_129 ),
	.sharein(Xd_0__inst_mult_16_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_136 ),
	.cout(Xd_0__inst_mult_16_137 ),
	.shareout(Xd_0__inst_mult_16_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_40 (
// Equation(s):
// Xd_0__inst_mult_17_132  = SUM(( (!din_a[124] & (((din_a[123] & din_b[122])))) # (din_a[124] & (!din_b[121] $ (((!din_a[123]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_17_126  ) + ( Xd_0__inst_mult_17_125  ))
// Xd_0__inst_mult_17_133  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[122])))) # (din_a[124] & (!din_b[121] $ (((!din_a[123]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_17_126  ) + ( Xd_0__inst_mult_17_125  ))
// Xd_0__inst_mult_17_134  = SHARE((din_a[124] & (din_b[121] & (din_a[123] & din_b[122]))))

	.dataa(!din_a[124]),
	.datab(!din_b[121]),
	.datac(!din_a[123]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_125 ),
	.sharein(Xd_0__inst_mult_17_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_132 ),
	.cout(Xd_0__inst_mult_17_133 ),
	.shareout(Xd_0__inst_mult_17_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_41 (
// Equation(s):
// Xd_0__inst_mult_17_136  = SUM(( (!din_a[122] & (((din_a[121] & din_b[124])))) # (din_a[122] & (!din_b[123] $ (((!din_a[121]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_130  ) + ( Xd_0__inst_mult_17_129  ))
// Xd_0__inst_mult_17_137  = CARRY(( (!din_a[122] & (((din_a[121] & din_b[124])))) # (din_a[122] & (!din_b[123] $ (((!din_a[121]) # (!din_b[124]))))) ) + ( Xd_0__inst_mult_17_130  ) + ( Xd_0__inst_mult_17_129  ))
// Xd_0__inst_mult_17_138  = SHARE((din_a[122] & (din_b[123] & (din_a[121] & din_b[124]))))

	.dataa(!din_a[122]),
	.datab(!din_b[123]),
	.datac(!din_a[121]),
	.datad(!din_b[124]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_129 ),
	.sharein(Xd_0__inst_mult_17_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_136 ),
	.cout(Xd_0__inst_mult_17_137 ),
	.shareout(Xd_0__inst_mult_17_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_40 (
// Equation(s):
// Xd_0__inst_mult_14_132  = SUM(( (!din_a[103] & (((din_a[102] & din_b[101])))) # (din_a[103] & (!din_b[100] $ (((!din_a[102]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_14_126  ) + ( Xd_0__inst_mult_14_125  ))
// Xd_0__inst_mult_14_133  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[101])))) # (din_a[103] & (!din_b[100] $ (((!din_a[102]) # (!din_b[101]))))) ) + ( Xd_0__inst_mult_14_126  ) + ( Xd_0__inst_mult_14_125  ))
// Xd_0__inst_mult_14_134  = SHARE((din_a[103] & (din_b[100] & (din_a[102] & din_b[101]))))

	.dataa(!din_a[103]),
	.datab(!din_b[100]),
	.datac(!din_a[102]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_125 ),
	.sharein(Xd_0__inst_mult_14_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_132 ),
	.cout(Xd_0__inst_mult_14_133 ),
	.shareout(Xd_0__inst_mult_14_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_41 (
// Equation(s):
// Xd_0__inst_mult_14_136  = SUM(( (!din_a[101] & (((din_a[100] & din_b[103])))) # (din_a[101] & (!din_b[102] $ (((!din_a[100]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_130  ) + ( Xd_0__inst_mult_14_129  ))
// Xd_0__inst_mult_14_137  = CARRY(( (!din_a[101] & (((din_a[100] & din_b[103])))) # (din_a[101] & (!din_b[102] $ (((!din_a[100]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_14_130  ) + ( Xd_0__inst_mult_14_129  ))
// Xd_0__inst_mult_14_138  = SHARE((din_a[101] & (din_b[102] & (din_a[100] & din_b[103]))))

	.dataa(!din_a[101]),
	.datab(!din_b[102]),
	.datac(!din_a[100]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_129 ),
	.sharein(Xd_0__inst_mult_14_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_136 ),
	.cout(Xd_0__inst_mult_14_137 ),
	.shareout(Xd_0__inst_mult_14_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_40 (
// Equation(s):
// Xd_0__inst_mult_15_132  = SUM(( (!din_a[110] & (((din_a[109] & din_b[108])))) # (din_a[110] & (!din_b[107] $ (((!din_a[109]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_15_126  ) + ( Xd_0__inst_mult_15_125  ))
// Xd_0__inst_mult_15_133  = CARRY(( (!din_a[110] & (((din_a[109] & din_b[108])))) # (din_a[110] & (!din_b[107] $ (((!din_a[109]) # (!din_b[108]))))) ) + ( Xd_0__inst_mult_15_126  ) + ( Xd_0__inst_mult_15_125  ))
// Xd_0__inst_mult_15_134  = SHARE((din_a[110] & (din_b[107] & (din_a[109] & din_b[108]))))

	.dataa(!din_a[110]),
	.datab(!din_b[107]),
	.datac(!din_a[109]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_125 ),
	.sharein(Xd_0__inst_mult_15_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_132 ),
	.cout(Xd_0__inst_mult_15_133 ),
	.shareout(Xd_0__inst_mult_15_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_41 (
// Equation(s):
// Xd_0__inst_mult_15_136  = SUM(( (!din_a[108] & (((din_a[107] & din_b[110])))) # (din_a[108] & (!din_b[109] $ (((!din_a[107]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_130  ) + ( Xd_0__inst_mult_15_129  ))
// Xd_0__inst_mult_15_137  = CARRY(( (!din_a[108] & (((din_a[107] & din_b[110])))) # (din_a[108] & (!din_b[109] $ (((!din_a[107]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_15_130  ) + ( Xd_0__inst_mult_15_129  ))
// Xd_0__inst_mult_15_138  = SHARE((din_a[108] & (din_b[109] & (din_a[107] & din_b[110]))))

	.dataa(!din_a[108]),
	.datab(!din_b[109]),
	.datac(!din_a[107]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_129 ),
	.sharein(Xd_0__inst_mult_15_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_136 ),
	.cout(Xd_0__inst_mult_15_137 ),
	.shareout(Xd_0__inst_mult_15_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_40 (
// Equation(s):
// Xd_0__inst_mult_12_132  = SUM(( (!din_a[89] & (((din_a[88] & din_b[87])))) # (din_a[89] & (!din_b[86] $ (((!din_a[88]) # (!din_b[87]))))) ) + ( Xd_0__inst_mult_12_126  ) + ( Xd_0__inst_mult_12_125  ))
// Xd_0__inst_mult_12_133  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[87])))) # (din_a[89] & (!din_b[86] $ (((!din_a[88]) # (!din_b[87]))))) ) + ( Xd_0__inst_mult_12_126  ) + ( Xd_0__inst_mult_12_125  ))
// Xd_0__inst_mult_12_134  = SHARE((din_a[89] & (din_b[86] & (din_a[88] & din_b[87]))))

	.dataa(!din_a[89]),
	.datab(!din_b[86]),
	.datac(!din_a[88]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_125 ),
	.sharein(Xd_0__inst_mult_12_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_132 ),
	.cout(Xd_0__inst_mult_12_133 ),
	.shareout(Xd_0__inst_mult_12_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_41 (
// Equation(s):
// Xd_0__inst_mult_12_136  = SUM(( (!din_a[87] & (((din_a[86] & din_b[89])))) # (din_a[87] & (!din_b[88] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_130  ) + ( Xd_0__inst_mult_12_129  ))
// Xd_0__inst_mult_12_137  = CARRY(( (!din_a[87] & (((din_a[86] & din_b[89])))) # (din_a[87] & (!din_b[88] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_12_130  ) + ( Xd_0__inst_mult_12_129  ))
// Xd_0__inst_mult_12_138  = SHARE((din_a[87] & (din_b[88] & (din_a[86] & din_b[89]))))

	.dataa(!din_a[87]),
	.datab(!din_b[88]),
	.datac(!din_a[86]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_129 ),
	.sharein(Xd_0__inst_mult_12_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_136 ),
	.cout(Xd_0__inst_mult_12_137 ),
	.shareout(Xd_0__inst_mult_12_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_40 (
// Equation(s):
// Xd_0__inst_mult_13_132  = SUM(( (!din_a[96] & (((din_a[95] & din_b[94])))) # (din_a[96] & (!din_b[93] $ (((!din_a[95]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_13_126  ) + ( Xd_0__inst_mult_13_125  ))
// Xd_0__inst_mult_13_133  = CARRY(( (!din_a[96] & (((din_a[95] & din_b[94])))) # (din_a[96] & (!din_b[93] $ (((!din_a[95]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_13_126  ) + ( Xd_0__inst_mult_13_125  ))
// Xd_0__inst_mult_13_134  = SHARE((din_a[96] & (din_b[93] & (din_a[95] & din_b[94]))))

	.dataa(!din_a[96]),
	.datab(!din_b[93]),
	.datac(!din_a[95]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_125 ),
	.sharein(Xd_0__inst_mult_13_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_132 ),
	.cout(Xd_0__inst_mult_13_133 ),
	.shareout(Xd_0__inst_mult_13_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_41 (
// Equation(s):
// Xd_0__inst_mult_13_136  = SUM(( (!din_a[94] & (((din_a[93] & din_b[96])))) # (din_a[94] & (!din_b[95] $ (((!din_a[93]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_130  ) + ( Xd_0__inst_mult_13_129  ))
// Xd_0__inst_mult_13_137  = CARRY(( (!din_a[94] & (((din_a[93] & din_b[96])))) # (din_a[94] & (!din_b[95] $ (((!din_a[93]) # (!din_b[96]))))) ) + ( Xd_0__inst_mult_13_130  ) + ( Xd_0__inst_mult_13_129  ))
// Xd_0__inst_mult_13_138  = SHARE((din_a[94] & (din_b[95] & (din_a[93] & din_b[96]))))

	.dataa(!din_a[94]),
	.datab(!din_b[95]),
	.datac(!din_a[93]),
	.datad(!din_b[96]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_129 ),
	.sharein(Xd_0__inst_mult_13_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_136 ),
	.cout(Xd_0__inst_mult_13_137 ),
	.shareout(Xd_0__inst_mult_13_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_40 (
// Equation(s):
// Xd_0__inst_mult_10_132  = SUM(( (!din_a[75] & (((din_a[74] & din_b[73])))) # (din_a[75] & (!din_b[72] $ (((!din_a[74]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_10_126  ) + ( Xd_0__inst_mult_10_125  ))
// Xd_0__inst_mult_10_133  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[73])))) # (din_a[75] & (!din_b[72] $ (((!din_a[74]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_10_126  ) + ( Xd_0__inst_mult_10_125  ))
// Xd_0__inst_mult_10_134  = SHARE((din_a[75] & (din_b[72] & (din_a[74] & din_b[73]))))

	.dataa(!din_a[75]),
	.datab(!din_b[72]),
	.datac(!din_a[74]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_125 ),
	.sharein(Xd_0__inst_mult_10_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_132 ),
	.cout(Xd_0__inst_mult_10_133 ),
	.shareout(Xd_0__inst_mult_10_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_41 (
// Equation(s):
// Xd_0__inst_mult_10_136  = SUM(( (!din_a[73] & (((din_a[72] & din_b[75])))) # (din_a[73] & (!din_b[74] $ (((!din_a[72]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_130  ) + ( Xd_0__inst_mult_10_129  ))
// Xd_0__inst_mult_10_137  = CARRY(( (!din_a[73] & (((din_a[72] & din_b[75])))) # (din_a[73] & (!din_b[74] $ (((!din_a[72]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_10_130  ) + ( Xd_0__inst_mult_10_129  ))
// Xd_0__inst_mult_10_138  = SHARE((din_a[73] & (din_b[74] & (din_a[72] & din_b[75]))))

	.dataa(!din_a[73]),
	.datab(!din_b[74]),
	.datac(!din_a[72]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_129 ),
	.sharein(Xd_0__inst_mult_10_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_136 ),
	.cout(Xd_0__inst_mult_10_137 ),
	.shareout(Xd_0__inst_mult_10_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_40 (
// Equation(s):
// Xd_0__inst_mult_11_132  = SUM(( (!din_a[82] & (((din_a[81] & din_b[80])))) # (din_a[82] & (!din_b[79] $ (((!din_a[81]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_11_126  ) + ( Xd_0__inst_mult_11_125  ))
// Xd_0__inst_mult_11_133  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[80])))) # (din_a[82] & (!din_b[79] $ (((!din_a[81]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_11_126  ) + ( Xd_0__inst_mult_11_125  ))
// Xd_0__inst_mult_11_134  = SHARE((din_a[82] & (din_b[79] & (din_a[81] & din_b[80]))))

	.dataa(!din_a[82]),
	.datab(!din_b[79]),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_125 ),
	.sharein(Xd_0__inst_mult_11_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_132 ),
	.cout(Xd_0__inst_mult_11_133 ),
	.shareout(Xd_0__inst_mult_11_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_41 (
// Equation(s):
// Xd_0__inst_mult_11_136  = SUM(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_130  ) + ( Xd_0__inst_mult_11_129  ))
// Xd_0__inst_mult_11_137  = CARRY(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_11_130  ) + ( Xd_0__inst_mult_11_129  ))
// Xd_0__inst_mult_11_138  = SHARE((din_a[80] & (din_b[81] & (din_a[79] & din_b[82]))))

	.dataa(!din_a[80]),
	.datab(!din_b[81]),
	.datac(!din_a[79]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_129 ),
	.sharein(Xd_0__inst_mult_11_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_136 ),
	.cout(Xd_0__inst_mult_11_137 ),
	.shareout(Xd_0__inst_mult_11_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_40 (
// Equation(s):
// Xd_0__inst_mult_8_132  = SUM(( (!din_a[61] & (((din_a[60] & din_b[59])))) # (din_a[61] & (!din_b[58] $ (((!din_a[60]) # (!din_b[59]))))) ) + ( Xd_0__inst_mult_8_126  ) + ( Xd_0__inst_mult_8_125  ))
// Xd_0__inst_mult_8_133  = CARRY(( (!din_a[61] & (((din_a[60] & din_b[59])))) # (din_a[61] & (!din_b[58] $ (((!din_a[60]) # (!din_b[59]))))) ) + ( Xd_0__inst_mult_8_126  ) + ( Xd_0__inst_mult_8_125  ))
// Xd_0__inst_mult_8_134  = SHARE((din_a[61] & (din_b[58] & (din_a[60] & din_b[59]))))

	.dataa(!din_a[61]),
	.datab(!din_b[58]),
	.datac(!din_a[60]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_125 ),
	.sharein(Xd_0__inst_mult_8_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_132 ),
	.cout(Xd_0__inst_mult_8_133 ),
	.shareout(Xd_0__inst_mult_8_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_41 (
// Equation(s):
// Xd_0__inst_mult_8_136  = SUM(( (!din_a[59] & (((din_a[58] & din_b[61])))) # (din_a[59] & (!din_b[60] $ (((!din_a[58]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_130  ) + ( Xd_0__inst_mult_8_129  ))
// Xd_0__inst_mult_8_137  = CARRY(( (!din_a[59] & (((din_a[58] & din_b[61])))) # (din_a[59] & (!din_b[60] $ (((!din_a[58]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_8_130  ) + ( Xd_0__inst_mult_8_129  ))
// Xd_0__inst_mult_8_138  = SHARE((din_a[59] & (din_b[60] & (din_a[58] & din_b[61]))))

	.dataa(!din_a[59]),
	.datab(!din_b[60]),
	.datac(!din_a[58]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_129 ),
	.sharein(Xd_0__inst_mult_8_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_136 ),
	.cout(Xd_0__inst_mult_8_137 ),
	.shareout(Xd_0__inst_mult_8_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_40 (
// Equation(s):
// Xd_0__inst_mult_9_132  = SUM(( (!din_a[68] & (((din_a[67] & din_b[66])))) # (din_a[68] & (!din_b[65] $ (((!din_a[67]) # (!din_b[66]))))) ) + ( Xd_0__inst_mult_9_126  ) + ( Xd_0__inst_mult_9_125  ))
// Xd_0__inst_mult_9_133  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[66])))) # (din_a[68] & (!din_b[65] $ (((!din_a[67]) # (!din_b[66]))))) ) + ( Xd_0__inst_mult_9_126  ) + ( Xd_0__inst_mult_9_125  ))
// Xd_0__inst_mult_9_134  = SHARE((din_a[68] & (din_b[65] & (din_a[67] & din_b[66]))))

	.dataa(!din_a[68]),
	.datab(!din_b[65]),
	.datac(!din_a[67]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_125 ),
	.sharein(Xd_0__inst_mult_9_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_132 ),
	.cout(Xd_0__inst_mult_9_133 ),
	.shareout(Xd_0__inst_mult_9_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_41 (
// Equation(s):
// Xd_0__inst_mult_9_136  = SUM(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_130  ) + ( Xd_0__inst_mult_9_129  ))
// Xd_0__inst_mult_9_137  = CARRY(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_9_130  ) + ( Xd_0__inst_mult_9_129  ))
// Xd_0__inst_mult_9_138  = SHARE((din_a[66] & (din_b[67] & (din_a[65] & din_b[68]))))

	.dataa(!din_a[66]),
	.datab(!din_b[67]),
	.datac(!din_a[65]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_129 ),
	.sharein(Xd_0__inst_mult_9_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_136 ),
	.cout(Xd_0__inst_mult_9_137 ),
	.shareout(Xd_0__inst_mult_9_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_40 (
// Equation(s):
// Xd_0__inst_mult_6_132  = SUM(( (!din_a[47] & (((din_a[46] & din_b[45])))) # (din_a[47] & (!din_b[44] $ (((!din_a[46]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_6_126  ) + ( Xd_0__inst_mult_6_125  ))
// Xd_0__inst_mult_6_133  = CARRY(( (!din_a[47] & (((din_a[46] & din_b[45])))) # (din_a[47] & (!din_b[44] $ (((!din_a[46]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_6_126  ) + ( Xd_0__inst_mult_6_125  ))
// Xd_0__inst_mult_6_134  = SHARE((din_a[47] & (din_b[44] & (din_a[46] & din_b[45]))))

	.dataa(!din_a[47]),
	.datab(!din_b[44]),
	.datac(!din_a[46]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_125 ),
	.sharein(Xd_0__inst_mult_6_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_132 ),
	.cout(Xd_0__inst_mult_6_133 ),
	.shareout(Xd_0__inst_mult_6_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_41 (
// Equation(s):
// Xd_0__inst_mult_6_136  = SUM(( (!din_a[45] & (((din_a[44] & din_b[47])))) # (din_a[45] & (!din_b[46] $ (((!din_a[44]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_130  ) + ( Xd_0__inst_mult_6_129  ))
// Xd_0__inst_mult_6_137  = CARRY(( (!din_a[45] & (((din_a[44] & din_b[47])))) # (din_a[45] & (!din_b[46] $ (((!din_a[44]) # (!din_b[47]))))) ) + ( Xd_0__inst_mult_6_130  ) + ( Xd_0__inst_mult_6_129  ))
// Xd_0__inst_mult_6_138  = SHARE((din_a[45] & (din_b[46] & (din_a[44] & din_b[47]))))

	.dataa(!din_a[45]),
	.datab(!din_b[46]),
	.datac(!din_a[44]),
	.datad(!din_b[47]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_129 ),
	.sharein(Xd_0__inst_mult_6_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_136 ),
	.cout(Xd_0__inst_mult_6_137 ),
	.shareout(Xd_0__inst_mult_6_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_40 (
// Equation(s):
// Xd_0__inst_mult_7_132  = SUM(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_7_126  ) + ( Xd_0__inst_mult_7_125  ))
// Xd_0__inst_mult_7_133  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_7_126  ) + ( Xd_0__inst_mult_7_125  ))
// Xd_0__inst_mult_7_134  = SHARE((din_a[54] & (din_b[51] & (din_a[53] & din_b[52]))))

	.dataa(!din_a[54]),
	.datab(!din_b[51]),
	.datac(!din_a[53]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_125 ),
	.sharein(Xd_0__inst_mult_7_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_132 ),
	.cout(Xd_0__inst_mult_7_133 ),
	.shareout(Xd_0__inst_mult_7_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_41 (
// Equation(s):
// Xd_0__inst_mult_7_136  = SUM(( (!din_a[52] & (((din_a[51] & din_b[54])))) # (din_a[52] & (!din_b[53] $ (((!din_a[51]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_130  ) + ( Xd_0__inst_mult_7_129  ))
// Xd_0__inst_mult_7_137  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[54])))) # (din_a[52] & (!din_b[53] $ (((!din_a[51]) # (!din_b[54]))))) ) + ( Xd_0__inst_mult_7_130  ) + ( Xd_0__inst_mult_7_129  ))
// Xd_0__inst_mult_7_138  = SHARE((din_a[52] & (din_b[53] & (din_a[51] & din_b[54]))))

	.dataa(!din_a[52]),
	.datab(!din_b[53]),
	.datac(!din_a[51]),
	.datad(!din_b[54]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_129 ),
	.sharein(Xd_0__inst_mult_7_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_136 ),
	.cout(Xd_0__inst_mult_7_137 ),
	.shareout(Xd_0__inst_mult_7_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_40 (
// Equation(s):
// Xd_0__inst_mult_4_132  = SUM(( (!din_a[33] & (((din_a[32] & din_b[31])))) # (din_a[33] & (!din_b[30] $ (((!din_a[32]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_4_126  ) + ( Xd_0__inst_mult_4_125  ))
// Xd_0__inst_mult_4_133  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[31])))) # (din_a[33] & (!din_b[30] $ (((!din_a[32]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_4_126  ) + ( Xd_0__inst_mult_4_125  ))
// Xd_0__inst_mult_4_134  = SHARE((din_a[33] & (din_b[30] & (din_a[32] & din_b[31]))))

	.dataa(!din_a[33]),
	.datab(!din_b[30]),
	.datac(!din_a[32]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_125 ),
	.sharein(Xd_0__inst_mult_4_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_132 ),
	.cout(Xd_0__inst_mult_4_133 ),
	.shareout(Xd_0__inst_mult_4_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_41 (
// Equation(s):
// Xd_0__inst_mult_4_136  = SUM(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_130  ) + ( Xd_0__inst_mult_4_129  ))
// Xd_0__inst_mult_4_137  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_4_130  ) + ( Xd_0__inst_mult_4_129  ))
// Xd_0__inst_mult_4_138  = SHARE((din_a[31] & (din_b[32] & (din_a[30] & din_b[33]))))

	.dataa(!din_a[31]),
	.datab(!din_b[32]),
	.datac(!din_a[30]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_129 ),
	.sharein(Xd_0__inst_mult_4_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_136 ),
	.cout(Xd_0__inst_mult_4_137 ),
	.shareout(Xd_0__inst_mult_4_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_40 (
// Equation(s):
// Xd_0__inst_mult_5_132  = SUM(( (!din_a[40] & (((din_a[39] & din_b[38])))) # (din_a[40] & (!din_b[37] $ (((!din_a[39]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_5_126  ) + ( Xd_0__inst_mult_5_125  ))
// Xd_0__inst_mult_5_133  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[38])))) # (din_a[40] & (!din_b[37] $ (((!din_a[39]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_5_126  ) + ( Xd_0__inst_mult_5_125  ))
// Xd_0__inst_mult_5_134  = SHARE((din_a[40] & (din_b[37] & (din_a[39] & din_b[38]))))

	.dataa(!din_a[40]),
	.datab(!din_b[37]),
	.datac(!din_a[39]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_125 ),
	.sharein(Xd_0__inst_mult_5_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_132 ),
	.cout(Xd_0__inst_mult_5_133 ),
	.shareout(Xd_0__inst_mult_5_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_41 (
// Equation(s):
// Xd_0__inst_mult_5_136  = SUM(( (!din_a[38] & (((din_a[37] & din_b[40])))) # (din_a[38] & (!din_b[39] $ (((!din_a[37]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_130  ) + ( Xd_0__inst_mult_5_129  ))
// Xd_0__inst_mult_5_137  = CARRY(( (!din_a[38] & (((din_a[37] & din_b[40])))) # (din_a[38] & (!din_b[39] $ (((!din_a[37]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_5_130  ) + ( Xd_0__inst_mult_5_129  ))
// Xd_0__inst_mult_5_138  = SHARE((din_a[38] & (din_b[39] & (din_a[37] & din_b[40]))))

	.dataa(!din_a[38]),
	.datab(!din_b[39]),
	.datac(!din_a[37]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_129 ),
	.sharein(Xd_0__inst_mult_5_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_136 ),
	.cout(Xd_0__inst_mult_5_137 ),
	.shareout(Xd_0__inst_mult_5_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_40 (
// Equation(s):
// Xd_0__inst_mult_2_132  = SUM(( (!din_a[19] & (((din_a[18] & din_b[17])))) # (din_a[19] & (!din_b[16] $ (((!din_a[18]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_2_126  ) + ( Xd_0__inst_mult_2_125  ))
// Xd_0__inst_mult_2_133  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[17])))) # (din_a[19] & (!din_b[16] $ (((!din_a[18]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_2_126  ) + ( Xd_0__inst_mult_2_125  ))
// Xd_0__inst_mult_2_134  = SHARE((din_a[19] & (din_b[16] & (din_a[18] & din_b[17]))))

	.dataa(!din_a[19]),
	.datab(!din_b[16]),
	.datac(!din_a[18]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_125 ),
	.sharein(Xd_0__inst_mult_2_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_132 ),
	.cout(Xd_0__inst_mult_2_133 ),
	.shareout(Xd_0__inst_mult_2_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_41 (
// Equation(s):
// Xd_0__inst_mult_2_136  = SUM(( (!din_a[17] & (((din_a[16] & din_b[19])))) # (din_a[17] & (!din_b[18] $ (((!din_a[16]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_130  ) + ( Xd_0__inst_mult_2_129  ))
// Xd_0__inst_mult_2_137  = CARRY(( (!din_a[17] & (((din_a[16] & din_b[19])))) # (din_a[17] & (!din_b[18] $ (((!din_a[16]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_2_130  ) + ( Xd_0__inst_mult_2_129  ))
// Xd_0__inst_mult_2_138  = SHARE((din_a[17] & (din_b[18] & (din_a[16] & din_b[19]))))

	.dataa(!din_a[17]),
	.datab(!din_b[18]),
	.datac(!din_a[16]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_129 ),
	.sharein(Xd_0__inst_mult_2_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_136 ),
	.cout(Xd_0__inst_mult_2_137 ),
	.shareout(Xd_0__inst_mult_2_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_40 (
// Equation(s):
// Xd_0__inst_mult_3_132  = SUM(( (!din_a[26] & (((din_a[25] & din_b[24])))) # (din_a[26] & (!din_b[23] $ (((!din_a[25]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_3_126  ) + ( Xd_0__inst_mult_3_125  ))
// Xd_0__inst_mult_3_133  = CARRY(( (!din_a[26] & (((din_a[25] & din_b[24])))) # (din_a[26] & (!din_b[23] $ (((!din_a[25]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_3_126  ) + ( Xd_0__inst_mult_3_125  ))
// Xd_0__inst_mult_3_134  = SHARE((din_a[26] & (din_b[23] & (din_a[25] & din_b[24]))))

	.dataa(!din_a[26]),
	.datab(!din_b[23]),
	.datac(!din_a[25]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_125 ),
	.sharein(Xd_0__inst_mult_3_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_132 ),
	.cout(Xd_0__inst_mult_3_133 ),
	.shareout(Xd_0__inst_mult_3_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_41 (
// Equation(s):
// Xd_0__inst_mult_3_136  = SUM(( (!din_a[24] & (((din_a[23] & din_b[26])))) # (din_a[24] & (!din_b[25] $ (((!din_a[23]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_130  ) + ( Xd_0__inst_mult_3_129  ))
// Xd_0__inst_mult_3_137  = CARRY(( (!din_a[24] & (((din_a[23] & din_b[26])))) # (din_a[24] & (!din_b[25] $ (((!din_a[23]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_3_130  ) + ( Xd_0__inst_mult_3_129  ))
// Xd_0__inst_mult_3_138  = SHARE((din_a[24] & (din_b[25] & (din_a[23] & din_b[26]))))

	.dataa(!din_a[24]),
	.datab(!din_b[25]),
	.datac(!din_a[23]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_129 ),
	.sharein(Xd_0__inst_mult_3_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_136 ),
	.cout(Xd_0__inst_mult_3_137 ),
	.shareout(Xd_0__inst_mult_3_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_40 (
// Equation(s):
// Xd_0__inst_mult_0_132  = SUM(( (!din_a[5] & (((din_a[4] & din_b[3])))) # (din_a[5] & (!din_b[2] $ (((!din_a[4]) # (!din_b[3]))))) ) + ( Xd_0__inst_mult_0_126  ) + ( Xd_0__inst_mult_0_125  ))
// Xd_0__inst_mult_0_133  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[3])))) # (din_a[5] & (!din_b[2] $ (((!din_a[4]) # (!din_b[3]))))) ) + ( Xd_0__inst_mult_0_126  ) + ( Xd_0__inst_mult_0_125  ))
// Xd_0__inst_mult_0_134  = SHARE((din_a[5] & (din_b[2] & (din_a[4] & din_b[3]))))

	.dataa(!din_a[5]),
	.datab(!din_b[2]),
	.datac(!din_a[4]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_125 ),
	.sharein(Xd_0__inst_mult_0_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_132 ),
	.cout(Xd_0__inst_mult_0_133 ),
	.shareout(Xd_0__inst_mult_0_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_41 (
// Equation(s):
// Xd_0__inst_mult_0_136  = SUM(( (!din_a[3] & (((din_a[2] & din_b[5])))) # (din_a[3] & (!din_b[4] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_130  ) + ( Xd_0__inst_mult_0_129  ))
// Xd_0__inst_mult_0_137  = CARRY(( (!din_a[3] & (((din_a[2] & din_b[5])))) # (din_a[3] & (!din_b[4] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_130  ) + ( Xd_0__inst_mult_0_129  ))
// Xd_0__inst_mult_0_138  = SHARE((din_a[3] & (din_b[4] & (din_a[2] & din_b[5]))))

	.dataa(!din_a[3]),
	.datab(!din_b[4]),
	.datac(!din_a[2]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_129 ),
	.sharein(Xd_0__inst_mult_0_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_136 ),
	.cout(Xd_0__inst_mult_0_137 ),
	.shareout(Xd_0__inst_mult_0_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_40 (
// Equation(s):
// Xd_0__inst_mult_1_132  = SUM(( (!din_a[12] & (((din_a[11] & din_b[10])))) # (din_a[12] & (!din_b[9] $ (((!din_a[11]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_1_126  ) + ( Xd_0__inst_mult_1_125  ))
// Xd_0__inst_mult_1_133  = CARRY(( (!din_a[12] & (((din_a[11] & din_b[10])))) # (din_a[12] & (!din_b[9] $ (((!din_a[11]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_1_126  ) + ( Xd_0__inst_mult_1_125  ))
// Xd_0__inst_mult_1_134  = SHARE((din_a[12] & (din_b[9] & (din_a[11] & din_b[10]))))

	.dataa(!din_a[12]),
	.datab(!din_b[9]),
	.datac(!din_a[11]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_125 ),
	.sharein(Xd_0__inst_mult_1_126 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_132 ),
	.cout(Xd_0__inst_mult_1_133 ),
	.shareout(Xd_0__inst_mult_1_134 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_41 (
// Equation(s):
// Xd_0__inst_mult_1_136  = SUM(( (!din_a[10] & (((din_a[9] & din_b[12])))) # (din_a[10] & (!din_b[11] $ (((!din_a[9]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_130  ) + ( Xd_0__inst_mult_1_129  ))
// Xd_0__inst_mult_1_137  = CARRY(( (!din_a[10] & (((din_a[9] & din_b[12])))) # (din_a[10] & (!din_b[11] $ (((!din_a[9]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_130  ) + ( Xd_0__inst_mult_1_129  ))
// Xd_0__inst_mult_1_138  = SHARE((din_a[10] & (din_b[11] & (din_a[9] & din_b[12]))))

	.dataa(!din_a[10]),
	.datab(!din_b[11]),
	.datac(!din_a[9]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_129 ),
	.sharein(Xd_0__inst_mult_1_130 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_136 ),
	.cout(Xd_0__inst_mult_1_137 ),
	.shareout(Xd_0__inst_mult_1_138 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_42 (
// Equation(s):
// Xd_0__inst_mult_28_140  = SUM(( (!din_a[201] & (((din_a[200] & din_b[200])))) # (din_a[201] & (!din_b[199] $ (((!din_a[200]) # (!din_b[200]))))) ) + ( Xd_0__inst_mult_28_134  ) + ( Xd_0__inst_mult_28_133  ))
// Xd_0__inst_mult_28_141  = CARRY(( (!din_a[201] & (((din_a[200] & din_b[200])))) # (din_a[201] & (!din_b[199] $ (((!din_a[200]) # (!din_b[200]))))) ) + ( Xd_0__inst_mult_28_134  ) + ( Xd_0__inst_mult_28_133  ))
// Xd_0__inst_mult_28_142  = SHARE((din_a[201] & (din_b[199] & (din_a[200] & din_b[200]))))

	.dataa(!din_a[201]),
	.datab(!din_b[199]),
	.datac(!din_a[200]),
	.datad(!din_b[200]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_133 ),
	.sharein(Xd_0__inst_mult_28_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_140 ),
	.cout(Xd_0__inst_mult_28_141 ),
	.shareout(Xd_0__inst_mult_28_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_43 (
// Equation(s):
// Xd_0__inst_mult_28_144  = SUM(( (din_a[199] & din_b[201]) ) + ( Xd_0__inst_mult_28_138  ) + ( Xd_0__inst_mult_28_137  ))
// Xd_0__inst_mult_28_145  = CARRY(( (din_a[199] & din_b[201]) ) + ( Xd_0__inst_mult_28_138  ) + ( Xd_0__inst_mult_28_137  ))
// Xd_0__inst_mult_28_146  = SHARE(GND)

	.dataa(!din_a[199]),
	.datab(!din_b[201]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_137 ),
	.sharein(Xd_0__inst_mult_28_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_144 ),
	.cout(Xd_0__inst_mult_28_145 ),
	.shareout(Xd_0__inst_mult_28_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_42 (
// Equation(s):
// Xd_0__inst_mult_29_140  = SUM(( (!din_a[208] & (((din_a[207] & din_b[207])))) # (din_a[208] & (!din_b[206] $ (((!din_a[207]) # (!din_b[207]))))) ) + ( Xd_0__inst_mult_29_134  ) + ( Xd_0__inst_mult_29_133  ))
// Xd_0__inst_mult_29_141  = CARRY(( (!din_a[208] & (((din_a[207] & din_b[207])))) # (din_a[208] & (!din_b[206] $ (((!din_a[207]) # (!din_b[207]))))) ) + ( Xd_0__inst_mult_29_134  ) + ( Xd_0__inst_mult_29_133  ))
// Xd_0__inst_mult_29_142  = SHARE((din_a[208] & (din_b[206] & (din_a[207] & din_b[207]))))

	.dataa(!din_a[208]),
	.datab(!din_b[206]),
	.datac(!din_a[207]),
	.datad(!din_b[207]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_133 ),
	.sharein(Xd_0__inst_mult_29_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_140 ),
	.cout(Xd_0__inst_mult_29_141 ),
	.shareout(Xd_0__inst_mult_29_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_43 (
// Equation(s):
// Xd_0__inst_mult_29_144  = SUM(( (din_a[206] & din_b[208]) ) + ( Xd_0__inst_mult_29_138  ) + ( Xd_0__inst_mult_29_137  ))
// Xd_0__inst_mult_29_145  = CARRY(( (din_a[206] & din_b[208]) ) + ( Xd_0__inst_mult_29_138  ) + ( Xd_0__inst_mult_29_137  ))
// Xd_0__inst_mult_29_146  = SHARE(GND)

	.dataa(!din_a[206]),
	.datab(!din_b[208]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_137 ),
	.sharein(Xd_0__inst_mult_29_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_144 ),
	.cout(Xd_0__inst_mult_29_145 ),
	.shareout(Xd_0__inst_mult_29_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_42 (
// Equation(s):
// Xd_0__inst_mult_26_140  = SUM(( (!din_a[187] & (((din_a[186] & din_b[186])))) # (din_a[187] & (!din_b[185] $ (((!din_a[186]) # (!din_b[186]))))) ) + ( Xd_0__inst_mult_26_134  ) + ( Xd_0__inst_mult_26_133  ))
// Xd_0__inst_mult_26_141  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[186])))) # (din_a[187] & (!din_b[185] $ (((!din_a[186]) # (!din_b[186]))))) ) + ( Xd_0__inst_mult_26_134  ) + ( Xd_0__inst_mult_26_133  ))
// Xd_0__inst_mult_26_142  = SHARE((din_a[187] & (din_b[185] & (din_a[186] & din_b[186]))))

	.dataa(!din_a[187]),
	.datab(!din_b[185]),
	.datac(!din_a[186]),
	.datad(!din_b[186]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_133 ),
	.sharein(Xd_0__inst_mult_26_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_140 ),
	.cout(Xd_0__inst_mult_26_141 ),
	.shareout(Xd_0__inst_mult_26_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_43 (
// Equation(s):
// Xd_0__inst_mult_26_144  = SUM(( (din_a[185] & din_b[187]) ) + ( Xd_0__inst_mult_26_138  ) + ( Xd_0__inst_mult_26_137  ))
// Xd_0__inst_mult_26_145  = CARRY(( (din_a[185] & din_b[187]) ) + ( Xd_0__inst_mult_26_138  ) + ( Xd_0__inst_mult_26_137  ))
// Xd_0__inst_mult_26_146  = SHARE(GND)

	.dataa(!din_a[185]),
	.datab(!din_b[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_137 ),
	.sharein(Xd_0__inst_mult_26_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_144 ),
	.cout(Xd_0__inst_mult_26_145 ),
	.shareout(Xd_0__inst_mult_26_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_42 (
// Equation(s):
// Xd_0__inst_mult_27_140  = SUM(( (!din_a[194] & (((din_a[193] & din_b[193])))) # (din_a[194] & (!din_b[192] $ (((!din_a[193]) # (!din_b[193]))))) ) + ( Xd_0__inst_mult_27_134  ) + ( Xd_0__inst_mult_27_133  ))
// Xd_0__inst_mult_27_141  = CARRY(( (!din_a[194] & (((din_a[193] & din_b[193])))) # (din_a[194] & (!din_b[192] $ (((!din_a[193]) # (!din_b[193]))))) ) + ( Xd_0__inst_mult_27_134  ) + ( Xd_0__inst_mult_27_133  ))
// Xd_0__inst_mult_27_142  = SHARE((din_a[194] & (din_b[192] & (din_a[193] & din_b[193]))))

	.dataa(!din_a[194]),
	.datab(!din_b[192]),
	.datac(!din_a[193]),
	.datad(!din_b[193]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_133 ),
	.sharein(Xd_0__inst_mult_27_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_140 ),
	.cout(Xd_0__inst_mult_27_141 ),
	.shareout(Xd_0__inst_mult_27_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_43 (
// Equation(s):
// Xd_0__inst_mult_27_144  = SUM(( (din_a[192] & din_b[194]) ) + ( Xd_0__inst_mult_27_138  ) + ( Xd_0__inst_mult_27_137  ))
// Xd_0__inst_mult_27_145  = CARRY(( (din_a[192] & din_b[194]) ) + ( Xd_0__inst_mult_27_138  ) + ( Xd_0__inst_mult_27_137  ))
// Xd_0__inst_mult_27_146  = SHARE(GND)

	.dataa(!din_a[192]),
	.datab(!din_b[194]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_137 ),
	.sharein(Xd_0__inst_mult_27_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_144 ),
	.cout(Xd_0__inst_mult_27_145 ),
	.shareout(Xd_0__inst_mult_27_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_42 (
// Equation(s):
// Xd_0__inst_mult_24_140  = SUM(( (!din_a[173] & (((din_a[172] & din_b[172])))) # (din_a[173] & (!din_b[171] $ (((!din_a[172]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_24_134  ) + ( Xd_0__inst_mult_24_133  ))
// Xd_0__inst_mult_24_141  = CARRY(( (!din_a[173] & (((din_a[172] & din_b[172])))) # (din_a[173] & (!din_b[171] $ (((!din_a[172]) # (!din_b[172]))))) ) + ( Xd_0__inst_mult_24_134  ) + ( Xd_0__inst_mult_24_133  ))
// Xd_0__inst_mult_24_142  = SHARE((din_a[173] & (din_b[171] & (din_a[172] & din_b[172]))))

	.dataa(!din_a[173]),
	.datab(!din_b[171]),
	.datac(!din_a[172]),
	.datad(!din_b[172]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_133 ),
	.sharein(Xd_0__inst_mult_24_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_140 ),
	.cout(Xd_0__inst_mult_24_141 ),
	.shareout(Xd_0__inst_mult_24_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_43 (
// Equation(s):
// Xd_0__inst_mult_24_144  = SUM(( (din_a[171] & din_b[173]) ) + ( Xd_0__inst_mult_24_138  ) + ( Xd_0__inst_mult_24_137  ))
// Xd_0__inst_mult_24_145  = CARRY(( (din_a[171] & din_b[173]) ) + ( Xd_0__inst_mult_24_138  ) + ( Xd_0__inst_mult_24_137  ))
// Xd_0__inst_mult_24_146  = SHARE(GND)

	.dataa(!din_a[171]),
	.datab(!din_b[173]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_137 ),
	.sharein(Xd_0__inst_mult_24_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_144 ),
	.cout(Xd_0__inst_mult_24_145 ),
	.shareout(Xd_0__inst_mult_24_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_43 (
// Equation(s):
// Xd_0__inst_mult_25_144  = SUM(( (!din_a[180] & (((din_a[179] & din_b[179])))) # (din_a[180] & (!din_b[178] $ (((!din_a[179]) # (!din_b[179]))))) ) + ( Xd_0__inst_mult_25_138  ) + ( Xd_0__inst_mult_25_137  ))
// Xd_0__inst_mult_25_145  = CARRY(( (!din_a[180] & (((din_a[179] & din_b[179])))) # (din_a[180] & (!din_b[178] $ (((!din_a[179]) # (!din_b[179]))))) ) + ( Xd_0__inst_mult_25_138  ) + ( Xd_0__inst_mult_25_137  ))
// Xd_0__inst_mult_25_146  = SHARE((din_a[180] & (din_b[178] & (din_a[179] & din_b[179]))))

	.dataa(!din_a[180]),
	.datab(!din_b[178]),
	.datac(!din_a[179]),
	.datad(!din_b[179]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_137 ),
	.sharein(Xd_0__inst_mult_25_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_144 ),
	.cout(Xd_0__inst_mult_25_145 ),
	.shareout(Xd_0__inst_mult_25_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_43 (
// Equation(s):
// Xd_0__inst_mult_22_144  = SUM(( (!din_a[159] & (((din_a[158] & din_b[158])))) # (din_a[159] & (!din_b[157] $ (((!din_a[158]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_22_138  ) + ( Xd_0__inst_mult_22_137  ))
// Xd_0__inst_mult_22_145  = CARRY(( (!din_a[159] & (((din_a[158] & din_b[158])))) # (din_a[159] & (!din_b[157] $ (((!din_a[158]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_22_138  ) + ( Xd_0__inst_mult_22_137  ))
// Xd_0__inst_mult_22_146  = SHARE((din_a[159] & (din_b[157] & (din_a[158] & din_b[158]))))

	.dataa(!din_a[159]),
	.datab(!din_b[157]),
	.datac(!din_a[158]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_137 ),
	.sharein(Xd_0__inst_mult_22_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_144 ),
	.cout(Xd_0__inst_mult_22_145 ),
	.shareout(Xd_0__inst_mult_22_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_42 (
// Equation(s):
// Xd_0__inst_mult_23_140  = SUM(( (!din_a[166] & (((din_a[165] & din_b[165])))) # (din_a[166] & (!din_b[164] $ (((!din_a[165]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_23_134  ) + ( Xd_0__inst_mult_23_133  ))
// Xd_0__inst_mult_23_141  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[165])))) # (din_a[166] & (!din_b[164] $ (((!din_a[165]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_23_134  ) + ( Xd_0__inst_mult_23_133  ))
// Xd_0__inst_mult_23_142  = SHARE((din_a[166] & (din_b[164] & (din_a[165] & din_b[165]))))

	.dataa(!din_a[166]),
	.datab(!din_b[164]),
	.datac(!din_a[165]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_133 ),
	.sharein(Xd_0__inst_mult_23_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_140 ),
	.cout(Xd_0__inst_mult_23_141 ),
	.shareout(Xd_0__inst_mult_23_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_43 (
// Equation(s):
// Xd_0__inst_mult_23_144  = SUM(( (din_a[164] & din_b[166]) ) + ( Xd_0__inst_mult_23_138  ) + ( Xd_0__inst_mult_23_137  ))
// Xd_0__inst_mult_23_145  = CARRY(( (din_a[164] & din_b[166]) ) + ( Xd_0__inst_mult_23_138  ) + ( Xd_0__inst_mult_23_137  ))
// Xd_0__inst_mult_23_146  = SHARE(GND)

	.dataa(!din_a[164]),
	.datab(!din_b[166]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_137 ),
	.sharein(Xd_0__inst_mult_23_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_144 ),
	.cout(Xd_0__inst_mult_23_145 ),
	.shareout(Xd_0__inst_mult_23_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_42 (
// Equation(s):
// Xd_0__inst_mult_20_140  = SUM(( (!din_a[145] & (((din_a[144] & din_b[144])))) # (din_a[145] & (!din_b[143] $ (((!din_a[144]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_20_134  ) + ( Xd_0__inst_mult_20_133  ))
// Xd_0__inst_mult_20_141  = CARRY(( (!din_a[145] & (((din_a[144] & din_b[144])))) # (din_a[145] & (!din_b[143] $ (((!din_a[144]) # (!din_b[144]))))) ) + ( Xd_0__inst_mult_20_134  ) + ( Xd_0__inst_mult_20_133  ))
// Xd_0__inst_mult_20_142  = SHARE((din_a[145] & (din_b[143] & (din_a[144] & din_b[144]))))

	.dataa(!din_a[145]),
	.datab(!din_b[143]),
	.datac(!din_a[144]),
	.datad(!din_b[144]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_133 ),
	.sharein(Xd_0__inst_mult_20_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_140 ),
	.cout(Xd_0__inst_mult_20_141 ),
	.shareout(Xd_0__inst_mult_20_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_43 (
// Equation(s):
// Xd_0__inst_mult_20_144  = SUM(( (din_a[143] & din_b[145]) ) + ( Xd_0__inst_mult_20_138  ) + ( Xd_0__inst_mult_20_137  ))
// Xd_0__inst_mult_20_145  = CARRY(( (din_a[143] & din_b[145]) ) + ( Xd_0__inst_mult_20_138  ) + ( Xd_0__inst_mult_20_137  ))
// Xd_0__inst_mult_20_146  = SHARE(GND)

	.dataa(!din_a[143]),
	.datab(!din_b[145]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_137 ),
	.sharein(Xd_0__inst_mult_20_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_144 ),
	.cout(Xd_0__inst_mult_20_145 ),
	.shareout(Xd_0__inst_mult_20_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_42 (
// Equation(s):
// Xd_0__inst_mult_21_140  = SUM(( (!din_a[152] & (((din_a[151] & din_b[151])))) # (din_a[152] & (!din_b[150] $ (((!din_a[151]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_21_134  ) + ( Xd_0__inst_mult_21_133  ))
// Xd_0__inst_mult_21_141  = CARRY(( (!din_a[152] & (((din_a[151] & din_b[151])))) # (din_a[152] & (!din_b[150] $ (((!din_a[151]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_21_134  ) + ( Xd_0__inst_mult_21_133  ))
// Xd_0__inst_mult_21_142  = SHARE((din_a[152] & (din_b[150] & (din_a[151] & din_b[151]))))

	.dataa(!din_a[152]),
	.datab(!din_b[150]),
	.datac(!din_a[151]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_133 ),
	.sharein(Xd_0__inst_mult_21_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_140 ),
	.cout(Xd_0__inst_mult_21_141 ),
	.shareout(Xd_0__inst_mult_21_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_43 (
// Equation(s):
// Xd_0__inst_mult_21_144  = SUM(( (din_a[150] & din_b[152]) ) + ( Xd_0__inst_mult_21_138  ) + ( Xd_0__inst_mult_21_137  ))
// Xd_0__inst_mult_21_145  = CARRY(( (din_a[150] & din_b[152]) ) + ( Xd_0__inst_mult_21_138  ) + ( Xd_0__inst_mult_21_137  ))
// Xd_0__inst_mult_21_146  = SHARE(GND)

	.dataa(!din_a[150]),
	.datab(!din_b[152]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_137 ),
	.sharein(Xd_0__inst_mult_21_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_144 ),
	.cout(Xd_0__inst_mult_21_145 ),
	.shareout(Xd_0__inst_mult_21_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_42 (
// Equation(s):
// Xd_0__inst_mult_18_140  = SUM(( (!din_a[131] & (((din_a[130] & din_b[130])))) # (din_a[131] & (!din_b[129] $ (((!din_a[130]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_18_134  ) + ( Xd_0__inst_mult_18_133  ))
// Xd_0__inst_mult_18_141  = CARRY(( (!din_a[131] & (((din_a[130] & din_b[130])))) # (din_a[131] & (!din_b[129] $ (((!din_a[130]) # (!din_b[130]))))) ) + ( Xd_0__inst_mult_18_134  ) + ( Xd_0__inst_mult_18_133  ))
// Xd_0__inst_mult_18_142  = SHARE((din_a[131] & (din_b[129] & (din_a[130] & din_b[130]))))

	.dataa(!din_a[131]),
	.datab(!din_b[129]),
	.datac(!din_a[130]),
	.datad(!din_b[130]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_133 ),
	.sharein(Xd_0__inst_mult_18_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_140 ),
	.cout(Xd_0__inst_mult_18_141 ),
	.shareout(Xd_0__inst_mult_18_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_43 (
// Equation(s):
// Xd_0__inst_mult_18_144  = SUM(( (din_a[129] & din_b[131]) ) + ( Xd_0__inst_mult_18_138  ) + ( Xd_0__inst_mult_18_137  ))
// Xd_0__inst_mult_18_145  = CARRY(( (din_a[129] & din_b[131]) ) + ( Xd_0__inst_mult_18_138  ) + ( Xd_0__inst_mult_18_137  ))
// Xd_0__inst_mult_18_146  = SHARE(GND)

	.dataa(!din_a[129]),
	.datab(!din_b[131]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_137 ),
	.sharein(Xd_0__inst_mult_18_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_144 ),
	.cout(Xd_0__inst_mult_18_145 ),
	.shareout(Xd_0__inst_mult_18_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_42 (
// Equation(s):
// Xd_0__inst_mult_19_140  = SUM(( (!din_a[138] & (((din_a[137] & din_b[137])))) # (din_a[138] & (!din_b[136] $ (((!din_a[137]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_19_134  ) + ( Xd_0__inst_mult_19_133  ))
// Xd_0__inst_mult_19_141  = CARRY(( (!din_a[138] & (((din_a[137] & din_b[137])))) # (din_a[138] & (!din_b[136] $ (((!din_a[137]) # (!din_b[137]))))) ) + ( Xd_0__inst_mult_19_134  ) + ( Xd_0__inst_mult_19_133  ))
// Xd_0__inst_mult_19_142  = SHARE((din_a[138] & (din_b[136] & (din_a[137] & din_b[137]))))

	.dataa(!din_a[138]),
	.datab(!din_b[136]),
	.datac(!din_a[137]),
	.datad(!din_b[137]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_133 ),
	.sharein(Xd_0__inst_mult_19_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_140 ),
	.cout(Xd_0__inst_mult_19_141 ),
	.shareout(Xd_0__inst_mult_19_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_43 (
// Equation(s):
// Xd_0__inst_mult_19_144  = SUM(( (din_a[136] & din_b[138]) ) + ( Xd_0__inst_mult_19_138  ) + ( Xd_0__inst_mult_19_137  ))
// Xd_0__inst_mult_19_145  = CARRY(( (din_a[136] & din_b[138]) ) + ( Xd_0__inst_mult_19_138  ) + ( Xd_0__inst_mult_19_137  ))
// Xd_0__inst_mult_19_146  = SHARE(GND)

	.dataa(!din_a[136]),
	.datab(!din_b[138]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_137 ),
	.sharein(Xd_0__inst_mult_19_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_144 ),
	.cout(Xd_0__inst_mult_19_145 ),
	.shareout(Xd_0__inst_mult_19_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_42 (
// Equation(s):
// Xd_0__inst_mult_16_140  = SUM(( (!din_a[117] & (((din_a[116] & din_b[116])))) # (din_a[117] & (!din_b[115] $ (((!din_a[116]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_16_134  ) + ( Xd_0__inst_mult_16_133  ))
// Xd_0__inst_mult_16_141  = CARRY(( (!din_a[117] & (((din_a[116] & din_b[116])))) # (din_a[117] & (!din_b[115] $ (((!din_a[116]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_16_134  ) + ( Xd_0__inst_mult_16_133  ))
// Xd_0__inst_mult_16_142  = SHARE((din_a[117] & (din_b[115] & (din_a[116] & din_b[116]))))

	.dataa(!din_a[117]),
	.datab(!din_b[115]),
	.datac(!din_a[116]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_133 ),
	.sharein(Xd_0__inst_mult_16_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_140 ),
	.cout(Xd_0__inst_mult_16_141 ),
	.shareout(Xd_0__inst_mult_16_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_43 (
// Equation(s):
// Xd_0__inst_mult_16_144  = SUM(( (din_a[115] & din_b[117]) ) + ( Xd_0__inst_mult_16_138  ) + ( Xd_0__inst_mult_16_137  ))
// Xd_0__inst_mult_16_145  = CARRY(( (din_a[115] & din_b[117]) ) + ( Xd_0__inst_mult_16_138  ) + ( Xd_0__inst_mult_16_137  ))
// Xd_0__inst_mult_16_146  = SHARE(GND)

	.dataa(!din_a[115]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_137 ),
	.sharein(Xd_0__inst_mult_16_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_144 ),
	.cout(Xd_0__inst_mult_16_145 ),
	.shareout(Xd_0__inst_mult_16_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_42 (
// Equation(s):
// Xd_0__inst_mult_17_140  = SUM(( (!din_a[124] & (((din_a[123] & din_b[123])))) # (din_a[124] & (!din_b[122] $ (((!din_a[123]) # (!din_b[123]))))) ) + ( Xd_0__inst_mult_17_134  ) + ( Xd_0__inst_mult_17_133  ))
// Xd_0__inst_mult_17_141  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[123])))) # (din_a[124] & (!din_b[122] $ (((!din_a[123]) # (!din_b[123]))))) ) + ( Xd_0__inst_mult_17_134  ) + ( Xd_0__inst_mult_17_133  ))
// Xd_0__inst_mult_17_142  = SHARE((din_a[124] & (din_b[122] & (din_a[123] & din_b[123]))))

	.dataa(!din_a[124]),
	.datab(!din_b[122]),
	.datac(!din_a[123]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_133 ),
	.sharein(Xd_0__inst_mult_17_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_140 ),
	.cout(Xd_0__inst_mult_17_141 ),
	.shareout(Xd_0__inst_mult_17_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_43 (
// Equation(s):
// Xd_0__inst_mult_17_144  = SUM(( (din_a[122] & din_b[124]) ) + ( Xd_0__inst_mult_17_138  ) + ( Xd_0__inst_mult_17_137  ))
// Xd_0__inst_mult_17_145  = CARRY(( (din_a[122] & din_b[124]) ) + ( Xd_0__inst_mult_17_138  ) + ( Xd_0__inst_mult_17_137  ))
// Xd_0__inst_mult_17_146  = SHARE(GND)

	.dataa(!din_a[122]),
	.datab(!din_b[124]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_137 ),
	.sharein(Xd_0__inst_mult_17_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_144 ),
	.cout(Xd_0__inst_mult_17_145 ),
	.shareout(Xd_0__inst_mult_17_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_42 (
// Equation(s):
// Xd_0__inst_mult_14_140  = SUM(( (!din_a[103] & (((din_a[102] & din_b[102])))) # (din_a[103] & (!din_b[101] $ (((!din_a[102]) # (!din_b[102]))))) ) + ( Xd_0__inst_mult_14_134  ) + ( Xd_0__inst_mult_14_133  ))
// Xd_0__inst_mult_14_141  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[102])))) # (din_a[103] & (!din_b[101] $ (((!din_a[102]) # (!din_b[102]))))) ) + ( Xd_0__inst_mult_14_134  ) + ( Xd_0__inst_mult_14_133  ))
// Xd_0__inst_mult_14_142  = SHARE((din_a[103] & (din_b[101] & (din_a[102] & din_b[102]))))

	.dataa(!din_a[103]),
	.datab(!din_b[101]),
	.datac(!din_a[102]),
	.datad(!din_b[102]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_133 ),
	.sharein(Xd_0__inst_mult_14_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_140 ),
	.cout(Xd_0__inst_mult_14_141 ),
	.shareout(Xd_0__inst_mult_14_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_43 (
// Equation(s):
// Xd_0__inst_mult_14_144  = SUM(( (din_a[101] & din_b[103]) ) + ( Xd_0__inst_mult_14_138  ) + ( Xd_0__inst_mult_14_137  ))
// Xd_0__inst_mult_14_145  = CARRY(( (din_a[101] & din_b[103]) ) + ( Xd_0__inst_mult_14_138  ) + ( Xd_0__inst_mult_14_137  ))
// Xd_0__inst_mult_14_146  = SHARE(GND)

	.dataa(!din_a[101]),
	.datab(!din_b[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_137 ),
	.sharein(Xd_0__inst_mult_14_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_144 ),
	.cout(Xd_0__inst_mult_14_145 ),
	.shareout(Xd_0__inst_mult_14_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_42 (
// Equation(s):
// Xd_0__inst_mult_15_140  = SUM(( (!din_a[110] & (((din_a[109] & din_b[109])))) # (din_a[110] & (!din_b[108] $ (((!din_a[109]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_15_134  ) + ( Xd_0__inst_mult_15_133  ))
// Xd_0__inst_mult_15_141  = CARRY(( (!din_a[110] & (((din_a[109] & din_b[109])))) # (din_a[110] & (!din_b[108] $ (((!din_a[109]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_15_134  ) + ( Xd_0__inst_mult_15_133  ))
// Xd_0__inst_mult_15_142  = SHARE((din_a[110] & (din_b[108] & (din_a[109] & din_b[109]))))

	.dataa(!din_a[110]),
	.datab(!din_b[108]),
	.datac(!din_a[109]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_133 ),
	.sharein(Xd_0__inst_mult_15_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_140 ),
	.cout(Xd_0__inst_mult_15_141 ),
	.shareout(Xd_0__inst_mult_15_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_43 (
// Equation(s):
// Xd_0__inst_mult_15_144  = SUM(( (din_a[108] & din_b[110]) ) + ( Xd_0__inst_mult_15_138  ) + ( Xd_0__inst_mult_15_137  ))
// Xd_0__inst_mult_15_145  = CARRY(( (din_a[108] & din_b[110]) ) + ( Xd_0__inst_mult_15_138  ) + ( Xd_0__inst_mult_15_137  ))
// Xd_0__inst_mult_15_146  = SHARE(GND)

	.dataa(!din_a[108]),
	.datab(!din_b[110]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_137 ),
	.sharein(Xd_0__inst_mult_15_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_144 ),
	.cout(Xd_0__inst_mult_15_145 ),
	.shareout(Xd_0__inst_mult_15_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_42 (
// Equation(s):
// Xd_0__inst_mult_12_140  = SUM(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_12_134  ) + ( Xd_0__inst_mult_12_133  ))
// Xd_0__inst_mult_12_141  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_12_134  ) + ( Xd_0__inst_mult_12_133  ))
// Xd_0__inst_mult_12_142  = SHARE((din_a[89] & (din_b[87] & (din_a[88] & din_b[88]))))

	.dataa(!din_a[89]),
	.datab(!din_b[87]),
	.datac(!din_a[88]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_133 ),
	.sharein(Xd_0__inst_mult_12_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_140 ),
	.cout(Xd_0__inst_mult_12_141 ),
	.shareout(Xd_0__inst_mult_12_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_43 (
// Equation(s):
// Xd_0__inst_mult_12_144  = SUM(( (din_a[87] & din_b[89]) ) + ( Xd_0__inst_mult_12_138  ) + ( Xd_0__inst_mult_12_137  ))
// Xd_0__inst_mult_12_145  = CARRY(( (din_a[87] & din_b[89]) ) + ( Xd_0__inst_mult_12_138  ) + ( Xd_0__inst_mult_12_137  ))
// Xd_0__inst_mult_12_146  = SHARE(GND)

	.dataa(!din_a[87]),
	.datab(!din_b[89]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_137 ),
	.sharein(Xd_0__inst_mult_12_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_144 ),
	.cout(Xd_0__inst_mult_12_145 ),
	.shareout(Xd_0__inst_mult_12_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_42 (
// Equation(s):
// Xd_0__inst_mult_13_140  = SUM(( (!din_a[96] & (((din_a[95] & din_b[95])))) # (din_a[96] & (!din_b[94] $ (((!din_a[95]) # (!din_b[95]))))) ) + ( Xd_0__inst_mult_13_134  ) + ( Xd_0__inst_mult_13_133  ))
// Xd_0__inst_mult_13_141  = CARRY(( (!din_a[96] & (((din_a[95] & din_b[95])))) # (din_a[96] & (!din_b[94] $ (((!din_a[95]) # (!din_b[95]))))) ) + ( Xd_0__inst_mult_13_134  ) + ( Xd_0__inst_mult_13_133  ))
// Xd_0__inst_mult_13_142  = SHARE((din_a[96] & (din_b[94] & (din_a[95] & din_b[95]))))

	.dataa(!din_a[96]),
	.datab(!din_b[94]),
	.datac(!din_a[95]),
	.datad(!din_b[95]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_133 ),
	.sharein(Xd_0__inst_mult_13_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_140 ),
	.cout(Xd_0__inst_mult_13_141 ),
	.shareout(Xd_0__inst_mult_13_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_43 (
// Equation(s):
// Xd_0__inst_mult_13_144  = SUM(( (din_a[94] & din_b[96]) ) + ( Xd_0__inst_mult_13_138  ) + ( Xd_0__inst_mult_13_137  ))
// Xd_0__inst_mult_13_145  = CARRY(( (din_a[94] & din_b[96]) ) + ( Xd_0__inst_mult_13_138  ) + ( Xd_0__inst_mult_13_137  ))
// Xd_0__inst_mult_13_146  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[96]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_137 ),
	.sharein(Xd_0__inst_mult_13_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_144 ),
	.cout(Xd_0__inst_mult_13_145 ),
	.shareout(Xd_0__inst_mult_13_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_42 (
// Equation(s):
// Xd_0__inst_mult_10_140  = SUM(( (!din_a[75] & (((din_a[74] & din_b[74])))) # (din_a[75] & (!din_b[73] $ (((!din_a[74]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_10_134  ) + ( Xd_0__inst_mult_10_133  ))
// Xd_0__inst_mult_10_141  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[74])))) # (din_a[75] & (!din_b[73] $ (((!din_a[74]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_10_134  ) + ( Xd_0__inst_mult_10_133  ))
// Xd_0__inst_mult_10_142  = SHARE((din_a[75] & (din_b[73] & (din_a[74] & din_b[74]))))

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_133 ),
	.sharein(Xd_0__inst_mult_10_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_140 ),
	.cout(Xd_0__inst_mult_10_141 ),
	.shareout(Xd_0__inst_mult_10_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_43 (
// Equation(s):
// Xd_0__inst_mult_10_144  = SUM(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_10_138  ) + ( Xd_0__inst_mult_10_137  ))
// Xd_0__inst_mult_10_145  = CARRY(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_10_138  ) + ( Xd_0__inst_mult_10_137  ))
// Xd_0__inst_mult_10_146  = SHARE(GND)

	.dataa(!din_a[73]),
	.datab(!din_b[75]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_137 ),
	.sharein(Xd_0__inst_mult_10_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_144 ),
	.cout(Xd_0__inst_mult_10_145 ),
	.shareout(Xd_0__inst_mult_10_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_42 (
// Equation(s):
// Xd_0__inst_mult_11_140  = SUM(( (!din_a[82] & (((din_a[81] & din_b[81])))) # (din_a[82] & (!din_b[80] $ (((!din_a[81]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_11_134  ) + ( Xd_0__inst_mult_11_133  ))
// Xd_0__inst_mult_11_141  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[81])))) # (din_a[82] & (!din_b[80] $ (((!din_a[81]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_11_134  ) + ( Xd_0__inst_mult_11_133  ))
// Xd_0__inst_mult_11_142  = SHARE((din_a[82] & (din_b[80] & (din_a[81] & din_b[81]))))

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(!din_a[81]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_133 ),
	.sharein(Xd_0__inst_mult_11_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_140 ),
	.cout(Xd_0__inst_mult_11_141 ),
	.shareout(Xd_0__inst_mult_11_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_43 (
// Equation(s):
// Xd_0__inst_mult_11_144  = SUM(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_11_138  ) + ( Xd_0__inst_mult_11_137  ))
// Xd_0__inst_mult_11_145  = CARRY(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_11_138  ) + ( Xd_0__inst_mult_11_137  ))
// Xd_0__inst_mult_11_146  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_137 ),
	.sharein(Xd_0__inst_mult_11_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_144 ),
	.cout(Xd_0__inst_mult_11_145 ),
	.shareout(Xd_0__inst_mult_11_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_42 (
// Equation(s):
// Xd_0__inst_mult_8_140  = SUM(( (!din_a[61] & (((din_a[60] & din_b[60])))) # (din_a[61] & (!din_b[59] $ (((!din_a[60]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_8_134  ) + ( Xd_0__inst_mult_8_133  ))
// Xd_0__inst_mult_8_141  = CARRY(( (!din_a[61] & (((din_a[60] & din_b[60])))) # (din_a[61] & (!din_b[59] $ (((!din_a[60]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_8_134  ) + ( Xd_0__inst_mult_8_133  ))
// Xd_0__inst_mult_8_142  = SHARE((din_a[61] & (din_b[59] & (din_a[60] & din_b[60]))))

	.dataa(!din_a[61]),
	.datab(!din_b[59]),
	.datac(!din_a[60]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_133 ),
	.sharein(Xd_0__inst_mult_8_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_140 ),
	.cout(Xd_0__inst_mult_8_141 ),
	.shareout(Xd_0__inst_mult_8_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_43 (
// Equation(s):
// Xd_0__inst_mult_8_144  = SUM(( (din_a[59] & din_b[61]) ) + ( Xd_0__inst_mult_8_138  ) + ( Xd_0__inst_mult_8_137  ))
// Xd_0__inst_mult_8_145  = CARRY(( (din_a[59] & din_b[61]) ) + ( Xd_0__inst_mult_8_138  ) + ( Xd_0__inst_mult_8_137  ))
// Xd_0__inst_mult_8_146  = SHARE(GND)

	.dataa(!din_a[59]),
	.datab(!din_b[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_137 ),
	.sharein(Xd_0__inst_mult_8_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_144 ),
	.cout(Xd_0__inst_mult_8_145 ),
	.shareout(Xd_0__inst_mult_8_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_42 (
// Equation(s):
// Xd_0__inst_mult_9_140  = SUM(( (!din_a[68] & (((din_a[67] & din_b[67])))) # (din_a[68] & (!din_b[66] $ (((!din_a[67]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_9_134  ) + ( Xd_0__inst_mult_9_133  ))
// Xd_0__inst_mult_9_141  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[67])))) # (din_a[68] & (!din_b[66] $ (((!din_a[67]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_9_134  ) + ( Xd_0__inst_mult_9_133  ))
// Xd_0__inst_mult_9_142  = SHARE((din_a[68] & (din_b[66] & (din_a[67] & din_b[67]))))

	.dataa(!din_a[68]),
	.datab(!din_b[66]),
	.datac(!din_a[67]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_133 ),
	.sharein(Xd_0__inst_mult_9_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_140 ),
	.cout(Xd_0__inst_mult_9_141 ),
	.shareout(Xd_0__inst_mult_9_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_43 (
// Equation(s):
// Xd_0__inst_mult_9_144  = SUM(( (din_a[66] & din_b[68]) ) + ( Xd_0__inst_mult_9_138  ) + ( Xd_0__inst_mult_9_137  ))
// Xd_0__inst_mult_9_145  = CARRY(( (din_a[66] & din_b[68]) ) + ( Xd_0__inst_mult_9_138  ) + ( Xd_0__inst_mult_9_137  ))
// Xd_0__inst_mult_9_146  = SHARE(GND)

	.dataa(!din_a[66]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_137 ),
	.sharein(Xd_0__inst_mult_9_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_144 ),
	.cout(Xd_0__inst_mult_9_145 ),
	.shareout(Xd_0__inst_mult_9_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_42 (
// Equation(s):
// Xd_0__inst_mult_6_140  = SUM(( (!din_a[47] & (((din_a[46] & din_b[46])))) # (din_a[47] & (!din_b[45] $ (((!din_a[46]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_6_134  ) + ( Xd_0__inst_mult_6_133  ))
// Xd_0__inst_mult_6_141  = CARRY(( (!din_a[47] & (((din_a[46] & din_b[46])))) # (din_a[47] & (!din_b[45] $ (((!din_a[46]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_6_134  ) + ( Xd_0__inst_mult_6_133  ))
// Xd_0__inst_mult_6_142  = SHARE((din_a[47] & (din_b[45] & (din_a[46] & din_b[46]))))

	.dataa(!din_a[47]),
	.datab(!din_b[45]),
	.datac(!din_a[46]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_133 ),
	.sharein(Xd_0__inst_mult_6_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_140 ),
	.cout(Xd_0__inst_mult_6_141 ),
	.shareout(Xd_0__inst_mult_6_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_43 (
// Equation(s):
// Xd_0__inst_mult_6_144  = SUM(( (din_a[45] & din_b[47]) ) + ( Xd_0__inst_mult_6_138  ) + ( Xd_0__inst_mult_6_137  ))
// Xd_0__inst_mult_6_145  = CARRY(( (din_a[45] & din_b[47]) ) + ( Xd_0__inst_mult_6_138  ) + ( Xd_0__inst_mult_6_137  ))
// Xd_0__inst_mult_6_146  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_137 ),
	.sharein(Xd_0__inst_mult_6_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_144 ),
	.cout(Xd_0__inst_mult_6_145 ),
	.shareout(Xd_0__inst_mult_6_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_42 (
// Equation(s):
// Xd_0__inst_mult_7_140  = SUM(( (!din_a[54] & (((din_a[53] & din_b[53])))) # (din_a[54] & (!din_b[52] $ (((!din_a[53]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_7_134  ) + ( Xd_0__inst_mult_7_133  ))
// Xd_0__inst_mult_7_141  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[53])))) # (din_a[54] & (!din_b[52] $ (((!din_a[53]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_7_134  ) + ( Xd_0__inst_mult_7_133  ))
// Xd_0__inst_mult_7_142  = SHARE((din_a[54] & (din_b[52] & (din_a[53] & din_b[53]))))

	.dataa(!din_a[54]),
	.datab(!din_b[52]),
	.datac(!din_a[53]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_133 ),
	.sharein(Xd_0__inst_mult_7_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_140 ),
	.cout(Xd_0__inst_mult_7_141 ),
	.shareout(Xd_0__inst_mult_7_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_43 (
// Equation(s):
// Xd_0__inst_mult_7_144  = SUM(( (din_a[52] & din_b[54]) ) + ( Xd_0__inst_mult_7_138  ) + ( Xd_0__inst_mult_7_137  ))
// Xd_0__inst_mult_7_145  = CARRY(( (din_a[52] & din_b[54]) ) + ( Xd_0__inst_mult_7_138  ) + ( Xd_0__inst_mult_7_137  ))
// Xd_0__inst_mult_7_146  = SHARE(GND)

	.dataa(!din_a[52]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_137 ),
	.sharein(Xd_0__inst_mult_7_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_144 ),
	.cout(Xd_0__inst_mult_7_145 ),
	.shareout(Xd_0__inst_mult_7_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_42 (
// Equation(s):
// Xd_0__inst_mult_4_140  = SUM(( (!din_a[33] & (((din_a[32] & din_b[32])))) # (din_a[33] & (!din_b[31] $ (((!din_a[32]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_4_134  ) + ( Xd_0__inst_mult_4_133  ))
// Xd_0__inst_mult_4_141  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[32])))) # (din_a[33] & (!din_b[31] $ (((!din_a[32]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_4_134  ) + ( Xd_0__inst_mult_4_133  ))
// Xd_0__inst_mult_4_142  = SHARE((din_a[33] & (din_b[31] & (din_a[32] & din_b[32]))))

	.dataa(!din_a[33]),
	.datab(!din_b[31]),
	.datac(!din_a[32]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_133 ),
	.sharein(Xd_0__inst_mult_4_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_140 ),
	.cout(Xd_0__inst_mult_4_141 ),
	.shareout(Xd_0__inst_mult_4_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_43 (
// Equation(s):
// Xd_0__inst_mult_4_144  = SUM(( (din_a[31] & din_b[33]) ) + ( Xd_0__inst_mult_4_138  ) + ( Xd_0__inst_mult_4_137  ))
// Xd_0__inst_mult_4_145  = CARRY(( (din_a[31] & din_b[33]) ) + ( Xd_0__inst_mult_4_138  ) + ( Xd_0__inst_mult_4_137  ))
// Xd_0__inst_mult_4_146  = SHARE(GND)

	.dataa(!din_a[31]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_137 ),
	.sharein(Xd_0__inst_mult_4_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_144 ),
	.cout(Xd_0__inst_mult_4_145 ),
	.shareout(Xd_0__inst_mult_4_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_42 (
// Equation(s):
// Xd_0__inst_mult_5_140  = SUM(( (!din_a[40] & (((din_a[39] & din_b[39])))) # (din_a[40] & (!din_b[38] $ (((!din_a[39]) # (!din_b[39]))))) ) + ( Xd_0__inst_mult_5_134  ) + ( Xd_0__inst_mult_5_133  ))
// Xd_0__inst_mult_5_141  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[39])))) # (din_a[40] & (!din_b[38] $ (((!din_a[39]) # (!din_b[39]))))) ) + ( Xd_0__inst_mult_5_134  ) + ( Xd_0__inst_mult_5_133  ))
// Xd_0__inst_mult_5_142  = SHARE((din_a[40] & (din_b[38] & (din_a[39] & din_b[39]))))

	.dataa(!din_a[40]),
	.datab(!din_b[38]),
	.datac(!din_a[39]),
	.datad(!din_b[39]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_133 ),
	.sharein(Xd_0__inst_mult_5_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_140 ),
	.cout(Xd_0__inst_mult_5_141 ),
	.shareout(Xd_0__inst_mult_5_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_43 (
// Equation(s):
// Xd_0__inst_mult_5_144  = SUM(( (din_a[38] & din_b[40]) ) + ( Xd_0__inst_mult_5_138  ) + ( Xd_0__inst_mult_5_137  ))
// Xd_0__inst_mult_5_145  = CARRY(( (din_a[38] & din_b[40]) ) + ( Xd_0__inst_mult_5_138  ) + ( Xd_0__inst_mult_5_137  ))
// Xd_0__inst_mult_5_146  = SHARE(GND)

	.dataa(!din_a[38]),
	.datab(!din_b[40]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_137 ),
	.sharein(Xd_0__inst_mult_5_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_144 ),
	.cout(Xd_0__inst_mult_5_145 ),
	.shareout(Xd_0__inst_mult_5_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_42 (
// Equation(s):
// Xd_0__inst_mult_2_140  = SUM(( (!din_a[19] & (((din_a[18] & din_b[18])))) # (din_a[19] & (!din_b[17] $ (((!din_a[18]) # (!din_b[18]))))) ) + ( Xd_0__inst_mult_2_134  ) + ( Xd_0__inst_mult_2_133  ))
// Xd_0__inst_mult_2_141  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[18])))) # (din_a[19] & (!din_b[17] $ (((!din_a[18]) # (!din_b[18]))))) ) + ( Xd_0__inst_mult_2_134  ) + ( Xd_0__inst_mult_2_133  ))
// Xd_0__inst_mult_2_142  = SHARE((din_a[19] & (din_b[17] & (din_a[18] & din_b[18]))))

	.dataa(!din_a[19]),
	.datab(!din_b[17]),
	.datac(!din_a[18]),
	.datad(!din_b[18]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_133 ),
	.sharein(Xd_0__inst_mult_2_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_140 ),
	.cout(Xd_0__inst_mult_2_141 ),
	.shareout(Xd_0__inst_mult_2_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_43 (
// Equation(s):
// Xd_0__inst_mult_2_144  = SUM(( (din_a[17] & din_b[19]) ) + ( Xd_0__inst_mult_2_138  ) + ( Xd_0__inst_mult_2_137  ))
// Xd_0__inst_mult_2_145  = CARRY(( (din_a[17] & din_b[19]) ) + ( Xd_0__inst_mult_2_138  ) + ( Xd_0__inst_mult_2_137  ))
// Xd_0__inst_mult_2_146  = SHARE(GND)

	.dataa(!din_a[17]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_137 ),
	.sharein(Xd_0__inst_mult_2_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_144 ),
	.cout(Xd_0__inst_mult_2_145 ),
	.shareout(Xd_0__inst_mult_2_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_42 (
// Equation(s):
// Xd_0__inst_mult_3_140  = SUM(( (!din_a[26] & (((din_a[25] & din_b[25])))) # (din_a[26] & (!din_b[24] $ (((!din_a[25]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_3_134  ) + ( Xd_0__inst_mult_3_133  ))
// Xd_0__inst_mult_3_141  = CARRY(( (!din_a[26] & (((din_a[25] & din_b[25])))) # (din_a[26] & (!din_b[24] $ (((!din_a[25]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_3_134  ) + ( Xd_0__inst_mult_3_133  ))
// Xd_0__inst_mult_3_142  = SHARE((din_a[26] & (din_b[24] & (din_a[25] & din_b[25]))))

	.dataa(!din_a[26]),
	.datab(!din_b[24]),
	.datac(!din_a[25]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_133 ),
	.sharein(Xd_0__inst_mult_3_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_140 ),
	.cout(Xd_0__inst_mult_3_141 ),
	.shareout(Xd_0__inst_mult_3_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_43 (
// Equation(s):
// Xd_0__inst_mult_3_144  = SUM(( (din_a[24] & din_b[26]) ) + ( Xd_0__inst_mult_3_138  ) + ( Xd_0__inst_mult_3_137  ))
// Xd_0__inst_mult_3_145  = CARRY(( (din_a[24] & din_b[26]) ) + ( Xd_0__inst_mult_3_138  ) + ( Xd_0__inst_mult_3_137  ))
// Xd_0__inst_mult_3_146  = SHARE(GND)

	.dataa(!din_a[24]),
	.datab(!din_b[26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_137 ),
	.sharein(Xd_0__inst_mult_3_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_144 ),
	.cout(Xd_0__inst_mult_3_145 ),
	.shareout(Xd_0__inst_mult_3_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_42 (
// Equation(s):
// Xd_0__inst_mult_0_140  = SUM(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_134  ) + ( Xd_0__inst_mult_0_133  ))
// Xd_0__inst_mult_0_141  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_134  ) + ( Xd_0__inst_mult_0_133  ))
// Xd_0__inst_mult_0_142  = SHARE((din_a[5] & (din_b[3] & (din_a[4] & din_b[4]))))

	.dataa(!din_a[5]),
	.datab(!din_b[3]),
	.datac(!din_a[4]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_133 ),
	.sharein(Xd_0__inst_mult_0_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_140 ),
	.cout(Xd_0__inst_mult_0_141 ),
	.shareout(Xd_0__inst_mult_0_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_43 (
// Equation(s):
// Xd_0__inst_mult_0_144  = SUM(( (din_a[3] & din_b[5]) ) + ( Xd_0__inst_mult_0_138  ) + ( Xd_0__inst_mult_0_137  ))
// Xd_0__inst_mult_0_145  = CARRY(( (din_a[3] & din_b[5]) ) + ( Xd_0__inst_mult_0_138  ) + ( Xd_0__inst_mult_0_137  ))
// Xd_0__inst_mult_0_146  = SHARE(GND)

	.dataa(!din_a[3]),
	.datab(!din_b[5]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_137 ),
	.sharein(Xd_0__inst_mult_0_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_144 ),
	.cout(Xd_0__inst_mult_0_145 ),
	.shareout(Xd_0__inst_mult_0_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_42 (
// Equation(s):
// Xd_0__inst_mult_1_140  = SUM(( (!din_a[12] & (((din_a[11] & din_b[11])))) # (din_a[12] & (!din_b[10] $ (((!din_a[11]) # (!din_b[11]))))) ) + ( Xd_0__inst_mult_1_134  ) + ( Xd_0__inst_mult_1_133  ))
// Xd_0__inst_mult_1_141  = CARRY(( (!din_a[12] & (((din_a[11] & din_b[11])))) # (din_a[12] & (!din_b[10] $ (((!din_a[11]) # (!din_b[11]))))) ) + ( Xd_0__inst_mult_1_134  ) + ( Xd_0__inst_mult_1_133  ))
// Xd_0__inst_mult_1_142  = SHARE((din_a[12] & (din_b[10] & (din_a[11] & din_b[11]))))

	.dataa(!din_a[12]),
	.datab(!din_b[10]),
	.datac(!din_a[11]),
	.datad(!din_b[11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_133 ),
	.sharein(Xd_0__inst_mult_1_134 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_140 ),
	.cout(Xd_0__inst_mult_1_141 ),
	.shareout(Xd_0__inst_mult_1_142 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_43 (
// Equation(s):
// Xd_0__inst_mult_1_144  = SUM(( (din_a[10] & din_b[12]) ) + ( Xd_0__inst_mult_1_138  ) + ( Xd_0__inst_mult_1_137  ))
// Xd_0__inst_mult_1_145  = CARRY(( (din_a[10] & din_b[12]) ) + ( Xd_0__inst_mult_1_138  ) + ( Xd_0__inst_mult_1_137  ))
// Xd_0__inst_mult_1_146  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_137 ),
	.sharein(Xd_0__inst_mult_1_138 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_144 ),
	.cout(Xd_0__inst_mult_1_145 ),
	.shareout(Xd_0__inst_mult_1_146 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_44 (
// Equation(s):
// Xd_0__inst_mult_28_148  = SUM(( (din_a[201] & din_b[200]) ) + ( Xd_0__inst_mult_28_142  ) + ( Xd_0__inst_mult_28_141  ))
// Xd_0__inst_mult_28_149  = CARRY(( (din_a[201] & din_b[200]) ) + ( Xd_0__inst_mult_28_142  ) + ( Xd_0__inst_mult_28_141  ))
// Xd_0__inst_mult_28_150  = SHARE(GND)

	.dataa(!din_a[201]),
	.datab(!din_b[200]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_141 ),
	.sharein(Xd_0__inst_mult_28_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_148 ),
	.cout(Xd_0__inst_mult_28_149 ),
	.shareout(Xd_0__inst_mult_28_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_44 (
// Equation(s):
// Xd_0__inst_mult_29_148  = SUM(( (din_a[208] & din_b[207]) ) + ( Xd_0__inst_mult_29_142  ) + ( Xd_0__inst_mult_29_141  ))
// Xd_0__inst_mult_29_149  = CARRY(( (din_a[208] & din_b[207]) ) + ( Xd_0__inst_mult_29_142  ) + ( Xd_0__inst_mult_29_141  ))
// Xd_0__inst_mult_29_150  = SHARE(GND)

	.dataa(!din_a[208]),
	.datab(!din_b[207]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_141 ),
	.sharein(Xd_0__inst_mult_29_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_148 ),
	.cout(Xd_0__inst_mult_29_149 ),
	.shareout(Xd_0__inst_mult_29_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_44 (
// Equation(s):
// Xd_0__inst_mult_26_148  = SUM(( (din_a[187] & din_b[186]) ) + ( Xd_0__inst_mult_26_142  ) + ( Xd_0__inst_mult_26_141  ))
// Xd_0__inst_mult_26_149  = CARRY(( (din_a[187] & din_b[186]) ) + ( Xd_0__inst_mult_26_142  ) + ( Xd_0__inst_mult_26_141  ))
// Xd_0__inst_mult_26_150  = SHARE(GND)

	.dataa(!din_a[187]),
	.datab(!din_b[186]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_141 ),
	.sharein(Xd_0__inst_mult_26_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_148 ),
	.cout(Xd_0__inst_mult_26_149 ),
	.shareout(Xd_0__inst_mult_26_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_44 (
// Equation(s):
// Xd_0__inst_mult_27_148  = SUM(( (din_a[194] & din_b[193]) ) + ( Xd_0__inst_mult_27_142  ) + ( Xd_0__inst_mult_27_141  ))
// Xd_0__inst_mult_27_149  = CARRY(( (din_a[194] & din_b[193]) ) + ( Xd_0__inst_mult_27_142  ) + ( Xd_0__inst_mult_27_141  ))
// Xd_0__inst_mult_27_150  = SHARE(GND)

	.dataa(!din_a[194]),
	.datab(!din_b[193]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_141 ),
	.sharein(Xd_0__inst_mult_27_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_148 ),
	.cout(Xd_0__inst_mult_27_149 ),
	.shareout(Xd_0__inst_mult_27_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_44 (
// Equation(s):
// Xd_0__inst_mult_24_148  = SUM(( (din_a[173] & din_b[172]) ) + ( Xd_0__inst_mult_24_142  ) + ( Xd_0__inst_mult_24_141  ))
// Xd_0__inst_mult_24_149  = CARRY(( (din_a[173] & din_b[172]) ) + ( Xd_0__inst_mult_24_142  ) + ( Xd_0__inst_mult_24_141  ))
// Xd_0__inst_mult_24_150  = SHARE(GND)

	.dataa(!din_a[173]),
	.datab(!din_b[172]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_141 ),
	.sharein(Xd_0__inst_mult_24_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_148 ),
	.cout(Xd_0__inst_mult_24_149 ),
	.shareout(Xd_0__inst_mult_24_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_44 (
// Equation(s):
// Xd_0__inst_mult_25_148  = SUM(( (din_a[180] & din_b[179]) ) + ( Xd_0__inst_mult_25_146  ) + ( Xd_0__inst_mult_25_145  ))
// Xd_0__inst_mult_25_149  = CARRY(( (din_a[180] & din_b[179]) ) + ( Xd_0__inst_mult_25_146  ) + ( Xd_0__inst_mult_25_145  ))
// Xd_0__inst_mult_25_150  = SHARE(GND)

	.dataa(!din_a[180]),
	.datab(!din_b[179]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_145 ),
	.sharein(Xd_0__inst_mult_25_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_148 ),
	.cout(Xd_0__inst_mult_25_149 ),
	.shareout(Xd_0__inst_mult_25_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_44 (
// Equation(s):
// Xd_0__inst_mult_22_148  = SUM(( (din_a[159] & din_b[158]) ) + ( Xd_0__inst_mult_22_146  ) + ( Xd_0__inst_mult_22_145  ))
// Xd_0__inst_mult_22_149  = CARRY(( (din_a[159] & din_b[158]) ) + ( Xd_0__inst_mult_22_146  ) + ( Xd_0__inst_mult_22_145  ))
// Xd_0__inst_mult_22_150  = SHARE(GND)

	.dataa(!din_a[159]),
	.datab(!din_b[158]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_145 ),
	.sharein(Xd_0__inst_mult_22_146 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_148 ),
	.cout(Xd_0__inst_mult_22_149 ),
	.shareout(Xd_0__inst_mult_22_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_44 (
// Equation(s):
// Xd_0__inst_mult_23_148  = SUM(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_23_142  ) + ( Xd_0__inst_mult_23_141  ))
// Xd_0__inst_mult_23_149  = CARRY(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_23_142  ) + ( Xd_0__inst_mult_23_141  ))
// Xd_0__inst_mult_23_150  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_141 ),
	.sharein(Xd_0__inst_mult_23_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_148 ),
	.cout(Xd_0__inst_mult_23_149 ),
	.shareout(Xd_0__inst_mult_23_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_44 (
// Equation(s):
// Xd_0__inst_mult_20_148  = SUM(( (din_a[145] & din_b[144]) ) + ( Xd_0__inst_mult_20_142  ) + ( Xd_0__inst_mult_20_141  ))
// Xd_0__inst_mult_20_149  = CARRY(( (din_a[145] & din_b[144]) ) + ( Xd_0__inst_mult_20_142  ) + ( Xd_0__inst_mult_20_141  ))
// Xd_0__inst_mult_20_150  = SHARE(GND)

	.dataa(!din_a[145]),
	.datab(!din_b[144]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_141 ),
	.sharein(Xd_0__inst_mult_20_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_148 ),
	.cout(Xd_0__inst_mult_20_149 ),
	.shareout(Xd_0__inst_mult_20_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_44 (
// Equation(s):
// Xd_0__inst_mult_21_148  = SUM(( (din_a[152] & din_b[151]) ) + ( Xd_0__inst_mult_21_142  ) + ( Xd_0__inst_mult_21_141  ))
// Xd_0__inst_mult_21_149  = CARRY(( (din_a[152] & din_b[151]) ) + ( Xd_0__inst_mult_21_142  ) + ( Xd_0__inst_mult_21_141  ))
// Xd_0__inst_mult_21_150  = SHARE(GND)

	.dataa(!din_a[152]),
	.datab(!din_b[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_141 ),
	.sharein(Xd_0__inst_mult_21_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_148 ),
	.cout(Xd_0__inst_mult_21_149 ),
	.shareout(Xd_0__inst_mult_21_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_44 (
// Equation(s):
// Xd_0__inst_mult_18_148  = SUM(( (din_a[131] & din_b[130]) ) + ( Xd_0__inst_mult_18_142  ) + ( Xd_0__inst_mult_18_141  ))
// Xd_0__inst_mult_18_149  = CARRY(( (din_a[131] & din_b[130]) ) + ( Xd_0__inst_mult_18_142  ) + ( Xd_0__inst_mult_18_141  ))
// Xd_0__inst_mult_18_150  = SHARE(GND)

	.dataa(!din_a[131]),
	.datab(!din_b[130]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_141 ),
	.sharein(Xd_0__inst_mult_18_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_148 ),
	.cout(Xd_0__inst_mult_18_149 ),
	.shareout(Xd_0__inst_mult_18_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_44 (
// Equation(s):
// Xd_0__inst_mult_19_148  = SUM(( (din_a[138] & din_b[137]) ) + ( Xd_0__inst_mult_19_142  ) + ( Xd_0__inst_mult_19_141  ))
// Xd_0__inst_mult_19_149  = CARRY(( (din_a[138] & din_b[137]) ) + ( Xd_0__inst_mult_19_142  ) + ( Xd_0__inst_mult_19_141  ))
// Xd_0__inst_mult_19_150  = SHARE(GND)

	.dataa(!din_a[138]),
	.datab(!din_b[137]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_141 ),
	.sharein(Xd_0__inst_mult_19_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_148 ),
	.cout(Xd_0__inst_mult_19_149 ),
	.shareout(Xd_0__inst_mult_19_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_44 (
// Equation(s):
// Xd_0__inst_mult_16_148  = SUM(( (din_a[117] & din_b[116]) ) + ( Xd_0__inst_mult_16_142  ) + ( Xd_0__inst_mult_16_141  ))
// Xd_0__inst_mult_16_149  = CARRY(( (din_a[117] & din_b[116]) ) + ( Xd_0__inst_mult_16_142  ) + ( Xd_0__inst_mult_16_141  ))
// Xd_0__inst_mult_16_150  = SHARE(GND)

	.dataa(!din_a[117]),
	.datab(!din_b[116]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_141 ),
	.sharein(Xd_0__inst_mult_16_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_148 ),
	.cout(Xd_0__inst_mult_16_149 ),
	.shareout(Xd_0__inst_mult_16_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_44 (
// Equation(s):
// Xd_0__inst_mult_17_148  = SUM(( (din_a[124] & din_b[123]) ) + ( Xd_0__inst_mult_17_142  ) + ( Xd_0__inst_mult_17_141  ))
// Xd_0__inst_mult_17_149  = CARRY(( (din_a[124] & din_b[123]) ) + ( Xd_0__inst_mult_17_142  ) + ( Xd_0__inst_mult_17_141  ))
// Xd_0__inst_mult_17_150  = SHARE(GND)

	.dataa(!din_a[124]),
	.datab(!din_b[123]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_141 ),
	.sharein(Xd_0__inst_mult_17_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_148 ),
	.cout(Xd_0__inst_mult_17_149 ),
	.shareout(Xd_0__inst_mult_17_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_44 (
// Equation(s):
// Xd_0__inst_mult_14_148  = SUM(( (din_a[103] & din_b[102]) ) + ( Xd_0__inst_mult_14_142  ) + ( Xd_0__inst_mult_14_141  ))
// Xd_0__inst_mult_14_149  = CARRY(( (din_a[103] & din_b[102]) ) + ( Xd_0__inst_mult_14_142  ) + ( Xd_0__inst_mult_14_141  ))
// Xd_0__inst_mult_14_150  = SHARE(GND)

	.dataa(!din_a[103]),
	.datab(!din_b[102]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_141 ),
	.sharein(Xd_0__inst_mult_14_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_148 ),
	.cout(Xd_0__inst_mult_14_149 ),
	.shareout(Xd_0__inst_mult_14_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_44 (
// Equation(s):
// Xd_0__inst_mult_15_148  = SUM(( (din_a[110] & din_b[109]) ) + ( Xd_0__inst_mult_15_142  ) + ( Xd_0__inst_mult_15_141  ))
// Xd_0__inst_mult_15_149  = CARRY(( (din_a[110] & din_b[109]) ) + ( Xd_0__inst_mult_15_142  ) + ( Xd_0__inst_mult_15_141  ))
// Xd_0__inst_mult_15_150  = SHARE(GND)

	.dataa(!din_a[110]),
	.datab(!din_b[109]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_141 ),
	.sharein(Xd_0__inst_mult_15_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_148 ),
	.cout(Xd_0__inst_mult_15_149 ),
	.shareout(Xd_0__inst_mult_15_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_44 (
// Equation(s):
// Xd_0__inst_mult_12_148  = SUM(( (din_a[89] & din_b[88]) ) + ( Xd_0__inst_mult_12_142  ) + ( Xd_0__inst_mult_12_141  ))
// Xd_0__inst_mult_12_149  = CARRY(( (din_a[89] & din_b[88]) ) + ( Xd_0__inst_mult_12_142  ) + ( Xd_0__inst_mult_12_141  ))
// Xd_0__inst_mult_12_150  = SHARE(GND)

	.dataa(!din_a[89]),
	.datab(!din_b[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_141 ),
	.sharein(Xd_0__inst_mult_12_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_148 ),
	.cout(Xd_0__inst_mult_12_149 ),
	.shareout(Xd_0__inst_mult_12_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_44 (
// Equation(s):
// Xd_0__inst_mult_13_148  = SUM(( (din_a[96] & din_b[95]) ) + ( Xd_0__inst_mult_13_142  ) + ( Xd_0__inst_mult_13_141  ))
// Xd_0__inst_mult_13_149  = CARRY(( (din_a[96] & din_b[95]) ) + ( Xd_0__inst_mult_13_142  ) + ( Xd_0__inst_mult_13_141  ))
// Xd_0__inst_mult_13_150  = SHARE(GND)

	.dataa(!din_a[96]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_141 ),
	.sharein(Xd_0__inst_mult_13_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_148 ),
	.cout(Xd_0__inst_mult_13_149 ),
	.shareout(Xd_0__inst_mult_13_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_44 (
// Equation(s):
// Xd_0__inst_mult_10_148  = SUM(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_10_142  ) + ( Xd_0__inst_mult_10_141  ))
// Xd_0__inst_mult_10_149  = CARRY(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_10_142  ) + ( Xd_0__inst_mult_10_141  ))
// Xd_0__inst_mult_10_150  = SHARE(GND)

	.dataa(!din_a[75]),
	.datab(!din_b[74]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_141 ),
	.sharein(Xd_0__inst_mult_10_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_148 ),
	.cout(Xd_0__inst_mult_10_149 ),
	.shareout(Xd_0__inst_mult_10_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_44 (
// Equation(s):
// Xd_0__inst_mult_11_148  = SUM(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_11_142  ) + ( Xd_0__inst_mult_11_141  ))
// Xd_0__inst_mult_11_149  = CARRY(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_11_142  ) + ( Xd_0__inst_mult_11_141  ))
// Xd_0__inst_mult_11_150  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_141 ),
	.sharein(Xd_0__inst_mult_11_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_148 ),
	.cout(Xd_0__inst_mult_11_149 ),
	.shareout(Xd_0__inst_mult_11_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_44 (
// Equation(s):
// Xd_0__inst_mult_8_148  = SUM(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_8_142  ) + ( Xd_0__inst_mult_8_141  ))
// Xd_0__inst_mult_8_149  = CARRY(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_8_142  ) + ( Xd_0__inst_mult_8_141  ))
// Xd_0__inst_mult_8_150  = SHARE(GND)

	.dataa(!din_a[61]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_141 ),
	.sharein(Xd_0__inst_mult_8_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_148 ),
	.cout(Xd_0__inst_mult_8_149 ),
	.shareout(Xd_0__inst_mult_8_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_44 (
// Equation(s):
// Xd_0__inst_mult_9_148  = SUM(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_9_142  ) + ( Xd_0__inst_mult_9_141  ))
// Xd_0__inst_mult_9_149  = CARRY(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_9_142  ) + ( Xd_0__inst_mult_9_141  ))
// Xd_0__inst_mult_9_150  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_141 ),
	.sharein(Xd_0__inst_mult_9_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_148 ),
	.cout(Xd_0__inst_mult_9_149 ),
	.shareout(Xd_0__inst_mult_9_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_44 (
// Equation(s):
// Xd_0__inst_mult_6_148  = SUM(( (din_a[47] & din_b[46]) ) + ( Xd_0__inst_mult_6_142  ) + ( Xd_0__inst_mult_6_141  ))
// Xd_0__inst_mult_6_149  = CARRY(( (din_a[47] & din_b[46]) ) + ( Xd_0__inst_mult_6_142  ) + ( Xd_0__inst_mult_6_141  ))
// Xd_0__inst_mult_6_150  = SHARE(GND)

	.dataa(!din_a[47]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_141 ),
	.sharein(Xd_0__inst_mult_6_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_148 ),
	.cout(Xd_0__inst_mult_6_149 ),
	.shareout(Xd_0__inst_mult_6_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_44 (
// Equation(s):
// Xd_0__inst_mult_7_148  = SUM(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_7_142  ) + ( Xd_0__inst_mult_7_141  ))
// Xd_0__inst_mult_7_149  = CARRY(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_7_142  ) + ( Xd_0__inst_mult_7_141  ))
// Xd_0__inst_mult_7_150  = SHARE(GND)

	.dataa(!din_a[54]),
	.datab(!din_b[53]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_141 ),
	.sharein(Xd_0__inst_mult_7_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_148 ),
	.cout(Xd_0__inst_mult_7_149 ),
	.shareout(Xd_0__inst_mult_7_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_44 (
// Equation(s):
// Xd_0__inst_mult_4_148  = SUM(( (din_a[33] & din_b[32]) ) + ( Xd_0__inst_mult_4_142  ) + ( Xd_0__inst_mult_4_141  ))
// Xd_0__inst_mult_4_149  = CARRY(( (din_a[33] & din_b[32]) ) + ( Xd_0__inst_mult_4_142  ) + ( Xd_0__inst_mult_4_141  ))
// Xd_0__inst_mult_4_150  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_141 ),
	.sharein(Xd_0__inst_mult_4_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_148 ),
	.cout(Xd_0__inst_mult_4_149 ),
	.shareout(Xd_0__inst_mult_4_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_44 (
// Equation(s):
// Xd_0__inst_mult_5_148  = SUM(( (din_a[40] & din_b[39]) ) + ( Xd_0__inst_mult_5_142  ) + ( Xd_0__inst_mult_5_141  ))
// Xd_0__inst_mult_5_149  = CARRY(( (din_a[40] & din_b[39]) ) + ( Xd_0__inst_mult_5_142  ) + ( Xd_0__inst_mult_5_141  ))
// Xd_0__inst_mult_5_150  = SHARE(GND)

	.dataa(!din_a[40]),
	.datab(!din_b[39]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_141 ),
	.sharein(Xd_0__inst_mult_5_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_148 ),
	.cout(Xd_0__inst_mult_5_149 ),
	.shareout(Xd_0__inst_mult_5_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_44 (
// Equation(s):
// Xd_0__inst_mult_2_148  = SUM(( (din_a[19] & din_b[18]) ) + ( Xd_0__inst_mult_2_142  ) + ( Xd_0__inst_mult_2_141  ))
// Xd_0__inst_mult_2_149  = CARRY(( (din_a[19] & din_b[18]) ) + ( Xd_0__inst_mult_2_142  ) + ( Xd_0__inst_mult_2_141  ))
// Xd_0__inst_mult_2_150  = SHARE(GND)

	.dataa(!din_a[19]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_141 ),
	.sharein(Xd_0__inst_mult_2_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_148 ),
	.cout(Xd_0__inst_mult_2_149 ),
	.shareout(Xd_0__inst_mult_2_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_44 (
// Equation(s):
// Xd_0__inst_mult_3_148  = SUM(( (din_a[26] & din_b[25]) ) + ( Xd_0__inst_mult_3_142  ) + ( Xd_0__inst_mult_3_141  ))
// Xd_0__inst_mult_3_149  = CARRY(( (din_a[26] & din_b[25]) ) + ( Xd_0__inst_mult_3_142  ) + ( Xd_0__inst_mult_3_141  ))
// Xd_0__inst_mult_3_150  = SHARE(GND)

	.dataa(!din_a[26]),
	.datab(!din_b[25]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_141 ),
	.sharein(Xd_0__inst_mult_3_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_148 ),
	.cout(Xd_0__inst_mult_3_149 ),
	.shareout(Xd_0__inst_mult_3_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_44 (
// Equation(s):
// Xd_0__inst_mult_0_148  = SUM(( (din_a[5] & din_b[4]) ) + ( Xd_0__inst_mult_0_142  ) + ( Xd_0__inst_mult_0_141  ))
// Xd_0__inst_mult_0_149  = CARRY(( (din_a[5] & din_b[4]) ) + ( Xd_0__inst_mult_0_142  ) + ( Xd_0__inst_mult_0_141  ))
// Xd_0__inst_mult_0_150  = SHARE(GND)

	.dataa(!din_a[5]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_141 ),
	.sharein(Xd_0__inst_mult_0_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_148 ),
	.cout(Xd_0__inst_mult_0_149 ),
	.shareout(Xd_0__inst_mult_0_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_44 (
// Equation(s):
// Xd_0__inst_mult_1_148  = SUM(( (din_a[12] & din_b[11]) ) + ( Xd_0__inst_mult_1_142  ) + ( Xd_0__inst_mult_1_141  ))
// Xd_0__inst_mult_1_149  = CARRY(( (din_a[12] & din_b[11]) ) + ( Xd_0__inst_mult_1_142  ) + ( Xd_0__inst_mult_1_141  ))
// Xd_0__inst_mult_1_150  = SHARE(GND)

	.dataa(!din_a[12]),
	.datab(!din_b[11]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_141 ),
	.sharein(Xd_0__inst_mult_1_142 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_148 ),
	.cout(Xd_0__inst_mult_1_149 ),
	.shareout(Xd_0__inst_mult_1_150 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_45 (
// Equation(s):
// Xd_0__inst_mult_28_152  = SUM(( GND ) + ( Xd_0__inst_mult_28_150  ) + ( Xd_0__inst_mult_28_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_149 ),
	.sharein(Xd_0__inst_mult_28_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_45 (
// Equation(s):
// Xd_0__inst_mult_29_152  = SUM(( GND ) + ( Xd_0__inst_mult_29_150  ) + ( Xd_0__inst_mult_29_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_149 ),
	.sharein(Xd_0__inst_mult_29_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_45 (
// Equation(s):
// Xd_0__inst_mult_26_152  = SUM(( GND ) + ( Xd_0__inst_mult_26_150  ) + ( Xd_0__inst_mult_26_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_149 ),
	.sharein(Xd_0__inst_mult_26_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_45 (
// Equation(s):
// Xd_0__inst_mult_27_152  = SUM(( GND ) + ( Xd_0__inst_mult_27_150  ) + ( Xd_0__inst_mult_27_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_149 ),
	.sharein(Xd_0__inst_mult_27_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_45 (
// Equation(s):
// Xd_0__inst_mult_24_152  = SUM(( GND ) + ( Xd_0__inst_mult_24_150  ) + ( Xd_0__inst_mult_24_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_149 ),
	.sharein(Xd_0__inst_mult_24_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_45 (
// Equation(s):
// Xd_0__inst_mult_25_152  = SUM(( GND ) + ( Xd_0__inst_mult_25_150  ) + ( Xd_0__inst_mult_25_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_149 ),
	.sharein(Xd_0__inst_mult_25_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_45 (
// Equation(s):
// Xd_0__inst_mult_22_152  = SUM(( GND ) + ( Xd_0__inst_mult_22_150  ) + ( Xd_0__inst_mult_22_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_149 ),
	.sharein(Xd_0__inst_mult_22_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_45 (
// Equation(s):
// Xd_0__inst_mult_23_152  = SUM(( GND ) + ( Xd_0__inst_mult_23_150  ) + ( Xd_0__inst_mult_23_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_149 ),
	.sharein(Xd_0__inst_mult_23_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_45 (
// Equation(s):
// Xd_0__inst_mult_20_152  = SUM(( GND ) + ( Xd_0__inst_mult_20_150  ) + ( Xd_0__inst_mult_20_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_149 ),
	.sharein(Xd_0__inst_mult_20_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_45 (
// Equation(s):
// Xd_0__inst_mult_21_152  = SUM(( GND ) + ( Xd_0__inst_mult_21_150  ) + ( Xd_0__inst_mult_21_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_149 ),
	.sharein(Xd_0__inst_mult_21_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_45 (
// Equation(s):
// Xd_0__inst_mult_18_152  = SUM(( GND ) + ( Xd_0__inst_mult_18_150  ) + ( Xd_0__inst_mult_18_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_149 ),
	.sharein(Xd_0__inst_mult_18_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_45 (
// Equation(s):
// Xd_0__inst_mult_19_152  = SUM(( GND ) + ( Xd_0__inst_mult_19_150  ) + ( Xd_0__inst_mult_19_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_149 ),
	.sharein(Xd_0__inst_mult_19_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_45 (
// Equation(s):
// Xd_0__inst_mult_16_152  = SUM(( GND ) + ( Xd_0__inst_mult_16_150  ) + ( Xd_0__inst_mult_16_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_149 ),
	.sharein(Xd_0__inst_mult_16_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_45 (
// Equation(s):
// Xd_0__inst_mult_17_152  = SUM(( GND ) + ( Xd_0__inst_mult_17_150  ) + ( Xd_0__inst_mult_17_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_149 ),
	.sharein(Xd_0__inst_mult_17_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_45 (
// Equation(s):
// Xd_0__inst_mult_14_152  = SUM(( GND ) + ( Xd_0__inst_mult_14_150  ) + ( Xd_0__inst_mult_14_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_149 ),
	.sharein(Xd_0__inst_mult_14_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_45 (
// Equation(s):
// Xd_0__inst_mult_15_152  = SUM(( GND ) + ( Xd_0__inst_mult_15_150  ) + ( Xd_0__inst_mult_15_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_149 ),
	.sharein(Xd_0__inst_mult_15_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_45 (
// Equation(s):
// Xd_0__inst_mult_12_152  = SUM(( GND ) + ( Xd_0__inst_mult_12_150  ) + ( Xd_0__inst_mult_12_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_149 ),
	.sharein(Xd_0__inst_mult_12_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_45 (
// Equation(s):
// Xd_0__inst_mult_13_152  = SUM(( GND ) + ( Xd_0__inst_mult_13_150  ) + ( Xd_0__inst_mult_13_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_149 ),
	.sharein(Xd_0__inst_mult_13_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_45 (
// Equation(s):
// Xd_0__inst_mult_10_152  = SUM(( GND ) + ( Xd_0__inst_mult_10_150  ) + ( Xd_0__inst_mult_10_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_149 ),
	.sharein(Xd_0__inst_mult_10_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_45 (
// Equation(s):
// Xd_0__inst_mult_11_152  = SUM(( GND ) + ( Xd_0__inst_mult_11_150  ) + ( Xd_0__inst_mult_11_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_149 ),
	.sharein(Xd_0__inst_mult_11_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_45 (
// Equation(s):
// Xd_0__inst_mult_8_152  = SUM(( GND ) + ( Xd_0__inst_mult_8_150  ) + ( Xd_0__inst_mult_8_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_149 ),
	.sharein(Xd_0__inst_mult_8_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_45 (
// Equation(s):
// Xd_0__inst_mult_9_152  = SUM(( GND ) + ( Xd_0__inst_mult_9_150  ) + ( Xd_0__inst_mult_9_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_149 ),
	.sharein(Xd_0__inst_mult_9_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_45 (
// Equation(s):
// Xd_0__inst_mult_6_152  = SUM(( GND ) + ( Xd_0__inst_mult_6_150  ) + ( Xd_0__inst_mult_6_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_149 ),
	.sharein(Xd_0__inst_mult_6_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_45 (
// Equation(s):
// Xd_0__inst_mult_7_152  = SUM(( GND ) + ( Xd_0__inst_mult_7_150  ) + ( Xd_0__inst_mult_7_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_149 ),
	.sharein(Xd_0__inst_mult_7_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_45 (
// Equation(s):
// Xd_0__inst_mult_4_152  = SUM(( GND ) + ( Xd_0__inst_mult_4_150  ) + ( Xd_0__inst_mult_4_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_149 ),
	.sharein(Xd_0__inst_mult_4_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_45 (
// Equation(s):
// Xd_0__inst_mult_5_152  = SUM(( GND ) + ( Xd_0__inst_mult_5_150  ) + ( Xd_0__inst_mult_5_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_149 ),
	.sharein(Xd_0__inst_mult_5_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_45 (
// Equation(s):
// Xd_0__inst_mult_2_152  = SUM(( GND ) + ( Xd_0__inst_mult_2_150  ) + ( Xd_0__inst_mult_2_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_149 ),
	.sharein(Xd_0__inst_mult_2_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_45 (
// Equation(s):
// Xd_0__inst_mult_3_152  = SUM(( GND ) + ( Xd_0__inst_mult_3_150  ) + ( Xd_0__inst_mult_3_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_149 ),
	.sharein(Xd_0__inst_mult_3_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_45 (
// Equation(s):
// Xd_0__inst_mult_0_152  = SUM(( GND ) + ( Xd_0__inst_mult_0_150  ) + ( Xd_0__inst_mult_0_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_149 ),
	.sharein(Xd_0__inst_mult_0_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_45 (
// Equation(s):
// Xd_0__inst_mult_1_152  = SUM(( GND ) + ( Xd_0__inst_mult_1_150  ) + ( Xd_0__inst_mult_1_149  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_149 ),
	.sharein(Xd_0__inst_mult_1_150 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_152 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_46 (
// Equation(s):
// Xd_0__inst_mult_28_157  = CARRY(( (din_a[198] & din_b[198]) ) + ( Xd_0__inst_mult_28_162  ) + ( Xd_0__inst_mult_28_161  ))
// Xd_0__inst_mult_28_158  = SHARE((din_a[197] & din_b[199]))

	.dataa(!din_a[198]),
	.datab(!din_b[198]),
	.datac(!din_a[197]),
	.datad(!din_b[199]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_161 ),
	.sharein(Xd_0__inst_mult_28_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_157 ),
	.shareout(Xd_0__inst_mult_28_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_46 (
// Equation(s):
// Xd_0__inst_mult_29_157  = CARRY(( (din_a[205] & din_b[205]) ) + ( Xd_0__inst_mult_29_162  ) + ( Xd_0__inst_mult_29_161  ))
// Xd_0__inst_mult_29_158  = SHARE((din_a[204] & din_b[206]))

	.dataa(!din_a[205]),
	.datab(!din_b[205]),
	.datac(!din_a[204]),
	.datad(!din_b[206]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_161 ),
	.sharein(Xd_0__inst_mult_29_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_157 ),
	.shareout(Xd_0__inst_mult_29_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_46 (
// Equation(s):
// Xd_0__inst_mult_26_157  = CARRY(( (din_a[184] & din_b[184]) ) + ( Xd_0__inst_mult_26_162  ) + ( Xd_0__inst_mult_26_161  ))
// Xd_0__inst_mult_26_158  = SHARE((din_a[183] & din_b[185]))

	.dataa(!din_a[184]),
	.datab(!din_b[184]),
	.datac(!din_a[183]),
	.datad(!din_b[185]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_161 ),
	.sharein(Xd_0__inst_mult_26_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_157 ),
	.shareout(Xd_0__inst_mult_26_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_46 (
// Equation(s):
// Xd_0__inst_mult_27_157  = CARRY(( (din_a[191] & din_b[191]) ) + ( Xd_0__inst_mult_27_162  ) + ( Xd_0__inst_mult_27_161  ))
// Xd_0__inst_mult_27_158  = SHARE((din_a[190] & din_b[192]))

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(!din_a[190]),
	.datad(!din_b[192]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_161 ),
	.sharein(Xd_0__inst_mult_27_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_157 ),
	.shareout(Xd_0__inst_mult_27_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_46 (
// Equation(s):
// Xd_0__inst_mult_24_157  = CARRY(( (din_a[170] & din_b[170]) ) + ( Xd_0__inst_mult_24_162  ) + ( Xd_0__inst_mult_24_161  ))
// Xd_0__inst_mult_24_158  = SHARE((din_a[169] & din_b[171]))

	.dataa(!din_a[170]),
	.datab(!din_b[170]),
	.datac(!din_a[169]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_161 ),
	.sharein(Xd_0__inst_mult_24_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_157 ),
	.shareout(Xd_0__inst_mult_24_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_46 (
// Equation(s):
// Xd_0__inst_mult_25_157  = CARRY(( (din_a[177] & din_b[177]) ) + ( Xd_0__inst_mult_25_162  ) + ( Xd_0__inst_mult_25_161  ))
// Xd_0__inst_mult_25_158  = SHARE((din_a[176] & din_b[178]))

	.dataa(!din_a[177]),
	.datab(!din_b[177]),
	.datac(!din_a[176]),
	.datad(!din_b[178]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_161 ),
	.sharein(Xd_0__inst_mult_25_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_157 ),
	.shareout(Xd_0__inst_mult_25_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_46 (
// Equation(s):
// Xd_0__inst_mult_22_157  = CARRY(( (din_a[156] & din_b[156]) ) + ( Xd_0__inst_mult_22_162  ) + ( Xd_0__inst_mult_22_161  ))
// Xd_0__inst_mult_22_158  = SHARE((din_a[155] & din_b[157]))

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(!din_a[155]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_161 ),
	.sharein(Xd_0__inst_mult_22_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_157 ),
	.shareout(Xd_0__inst_mult_22_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_46 (
// Equation(s):
// Xd_0__inst_mult_23_157  = CARRY(( (din_a[163] & din_b[163]) ) + ( Xd_0__inst_mult_23_162  ) + ( Xd_0__inst_mult_23_161  ))
// Xd_0__inst_mult_23_158  = SHARE((din_a[162] & din_b[164]))

	.dataa(!din_a[163]),
	.datab(!din_b[163]),
	.datac(!din_a[162]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_161 ),
	.sharein(Xd_0__inst_mult_23_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_157 ),
	.shareout(Xd_0__inst_mult_23_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_46 (
// Equation(s):
// Xd_0__inst_mult_20_157  = CARRY(( (din_a[142] & din_b[142]) ) + ( Xd_0__inst_mult_20_162  ) + ( Xd_0__inst_mult_20_161  ))
// Xd_0__inst_mult_20_158  = SHARE((din_a[141] & din_b[143]))

	.dataa(!din_a[142]),
	.datab(!din_b[142]),
	.datac(!din_a[141]),
	.datad(!din_b[143]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_161 ),
	.sharein(Xd_0__inst_mult_20_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_157 ),
	.shareout(Xd_0__inst_mult_20_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_46 (
// Equation(s):
// Xd_0__inst_mult_21_157  = CARRY(( (din_a[149] & din_b[149]) ) + ( Xd_0__inst_mult_21_162  ) + ( Xd_0__inst_mult_21_161  ))
// Xd_0__inst_mult_21_158  = SHARE((din_a[148] & din_b[150]))

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(!din_a[148]),
	.datad(!din_b[150]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_161 ),
	.sharein(Xd_0__inst_mult_21_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_157 ),
	.shareout(Xd_0__inst_mult_21_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_46 (
// Equation(s):
// Xd_0__inst_mult_18_157  = CARRY(( (din_a[128] & din_b[128]) ) + ( Xd_0__inst_mult_18_162  ) + ( Xd_0__inst_mult_18_161  ))
// Xd_0__inst_mult_18_158  = SHARE((din_a[127] & din_b[129]))

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(!din_a[127]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_161 ),
	.sharein(Xd_0__inst_mult_18_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_157 ),
	.shareout(Xd_0__inst_mult_18_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_46 (
// Equation(s):
// Xd_0__inst_mult_19_157  = CARRY(( (din_a[135] & din_b[135]) ) + ( Xd_0__inst_mult_19_162  ) + ( Xd_0__inst_mult_19_161  ))
// Xd_0__inst_mult_19_158  = SHARE((din_a[134] & din_b[136]))

	.dataa(!din_a[135]),
	.datab(!din_b[135]),
	.datac(!din_a[134]),
	.datad(!din_b[136]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_161 ),
	.sharein(Xd_0__inst_mult_19_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_157 ),
	.shareout(Xd_0__inst_mult_19_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_47 (
// Equation(s):
// Xd_0__inst_mult_30_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_30_162  = SHARE((din_a[212] & din_b[212]))

	.dataa(!din_a[212]),
	.datab(!din_b[212]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_161 ),
	.shareout(Xd_0__inst_mult_30_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_47 (
// Equation(s):
// Xd_0__inst_mult_31_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_31_162  = SHARE((din_a[219] & din_b[219]))

	.dataa(!din_a[219]),
	.datab(!din_b[219]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_161 ),
	.shareout(Xd_0__inst_mult_31_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_46 (
// Equation(s):
// Xd_0__inst_mult_16_157  = CARRY(( (din_a[114] & din_b[114]) ) + ( Xd_0__inst_mult_16_162  ) + ( Xd_0__inst_mult_16_161  ))
// Xd_0__inst_mult_16_158  = SHARE((din_a[113] & din_b[115]))

	.dataa(!din_a[114]),
	.datab(!din_b[114]),
	.datac(!din_a[113]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_161 ),
	.sharein(Xd_0__inst_mult_16_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_157 ),
	.shareout(Xd_0__inst_mult_16_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_46 (
// Equation(s):
// Xd_0__inst_mult_17_157  = CARRY(( (din_a[121] & din_b[121]) ) + ( Xd_0__inst_mult_17_162  ) + ( Xd_0__inst_mult_17_161  ))
// Xd_0__inst_mult_17_158  = SHARE((din_a[120] & din_b[122]))

	.dataa(!din_a[121]),
	.datab(!din_b[121]),
	.datac(!din_a[120]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_161 ),
	.sharein(Xd_0__inst_mult_17_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_157 ),
	.shareout(Xd_0__inst_mult_17_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_46 (
// Equation(s):
// Xd_0__inst_mult_14_157  = CARRY(( (din_a[100] & din_b[100]) ) + ( Xd_0__inst_mult_14_162  ) + ( Xd_0__inst_mult_14_161  ))
// Xd_0__inst_mult_14_158  = SHARE((din_a[99] & din_b[101]))

	.dataa(!din_a[100]),
	.datab(!din_b[100]),
	.datac(!din_a[99]),
	.datad(!din_b[101]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_161 ),
	.sharein(Xd_0__inst_mult_14_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_157 ),
	.shareout(Xd_0__inst_mult_14_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_46 (
// Equation(s):
// Xd_0__inst_mult_15_157  = CARRY(( (din_a[107] & din_b[107]) ) + ( Xd_0__inst_mult_15_162  ) + ( Xd_0__inst_mult_15_161  ))
// Xd_0__inst_mult_15_158  = SHARE((din_a[106] & din_b[108]))

	.dataa(!din_a[107]),
	.datab(!din_b[107]),
	.datac(!din_a[106]),
	.datad(!din_b[108]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_161 ),
	.sharein(Xd_0__inst_mult_15_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_157 ),
	.shareout(Xd_0__inst_mult_15_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_46 (
// Equation(s):
// Xd_0__inst_mult_12_157  = CARRY(( (din_a[86] & din_b[86]) ) + ( Xd_0__inst_mult_12_162  ) + ( Xd_0__inst_mult_12_161  ))
// Xd_0__inst_mult_12_158  = SHARE((din_a[85] & din_b[87]))

	.dataa(!din_a[86]),
	.datab(!din_b[86]),
	.datac(!din_a[85]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_161 ),
	.sharein(Xd_0__inst_mult_12_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_157 ),
	.shareout(Xd_0__inst_mult_12_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_46 (
// Equation(s):
// Xd_0__inst_mult_13_157  = CARRY(( (din_a[93] & din_b[93]) ) + ( Xd_0__inst_mult_13_162  ) + ( Xd_0__inst_mult_13_161  ))
// Xd_0__inst_mult_13_158  = SHARE((din_a[92] & din_b[94]))

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(!din_a[92]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_161 ),
	.sharein(Xd_0__inst_mult_13_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_157 ),
	.shareout(Xd_0__inst_mult_13_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_46 (
// Equation(s):
// Xd_0__inst_mult_10_157  = CARRY(( (din_a[72] & din_b[72]) ) + ( Xd_0__inst_mult_10_162  ) + ( Xd_0__inst_mult_10_161  ))
// Xd_0__inst_mult_10_158  = SHARE((din_a[71] & din_b[73]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_a[71]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_161 ),
	.sharein(Xd_0__inst_mult_10_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_157 ),
	.shareout(Xd_0__inst_mult_10_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_46 (
// Equation(s):
// Xd_0__inst_mult_11_157  = CARRY(( (din_a[79] & din_b[79]) ) + ( Xd_0__inst_mult_11_162  ) + ( Xd_0__inst_mult_11_161  ))
// Xd_0__inst_mult_11_158  = SHARE((din_a[78] & din_b[80]))

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(!din_a[78]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_161 ),
	.sharein(Xd_0__inst_mult_11_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_157 ),
	.shareout(Xd_0__inst_mult_11_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_46 (
// Equation(s):
// Xd_0__inst_mult_8_157  = CARRY(( (din_a[58] & din_b[58]) ) + ( Xd_0__inst_mult_8_162  ) + ( Xd_0__inst_mult_8_161  ))
// Xd_0__inst_mult_8_158  = SHARE((din_a[57] & din_b[59]))

	.dataa(!din_a[58]),
	.datab(!din_b[58]),
	.datac(!din_a[57]),
	.datad(!din_b[59]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_161 ),
	.sharein(Xd_0__inst_mult_8_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_157 ),
	.shareout(Xd_0__inst_mult_8_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_46 (
// Equation(s):
// Xd_0__inst_mult_9_157  = CARRY(( (din_a[65] & din_b[65]) ) + ( Xd_0__inst_mult_9_162  ) + ( Xd_0__inst_mult_9_161  ))
// Xd_0__inst_mult_9_158  = SHARE((din_a[64] & din_b[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(!din_a[64]),
	.datad(!din_b[66]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_161 ),
	.sharein(Xd_0__inst_mult_9_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_157 ),
	.shareout(Xd_0__inst_mult_9_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_46 (
// Equation(s):
// Xd_0__inst_mult_6_157  = CARRY(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_6_162  ) + ( Xd_0__inst_mult_6_161  ))
// Xd_0__inst_mult_6_158  = SHARE((din_a[43] & din_b[45]))

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(!din_a[43]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_161 ),
	.sharein(Xd_0__inst_mult_6_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_157 ),
	.shareout(Xd_0__inst_mult_6_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_46 (
// Equation(s):
// Xd_0__inst_mult_7_157  = CARRY(( (din_a[51] & din_b[51]) ) + ( Xd_0__inst_mult_7_162  ) + ( Xd_0__inst_mult_7_161  ))
// Xd_0__inst_mult_7_158  = SHARE((din_a[50] & din_b[52]))

	.dataa(!din_a[51]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_161 ),
	.sharein(Xd_0__inst_mult_7_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_157 ),
	.shareout(Xd_0__inst_mult_7_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_46 (
// Equation(s):
// Xd_0__inst_mult_4_157  = CARRY(( (din_a[30] & din_b[30]) ) + ( Xd_0__inst_mult_4_162  ) + ( Xd_0__inst_mult_4_161  ))
// Xd_0__inst_mult_4_158  = SHARE((din_a[29] & din_b[31]))

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(!din_a[29]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_161 ),
	.sharein(Xd_0__inst_mult_4_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_157 ),
	.shareout(Xd_0__inst_mult_4_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_46 (
// Equation(s):
// Xd_0__inst_mult_5_157  = CARRY(( (din_a[37] & din_b[37]) ) + ( Xd_0__inst_mult_5_162  ) + ( Xd_0__inst_mult_5_161  ))
// Xd_0__inst_mult_5_158  = SHARE((din_a[36] & din_b[38]))

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[36]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_161 ),
	.sharein(Xd_0__inst_mult_5_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_157 ),
	.shareout(Xd_0__inst_mult_5_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_46 (
// Equation(s):
// Xd_0__inst_mult_2_157  = CARRY(( (din_a[16] & din_b[16]) ) + ( Xd_0__inst_mult_2_162  ) + ( Xd_0__inst_mult_2_161  ))
// Xd_0__inst_mult_2_158  = SHARE((din_a[15] & din_b[17]))

	.dataa(!din_a[16]),
	.datab(!din_b[16]),
	.datac(!din_a[15]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_161 ),
	.sharein(Xd_0__inst_mult_2_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_157 ),
	.shareout(Xd_0__inst_mult_2_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_46 (
// Equation(s):
// Xd_0__inst_mult_3_157  = CARRY(( (din_a[23] & din_b[23]) ) + ( Xd_0__inst_mult_3_162  ) + ( Xd_0__inst_mult_3_161  ))
// Xd_0__inst_mult_3_158  = SHARE((din_a[22] & din_b[24]))

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(!din_a[22]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_161 ),
	.sharein(Xd_0__inst_mult_3_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_157 ),
	.shareout(Xd_0__inst_mult_3_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_46 (
// Equation(s):
// Xd_0__inst_mult_0_157  = CARRY(( (din_a[2] & din_b[2]) ) + ( Xd_0__inst_mult_0_162  ) + ( Xd_0__inst_mult_0_161  ))
// Xd_0__inst_mult_0_158  = SHARE((din_a[1] & din_b[3]))

	.dataa(!din_a[2]),
	.datab(!din_b[2]),
	.datac(!din_a[1]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_161 ),
	.sharein(Xd_0__inst_mult_0_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_157 ),
	.shareout(Xd_0__inst_mult_0_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_46 (
// Equation(s):
// Xd_0__inst_mult_1_157  = CARRY(( (din_a[9] & din_b[9]) ) + ( Xd_0__inst_mult_1_162  ) + ( Xd_0__inst_mult_1_161  ))
// Xd_0__inst_mult_1_158  = SHARE((din_a[8] & din_b[10]))

	.dataa(!din_a[9]),
	.datab(!din_b[9]),
	.datac(!din_a[8]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_161 ),
	.sharein(Xd_0__inst_mult_1_162 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_157 ),
	.shareout(Xd_0__inst_mult_1_158 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_47 (
// Equation(s):
// Xd_0__inst_mult_28_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_28_162  = SHARE((din_a[198] & din_b[198]))

	.dataa(!din_a[198]),
	.datab(!din_b[198]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_161 ),
	.shareout(Xd_0__inst_mult_28_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_47 (
// Equation(s):
// Xd_0__inst_mult_29_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_29_162  = SHARE((din_a[205] & din_b[205]))

	.dataa(!din_a[205]),
	.datab(!din_b[205]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_161 ),
	.shareout(Xd_0__inst_mult_29_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_47 (
// Equation(s):
// Xd_0__inst_mult_26_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_26_162  = SHARE((din_a[184] & din_b[184]))

	.dataa(!din_a[184]),
	.datab(!din_b[184]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_161 ),
	.shareout(Xd_0__inst_mult_26_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_47 (
// Equation(s):
// Xd_0__inst_mult_27_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_27_162  = SHARE((din_a[191] & din_b[191]))

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_161 ),
	.shareout(Xd_0__inst_mult_27_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_47 (
// Equation(s):
// Xd_0__inst_mult_24_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_24_162  = SHARE((din_a[170] & din_b[170]))

	.dataa(!din_a[170]),
	.datab(!din_b[170]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_161 ),
	.shareout(Xd_0__inst_mult_24_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_47 (
// Equation(s):
// Xd_0__inst_mult_25_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_25_162  = SHARE((din_a[177] & din_b[177]))

	.dataa(!din_a[177]),
	.datab(!din_b[177]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_161 ),
	.shareout(Xd_0__inst_mult_25_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_47 (
// Equation(s):
// Xd_0__inst_mult_22_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_22_162  = SHARE((din_a[156] & din_b[156]))

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_161 ),
	.shareout(Xd_0__inst_mult_22_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_47 (
// Equation(s):
// Xd_0__inst_mult_23_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_23_162  = SHARE((din_a[163] & din_b[163]))

	.dataa(!din_a[163]),
	.datab(!din_b[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_161 ),
	.shareout(Xd_0__inst_mult_23_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_47 (
// Equation(s):
// Xd_0__inst_mult_20_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_20_162  = SHARE((din_a[142] & din_b[142]))

	.dataa(!din_a[142]),
	.datab(!din_b[142]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_161 ),
	.shareout(Xd_0__inst_mult_20_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_47 (
// Equation(s):
// Xd_0__inst_mult_21_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_21_162  = SHARE((din_a[149] & din_b[149]))

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_161 ),
	.shareout(Xd_0__inst_mult_21_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_47 (
// Equation(s):
// Xd_0__inst_mult_18_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_18_162  = SHARE((din_a[128] & din_b[128]))

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_161 ),
	.shareout(Xd_0__inst_mult_18_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_47 (
// Equation(s):
// Xd_0__inst_mult_19_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_19_162  = SHARE((din_a[135] & din_b[135]))

	.dataa(!din_a[135]),
	.datab(!din_b[135]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_161 ),
	.shareout(Xd_0__inst_mult_19_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_47 (
// Equation(s):
// Xd_0__inst_mult_16_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_16_162  = SHARE((din_a[114] & din_b[114]))

	.dataa(!din_a[114]),
	.datab(!din_b[114]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_161 ),
	.shareout(Xd_0__inst_mult_16_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_47 (
// Equation(s):
// Xd_0__inst_mult_17_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_17_162  = SHARE((din_a[121] & din_b[121]))

	.dataa(!din_a[121]),
	.datab(!din_b[121]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_161 ),
	.shareout(Xd_0__inst_mult_17_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_47 (
// Equation(s):
// Xd_0__inst_mult_14_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_14_162  = SHARE((din_a[100] & din_b[100]))

	.dataa(!din_a[100]),
	.datab(!din_b[100]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_161 ),
	.shareout(Xd_0__inst_mult_14_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_47 (
// Equation(s):
// Xd_0__inst_mult_15_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_15_162  = SHARE((din_a[107] & din_b[107]))

	.dataa(!din_a[107]),
	.datab(!din_b[107]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_161 ),
	.shareout(Xd_0__inst_mult_15_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_47 (
// Equation(s):
// Xd_0__inst_mult_12_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_162  = SHARE((din_a[86] & din_b[86]))

	.dataa(!din_a[86]),
	.datab(!din_b[86]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_161 ),
	.shareout(Xd_0__inst_mult_12_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_47 (
// Equation(s):
// Xd_0__inst_mult_13_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_13_162  = SHARE((din_a[93] & din_b[93]))

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_161 ),
	.shareout(Xd_0__inst_mult_13_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_47 (
// Equation(s):
// Xd_0__inst_mult_10_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_10_162  = SHARE((din_a[72] & din_b[72]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_161 ),
	.shareout(Xd_0__inst_mult_10_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_47 (
// Equation(s):
// Xd_0__inst_mult_11_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_162  = SHARE((din_a[79] & din_b[79]))

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_161 ),
	.shareout(Xd_0__inst_mult_11_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_47 (
// Equation(s):
// Xd_0__inst_mult_8_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_8_162  = SHARE((din_a[58] & din_b[58]))

	.dataa(!din_a[58]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_161 ),
	.shareout(Xd_0__inst_mult_8_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_47 (
// Equation(s):
// Xd_0__inst_mult_9_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_9_162  = SHARE((din_a[65] & din_b[65]))

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_161 ),
	.shareout(Xd_0__inst_mult_9_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_47 (
// Equation(s):
// Xd_0__inst_mult_6_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_162  = SHARE((din_a[44] & din_b[44]))

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_161 ),
	.shareout(Xd_0__inst_mult_6_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_47 (
// Equation(s):
// Xd_0__inst_mult_7_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_162  = SHARE((din_a[51] & din_b[51]))

	.dataa(!din_a[51]),
	.datab(!din_b[51]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_161 ),
	.shareout(Xd_0__inst_mult_7_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_47 (
// Equation(s):
// Xd_0__inst_mult_4_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_162  = SHARE((din_a[30] & din_b[30]))

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_161 ),
	.shareout(Xd_0__inst_mult_4_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_47 (
// Equation(s):
// Xd_0__inst_mult_5_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_162  = SHARE((din_a[37] & din_b[37]))

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_161 ),
	.shareout(Xd_0__inst_mult_5_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_47 (
// Equation(s):
// Xd_0__inst_mult_2_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_162  = SHARE((din_a[16] & din_b[16]))

	.dataa(!din_a[16]),
	.datab(!din_b[16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_161 ),
	.shareout(Xd_0__inst_mult_2_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_47 (
// Equation(s):
// Xd_0__inst_mult_3_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_162  = SHARE((din_a[23] & din_b[23]))

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_161 ),
	.shareout(Xd_0__inst_mult_3_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_47 (
// Equation(s):
// Xd_0__inst_mult_0_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_162  = SHARE((din_a[2] & din_b[2]))

	.dataa(!din_a[2]),
	.datab(!din_b[2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_161 ),
	.shareout(Xd_0__inst_mult_0_162 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_47 (
// Equation(s):
// Xd_0__inst_mult_1_161  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_162  = SHARE((din_a[9] & din_b[9]))

	.dataa(!din_a[9]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_161 ),
	.shareout(Xd_0__inst_mult_1_162 ));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__5__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__6__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__7__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__8__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__9__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__10__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__11__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__12__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__13__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_30_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [30]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_31_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [31]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_28_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [28]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_29_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [29]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_26_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [26]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_27_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [27]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_24_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_25_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_22_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_23_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_20_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_21_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_18_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_19_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_30_ (
	.clk(clk),
	.d(Xd_0__inst_i19_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [30]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_31_ (
	.clk(clk),
	.d(Xd_0__inst_i19_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [31]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_16_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_17_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_56 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_60 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_64 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_68 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_72 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_76 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_80 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_28_ (
	.clk(clk),
	.d(Xd_0__inst_i19_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [28]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_29_ (
	.clk(clk),
	.d(Xd_0__inst_i19_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [29]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_26_ (
	.clk(clk),
	.d(Xd_0__inst_i19_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [26]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_27_ (
	.clk(clk),
	.d(Xd_0__inst_i19_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [27]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_24_ (
	.clk(clk),
	.d(Xd_0__inst_i19_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_25_ (
	.clk(clk),
	.d(Xd_0__inst_i19_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_22_ (
	.clk(clk),
	.d(Xd_0__inst_i19_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_23_ (
	.clk(clk),
	.d(Xd_0__inst_i19_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_20_ (
	.clk(clk),
	.d(Xd_0__inst_i19_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_21_ (
	.clk(clk),
	.d(Xd_0__inst_i19_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_18_ (
	.clk(clk),
	.d(Xd_0__inst_i19_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_19_ (
	.clk(clk),
	.d(Xd_0__inst_i19_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_16_ (
	.clk(clk),
	.d(Xd_0__inst_i19_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_17_ (
	.clk(clk),
	.d(Xd_0__inst_i19_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_14_ (
	.clk(clk),
	.d(Xd_0__inst_i19_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_15_ (
	.clk(clk),
	.d(Xd_0__inst_i19_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_12_ (
	.clk(clk),
	.d(Xd_0__inst_i19_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_13_ (
	.clk(clk),
	.d(Xd_0__inst_i19_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_10_ (
	.clk(clk),
	.d(Xd_0__inst_i19_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_11_ (
	.clk(clk),
	.d(Xd_0__inst_i19_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_8_ (
	.clk(clk),
	.d(Xd_0__inst_i19_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_9_ (
	.clk(clk),
	.d(Xd_0__inst_i19_109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i19_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i19_105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i19_113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i19_117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i19_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i19_125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_84 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i19_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i19_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_96 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_96 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_92 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_2 (
	.clk(clk),
	.d(din_a[213]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_3 (
	.clk(clk),
	.d(din_b[210]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_2 (
	.clk(clk),
	.d(din_a[220]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_3 (
	.clk(clk),
	.d(din_b[217]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_7 (
	.clk(clk),
	.d(din_a[214]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_7 (
	.clk(clk),
	.d(din_a[221]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_1 (
	.clk(clk),
	.d(din_b[213]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_1 (
	.clk(clk),
	.d(din_b[220]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_18 (
	.clk(clk),
	.d(din_b[215]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_18 (
	.clk(clk),
	.d(din_b[222]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_19 (
	.clk(clk),
	.d(din_a[215]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_19 (
	.clk(clk),
	.d(din_a[222]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_2 (
	.clk(clk),
	.d(din_a[199]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_3 (
	.clk(clk),
	.d(din_b[196]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_2 (
	.clk(clk),
	.d(din_a[206]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_3 (
	.clk(clk),
	.d(din_b[203]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_2 (
	.clk(clk),
	.d(din_a[185]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_3 (
	.clk(clk),
	.d(din_b[182]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_2 (
	.clk(clk),
	.d(din_a[192]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_3 (
	.clk(clk),
	.d(din_b[189]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_2 (
	.clk(clk),
	.d(din_a[171]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_3 (
	.clk(clk),
	.d(din_b[168]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_2 (
	.clk(clk),
	.d(din_a[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_3 (
	.clk(clk),
	.d(din_b[175]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_2 (
	.clk(clk),
	.d(din_a[157]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_3 (
	.clk(clk),
	.d(din_b[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_2 (
	.clk(clk),
	.d(din_a[164]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_3 (
	.clk(clk),
	.d(din_b[161]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_2 (
	.clk(clk),
	.d(din_a[143]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_3 (
	.clk(clk),
	.d(din_b[140]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_2 (
	.clk(clk),
	.d(din_a[150]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_3 (
	.clk(clk),
	.d(din_b[147]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_2 (
	.clk(clk),
	.d(din_a[129]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_3 (
	.clk(clk),
	.d(din_b[126]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_2 (
	.clk(clk),
	.d(din_a[136]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_3 (
	.clk(clk),
	.d(din_b[133]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_0 (
	.clk(clk),
	.d(din_a[210]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_0 (
	.clk(clk),
	.d(din_a[217]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_2 (
	.clk(clk),
	.d(din_a[115]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_3 (
	.clk(clk),
	.d(din_b[112]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_2 (
	.clk(clk),
	.d(din_a[122]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_3 (
	.clk(clk),
	.d(din_b[119]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_2 (
	.clk(clk),
	.d(din_a[101]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_3 (
	.clk(clk),
	.d(din_b[98]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_2 (
	.clk(clk),
	.d(din_a[108]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_3 (
	.clk(clk),
	.d(din_b[105]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_2 (
	.clk(clk),
	.d(din_a[87]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_3 (
	.clk(clk),
	.d(din_b[84]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_2 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_3 (
	.clk(clk),
	.d(din_b[91]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_2 (
	.clk(clk),
	.d(din_a[73]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_3 (
	.clk(clk),
	.d(din_b[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_2 (
	.clk(clk),
	.d(din_a[80]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_3 (
	.clk(clk),
	.d(din_b[77]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_2 (
	.clk(clk),
	.d(din_a[59]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_3 (
	.clk(clk),
	.d(din_b[56]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_2 (
	.clk(clk),
	.d(din_a[66]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_3 (
	.clk(clk),
	.d(din_b[63]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(din_a[45]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(din_b[42]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(din_a[52]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(din_b[49]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(din_a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(din_b[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(din_a[38]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(din_b[35]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(din_a[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(din_b[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(din_a[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(din_b[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(din_a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(din_b[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(din_a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(din_b[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_7 (
	.clk(clk),
	.d(din_a[200]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_7 (
	.clk(clk),
	.d(din_a[207]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_7 (
	.clk(clk),
	.d(din_a[186]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_7 (
	.clk(clk),
	.d(din_a[193]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_7 (
	.clk(clk),
	.d(din_a[172]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_7 (
	.clk(clk),
	.d(din_a[179]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_7 (
	.clk(clk),
	.d(din_a[158]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_7 (
	.clk(clk),
	.d(din_a[165]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_7 (
	.clk(clk),
	.d(din_a[144]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_7 (
	.clk(clk),
	.d(din_a[151]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_7 (
	.clk(clk),
	.d(din_a[130]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_7 (
	.clk(clk),
	.d(din_a[137]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_7 (
	.clk(clk),
	.d(din_a[116]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_7 (
	.clk(clk),
	.d(din_a[123]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_7 (
	.clk(clk),
	.d(din_a[102]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_7 (
	.clk(clk),
	.d(din_a[109]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_7 (
	.clk(clk),
	.d(din_a[88]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_7 (
	.clk(clk),
	.d(din_a[95]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_7 (
	.clk(clk),
	.d(din_a[74]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_7 (
	.clk(clk),
	.d(din_a[81]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_7 (
	.clk(clk),
	.d(din_a[60]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_7 (
	.clk(clk),
	.d(din_a[67]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(din_a[53]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(din_a[32]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(din_a[39]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(din_a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(din_a[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(din_a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_108 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_112 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(din_a[11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_116 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_120 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_1 (
	.clk(clk),
	.d(din_b[199]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_1 (
	.clk(clk),
	.d(din_b[206]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_1 (
	.clk(clk),
	.d(din_b[185]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_1 (
	.clk(clk),
	.d(din_b[192]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_1 (
	.clk(clk),
	.d(din_b[171]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_1 (
	.clk(clk),
	.d(din_b[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_1 (
	.clk(clk),
	.d(din_b[157]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_1 (
	.clk(clk),
	.d(din_b[164]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_1 (
	.clk(clk),
	.d(din_b[143]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_1 (
	.clk(clk),
	.d(din_b[150]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_1 (
	.clk(clk),
	.d(din_b[129]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_1 (
	.clk(clk),
	.d(din_b[136]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_1 (
	.clk(clk),
	.d(din_b[115]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_1 (
	.clk(clk),
	.d(din_b[122]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_1 (
	.clk(clk),
	.d(din_b[101]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_1 (
	.clk(clk),
	.d(din_b[108]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_1 (
	.clk(clk),
	.d(din_b[87]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_1 (
	.clk(clk),
	.d(din_b[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_1 (
	.clk(clk),
	.d(din_b[73]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_1 (
	.clk(clk),
	.d(din_b[80]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_1 (
	.clk(clk),
	.d(din_b[59]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_1 (
	.clk(clk),
	.d(din_b[66]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(din_b[45]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(din_b[52]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(din_b[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(din_b[38]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(din_b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(din_b[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(din_b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_124 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_128 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(din_b[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_132 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_136 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_104 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_140 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_144 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_18 (
	.clk(clk),
	.d(din_b[201]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_18 (
	.clk(clk),
	.d(din_b[208]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_18 (
	.clk(clk),
	.d(din_b[187]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_18 (
	.clk(clk),
	.d(din_b[194]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_18 (
	.clk(clk),
	.d(din_b[173]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_18 (
	.clk(clk),
	.d(din_b[180]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_88 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_18 (
	.clk(clk),
	.d(din_b[159]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_18 (
	.clk(clk),
	.d(din_b[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_18 (
	.clk(clk),
	.d(din_b[145]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_18 (
	.clk(clk),
	.d(din_b[152]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_18 (
	.clk(clk),
	.d(din_b[131]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_18 (
	.clk(clk),
	.d(din_b[138]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_18 (
	.clk(clk),
	.d(din_b[117]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_18 (
	.clk(clk),
	.d(din_b[124]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_18 (
	.clk(clk),
	.d(din_b[103]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_18 (
	.clk(clk),
	.d(din_b[110]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_18 (
	.clk(clk),
	.d(din_b[89]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_18 (
	.clk(clk),
	.d(din_b[96]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_18 (
	.clk(clk),
	.d(din_b[75]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_18 (
	.clk(clk),
	.d(din_b[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_18 (
	.clk(clk),
	.d(din_b[61]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_18 (
	.clk(clk),
	.d(din_b[68]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_18 (
	.clk(clk),
	.d(din_b[47]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_18 (
	.clk(clk),
	.d(din_b[54]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_18 (
	.clk(clk),
	.d(din_b[33]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_18 (
	.clk(clk),
	.d(din_b[40]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_18 (
	.clk(clk),
	.d(din_b[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_18 (
	.clk(clk),
	.d(din_b[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_18 (
	.clk(clk),
	.d(din_b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_148 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_100 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_18 (
	.clk(clk),
	.d(din_b[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_19 (
	.clk(clk),
	.d(din_a[201]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_19 (
	.clk(clk),
	.d(din_a[208]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_19 (
	.clk(clk),
	.d(din_a[187]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_19 (
	.clk(clk),
	.d(din_a[194]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_19 (
	.clk(clk),
	.d(din_a[173]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_19 (
	.clk(clk),
	.d(din_a[180]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_19 (
	.clk(clk),
	.d(din_a[159]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_19 (
	.clk(clk),
	.d(din_a[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_19 (
	.clk(clk),
	.d(din_a[145]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_19 (
	.clk(clk),
	.d(din_a[152]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_19 (
	.clk(clk),
	.d(din_a[131]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_19 (
	.clk(clk),
	.d(din_a[138]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_19 (
	.clk(clk),
	.d(din_a[117]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_19 (
	.clk(clk),
	.d(din_a[124]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_19 (
	.clk(clk),
	.d(din_a[103]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_19 (
	.clk(clk),
	.d(din_a[110]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_19 (
	.clk(clk),
	.d(din_a[89]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_19 (
	.clk(clk),
	.d(din_a[96]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_19 (
	.clk(clk),
	.d(din_a[75]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_19 (
	.clk(clk),
	.d(din_a[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_19 (
	.clk(clk),
	.d(din_a[61]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_19 (
	.clk(clk),
	.d(din_a[68]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_19 (
	.clk(clk),
	.d(din_a[47]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_19 (
	.clk(clk),
	.d(din_a[54]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_19 (
	.clk(clk),
	.d(din_a[33]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_19 (
	.clk(clk),
	.d(din_a[40]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_19 (
	.clk(clk),
	.d(din_a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_19 (
	.clk(clk),
	.d(din_a[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_19 (
	.clk(clk),
	.d(din_a[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_19 (
	.clk(clk),
	.d(din_a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_152 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_0 (
	.clk(clk),
	.d(din_a[196]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_0 (
	.clk(clk),
	.d(din_a[203]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_0 (
	.clk(clk),
	.d(din_a[182]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_0 (
	.clk(clk),
	.d(din_a[189]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_0 (
	.clk(clk),
	.d(din_a[168]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_0 (
	.clk(clk),
	.d(din_a[175]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_0 (
	.clk(clk),
	.d(din_a[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_0 (
	.clk(clk),
	.d(din_a[161]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_0 (
	.clk(clk),
	.d(din_a[140]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_0 (
	.clk(clk),
	.d(din_a[147]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_0 (
	.clk(clk),
	.d(din_a[126]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_0 (
	.clk(clk),
	.d(din_a[133]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_0 (
	.clk(clk),
	.d(din_a[112]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_0 (
	.clk(clk),
	.d(din_a[119]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_0 (
	.clk(clk),
	.d(din_a[98]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_0 (
	.clk(clk),
	.d(din_a[105]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_0 (
	.clk(clk),
	.d(din_a[84]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_0 (
	.clk(clk),
	.d(din_a[91]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_0 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_0 (
	.clk(clk),
	.d(din_a[77]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_0 (
	.clk(clk),
	.d(din_a[56]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_0 (
	.clk(clk),
	.d(din_a[63]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(din_a[42]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(din_a[49]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(din_a[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(din_a[35]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(din_a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(din_a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(din_a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(din_a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ),
	.prn(vcc));

assign dout[0] = Xd_0__inst_inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_inst_dout [15];

assign dout[16] = Xd_0__inst_inst_inst_inst_dout [16];

assign dout[17] = Xd_0__inst_inst_inst_inst_dout [17];

endmodule
