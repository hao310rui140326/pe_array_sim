// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:31:28"

// 
// Device: Altera 10AX115S2F45I1SG Package FBGA1932
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_a10_6x6x32 (
	dout,
	clk,
	din_a,
	din_b);
output 	[15:0] dout;
input 	clk;
input 	[191:0] din_a;
input 	[191:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_inst_add_0_3 ;
wire Xd_0__inst_inst_inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_6 ;
wire Xd_0__inst_inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_10 ;
wire Xd_0__inst_inst_inst_inst_add_0_11 ;
wire Xd_0__inst_inst_inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_14 ;
wire Xd_0__inst_inst_inst_inst_add_0_15 ;
wire Xd_0__inst_inst_inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_18 ;
wire Xd_0__inst_inst_inst_inst_add_0_19 ;
wire Xd_0__inst_inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_inst_add_0_23 ;
wire Xd_0__inst_inst_inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_26 ;
wire Xd_0__inst_inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_30 ;
wire Xd_0__inst_inst_inst_inst_add_0_31 ;
wire Xd_0__inst_inst_inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_34 ;
wire Xd_0__inst_inst_inst_inst_add_0_35 ;
wire Xd_0__inst_inst_inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_38 ;
wire Xd_0__inst_inst_inst_inst_add_0_39 ;
wire Xd_0__inst_inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_inst_add_0_43 ;
wire Xd_0__inst_inst_inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_46 ;
wire Xd_0__inst_inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_50 ;
wire Xd_0__inst_inst_inst_inst_add_0_51 ;
wire Xd_0__inst_inst_inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_54 ;
wire Xd_0__inst_inst_inst_inst_add_0_55 ;
wire Xd_0__inst_inst_inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_inst_inst_add_0_58 ;
wire Xd_0__inst_inst_inst_inst_add_0_59 ;
wire Xd_0__inst_inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_mult_24_36 ;
wire Xd_0__inst_mult_24_37 ;
wire Xd_0__inst_mult_24_38 ;
wire Xd_0__inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_add_0_3 ;
wire Xd_0__inst_inst_inst_add_3_1_sumout ;
wire Xd_0__inst_inst_inst_add_3_2 ;
wire Xd_0__inst_inst_inst_add_3_3 ;
wire Xd_0__inst_mult_24_40 ;
wire Xd_0__inst_mult_24_41 ;
wire Xd_0__inst_mult_24_42 ;
wire Xd_0__inst_inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_inst_add_0_6 ;
wire Xd_0__inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_add_3_5_sumout ;
wire Xd_0__inst_inst_inst_add_3_6 ;
wire Xd_0__inst_inst_inst_add_3_7 ;
wire Xd_0__inst_inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_inst_add_0_10 ;
wire Xd_0__inst_inst_inst_add_0_11 ;
wire Xd_0__inst_inst_inst_add_3_9_sumout ;
wire Xd_0__inst_inst_inst_add_3_10 ;
wire Xd_0__inst_inst_inst_add_3_11 ;
wire Xd_0__inst_inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_inst_add_0_14 ;
wire Xd_0__inst_inst_inst_add_0_15 ;
wire Xd_0__inst_inst_inst_add_3_13_sumout ;
wire Xd_0__inst_inst_inst_add_3_14 ;
wire Xd_0__inst_inst_inst_add_3_15 ;
wire Xd_0__inst_inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_inst_add_0_18 ;
wire Xd_0__inst_inst_inst_add_0_19 ;
wire Xd_0__inst_inst_inst_add_3_17_sumout ;
wire Xd_0__inst_inst_inst_add_3_18 ;
wire Xd_0__inst_inst_inst_add_3_19 ;
wire Xd_0__inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_add_0_23 ;
wire Xd_0__inst_inst_inst_add_3_21_sumout ;
wire Xd_0__inst_inst_inst_add_3_22 ;
wire Xd_0__inst_inst_inst_add_3_23 ;
wire Xd_0__inst_inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_inst_add_0_26 ;
wire Xd_0__inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_add_3_25_sumout ;
wire Xd_0__inst_inst_inst_add_3_26 ;
wire Xd_0__inst_inst_inst_add_3_27 ;
wire Xd_0__inst_inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_inst_add_0_30 ;
wire Xd_0__inst_inst_inst_add_0_31 ;
wire Xd_0__inst_inst_inst_add_3_29_sumout ;
wire Xd_0__inst_inst_inst_add_3_30 ;
wire Xd_0__inst_inst_inst_add_3_31 ;
wire Xd_0__inst_inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_inst_add_0_34 ;
wire Xd_0__inst_inst_inst_add_0_35 ;
wire Xd_0__inst_inst_inst_add_3_33_sumout ;
wire Xd_0__inst_inst_inst_add_3_34 ;
wire Xd_0__inst_inst_inst_add_3_35 ;
wire Xd_0__inst_inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_inst_add_0_38 ;
wire Xd_0__inst_inst_inst_add_0_39 ;
wire Xd_0__inst_inst_inst_add_3_37_sumout ;
wire Xd_0__inst_inst_inst_add_3_38 ;
wire Xd_0__inst_inst_inst_add_3_39 ;
wire Xd_0__inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_add_0_43 ;
wire Xd_0__inst_inst_inst_add_3_41_sumout ;
wire Xd_0__inst_inst_inst_add_3_42 ;
wire Xd_0__inst_inst_inst_add_3_43 ;
wire Xd_0__inst_inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_inst_add_0_46 ;
wire Xd_0__inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_add_3_45_sumout ;
wire Xd_0__inst_inst_inst_add_3_46 ;
wire Xd_0__inst_inst_inst_add_3_47 ;
wire Xd_0__inst_inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_inst_add_0_50 ;
wire Xd_0__inst_inst_inst_add_0_51 ;
wire Xd_0__inst_inst_inst_add_3_49_sumout ;
wire Xd_0__inst_inst_inst_add_3_50 ;
wire Xd_0__inst_inst_inst_add_3_51 ;
wire Xd_0__inst_inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_inst_add_0_54 ;
wire Xd_0__inst_inst_inst_add_0_55 ;
wire Xd_0__inst_inst_inst_add_3_53_sumout ;
wire Xd_0__inst_inst_inst_add_3_54 ;
wire Xd_0__inst_inst_inst_add_3_55 ;
wire Xd_0__inst_inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_inst_add_0_58 ;
wire Xd_0__inst_inst_inst_add_0_59 ;
wire Xd_0__inst_inst_inst_add_3_57_sumout ;
wire Xd_0__inst_inst_inst_add_3_58 ;
wire Xd_0__inst_inst_inst_add_3_59 ;
wire Xd_0__inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_add_3_61_sumout ;
wire Xd_0__inst_mult_20_36 ;
wire Xd_0__inst_mult_20_37 ;
wire Xd_0__inst_mult_20_38 ;
wire Xd_0__inst_mult_23_36 ;
wire Xd_0__inst_mult_23_37 ;
wire Xd_0__inst_mult_23_38 ;
wire Xd_0__inst_mult_24_44 ;
wire Xd_0__inst_mult_24_45 ;
wire Xd_0__inst_inst_add_4_1_sumout ;
wire Xd_0__inst_inst_add_4_2 ;
wire Xd_0__inst_inst_add_4_3 ;
wire Xd_0__inst_inst_add_2_1_sumout ;
wire Xd_0__inst_inst_add_2_2 ;
wire Xd_0__inst_inst_add_2_3 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_inst_add_0_3 ;
wire Xd_0__inst_mult_20_40 ;
wire Xd_0__inst_mult_20_41 ;
wire Xd_0__inst_mult_20_42 ;
wire Xd_0__inst_inst_add_8_1_sumout ;
wire Xd_0__inst_inst_add_8_2 ;
wire Xd_0__inst_inst_add_8_3 ;
wire Xd_0__inst_inst_add_6_1_sumout ;
wire Xd_0__inst_inst_add_6_2 ;
wire Xd_0__inst_inst_add_6_3 ;
wire Xd_0__inst_mult_23_40 ;
wire Xd_0__inst_mult_23_41 ;
wire Xd_0__inst_mult_23_42 ;
wire Xd_0__inst_i17_1_sumout ;
wire Xd_0__inst_i17_2 ;
wire Xd_0__inst_i17_3 ;
wire Xd_0__inst_inst_add_4_5_sumout ;
wire Xd_0__inst_inst_add_4_6 ;
wire Xd_0__inst_inst_add_4_7 ;
wire Xd_0__inst_inst_add_2_5_sumout ;
wire Xd_0__inst_inst_add_2_6 ;
wire Xd_0__inst_inst_add_2_7 ;
wire Xd_0__inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_add_0_6 ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_8_5_sumout ;
wire Xd_0__inst_inst_add_8_6 ;
wire Xd_0__inst_inst_add_8_7 ;
wire Xd_0__inst_inst_add_6_5_sumout ;
wire Xd_0__inst_inst_add_6_6 ;
wire Xd_0__inst_inst_add_6_7 ;
wire Xd_0__inst_inst_add_4_9_sumout ;
wire Xd_0__inst_inst_add_4_10 ;
wire Xd_0__inst_inst_add_4_11 ;
wire Xd_0__inst_inst_add_2_9_sumout ;
wire Xd_0__inst_inst_add_2_10 ;
wire Xd_0__inst_inst_add_2_11 ;
wire Xd_0__inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_add_0_10 ;
wire Xd_0__inst_inst_add_0_11 ;
wire Xd_0__inst_inst_add_8_9_sumout ;
wire Xd_0__inst_inst_add_8_10 ;
wire Xd_0__inst_inst_add_8_11 ;
wire Xd_0__inst_inst_add_6_9_sumout ;
wire Xd_0__inst_inst_add_6_10 ;
wire Xd_0__inst_inst_add_6_11 ;
wire Xd_0__inst_inst_add_4_13_sumout ;
wire Xd_0__inst_inst_add_4_14 ;
wire Xd_0__inst_inst_add_4_15 ;
wire Xd_0__inst_inst_add_2_13_sumout ;
wire Xd_0__inst_inst_add_2_14 ;
wire Xd_0__inst_inst_add_2_15 ;
wire Xd_0__inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_add_0_14 ;
wire Xd_0__inst_inst_add_0_15 ;
wire Xd_0__inst_inst_add_8_13_sumout ;
wire Xd_0__inst_inst_add_8_14 ;
wire Xd_0__inst_inst_add_8_15 ;
wire Xd_0__inst_inst_add_6_13_sumout ;
wire Xd_0__inst_inst_add_6_14 ;
wire Xd_0__inst_inst_add_6_15 ;
wire Xd_0__inst_inst_add_4_17_sumout ;
wire Xd_0__inst_inst_add_4_18 ;
wire Xd_0__inst_inst_add_4_19 ;
wire Xd_0__inst_inst_add_2_17_sumout ;
wire Xd_0__inst_inst_add_2_18 ;
wire Xd_0__inst_inst_add_2_19 ;
wire Xd_0__inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_add_0_18 ;
wire Xd_0__inst_inst_add_0_19 ;
wire Xd_0__inst_inst_add_8_17_sumout ;
wire Xd_0__inst_inst_add_8_18 ;
wire Xd_0__inst_inst_add_8_19 ;
wire Xd_0__inst_inst_add_6_17_sumout ;
wire Xd_0__inst_inst_add_6_18 ;
wire Xd_0__inst_inst_add_6_19 ;
wire Xd_0__inst_inst_add_4_21_sumout ;
wire Xd_0__inst_inst_add_4_22 ;
wire Xd_0__inst_inst_add_4_23 ;
wire Xd_0__inst_inst_add_2_21_sumout ;
wire Xd_0__inst_inst_add_2_22 ;
wire Xd_0__inst_inst_add_2_23 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_0_23 ;
wire Xd_0__inst_inst_add_8_21_sumout ;
wire Xd_0__inst_inst_add_8_22 ;
wire Xd_0__inst_inst_add_8_23 ;
wire Xd_0__inst_inst_add_6_21_sumout ;
wire Xd_0__inst_inst_add_6_22 ;
wire Xd_0__inst_inst_add_6_23 ;
wire Xd_0__inst_inst_add_4_25_sumout ;
wire Xd_0__inst_inst_add_4_26 ;
wire Xd_0__inst_inst_add_4_27 ;
wire Xd_0__inst_inst_add_2_25_sumout ;
wire Xd_0__inst_inst_add_2_26 ;
wire Xd_0__inst_inst_add_2_27 ;
wire Xd_0__inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_add_0_26 ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_8_25_sumout ;
wire Xd_0__inst_inst_add_8_26 ;
wire Xd_0__inst_inst_add_8_27 ;
wire Xd_0__inst_inst_add_6_25_sumout ;
wire Xd_0__inst_inst_add_6_26 ;
wire Xd_0__inst_inst_add_6_27 ;
wire Xd_0__inst_inst_add_4_29_sumout ;
wire Xd_0__inst_inst_add_4_30 ;
wire Xd_0__inst_inst_add_4_31 ;
wire Xd_0__inst_inst_add_2_29_sumout ;
wire Xd_0__inst_inst_add_2_30 ;
wire Xd_0__inst_inst_add_2_31 ;
wire Xd_0__inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_add_0_30 ;
wire Xd_0__inst_inst_add_0_31 ;
wire Xd_0__inst_inst_add_8_29_sumout ;
wire Xd_0__inst_inst_add_8_30 ;
wire Xd_0__inst_inst_add_8_31 ;
wire Xd_0__inst_inst_add_6_29_sumout ;
wire Xd_0__inst_inst_add_6_30 ;
wire Xd_0__inst_inst_add_6_31 ;
wire Xd_0__inst_inst_add_4_33_sumout ;
wire Xd_0__inst_inst_add_4_34 ;
wire Xd_0__inst_inst_add_4_35 ;
wire Xd_0__inst_inst_add_2_33_sumout ;
wire Xd_0__inst_inst_add_2_34 ;
wire Xd_0__inst_inst_add_2_35 ;
wire Xd_0__inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_add_0_34 ;
wire Xd_0__inst_inst_add_0_35 ;
wire Xd_0__inst_inst_add_8_33_sumout ;
wire Xd_0__inst_inst_add_8_34 ;
wire Xd_0__inst_inst_add_8_35 ;
wire Xd_0__inst_inst_add_6_33_sumout ;
wire Xd_0__inst_inst_add_6_34 ;
wire Xd_0__inst_inst_add_6_35 ;
wire Xd_0__inst_inst_add_4_37_sumout ;
wire Xd_0__inst_inst_add_4_38 ;
wire Xd_0__inst_inst_add_4_39 ;
wire Xd_0__inst_inst_add_2_37_sumout ;
wire Xd_0__inst_inst_add_2_38 ;
wire Xd_0__inst_inst_add_2_39 ;
wire Xd_0__inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_add_0_38 ;
wire Xd_0__inst_inst_add_0_39 ;
wire Xd_0__inst_inst_add_8_37_sumout ;
wire Xd_0__inst_inst_add_8_38 ;
wire Xd_0__inst_inst_add_8_39 ;
wire Xd_0__inst_inst_add_6_37_sumout ;
wire Xd_0__inst_inst_add_6_38 ;
wire Xd_0__inst_inst_add_6_39 ;
wire Xd_0__inst_inst_add_4_41_sumout ;
wire Xd_0__inst_inst_add_4_42 ;
wire Xd_0__inst_inst_add_4_43 ;
wire Xd_0__inst_inst_add_2_41_sumout ;
wire Xd_0__inst_inst_add_2_42 ;
wire Xd_0__inst_inst_add_2_43 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_0_43 ;
wire Xd_0__inst_inst_add_8_41_sumout ;
wire Xd_0__inst_inst_add_8_42 ;
wire Xd_0__inst_inst_add_8_43 ;
wire Xd_0__inst_inst_add_6_41_sumout ;
wire Xd_0__inst_inst_add_6_42 ;
wire Xd_0__inst_inst_add_6_43 ;
wire Xd_0__inst_inst_add_4_45_sumout ;
wire Xd_0__inst_inst_add_4_46 ;
wire Xd_0__inst_inst_add_4_47 ;
wire Xd_0__inst_inst_add_2_45_sumout ;
wire Xd_0__inst_inst_add_2_46 ;
wire Xd_0__inst_inst_add_2_47 ;
wire Xd_0__inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_add_0_46 ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_8_45_sumout ;
wire Xd_0__inst_inst_add_8_46 ;
wire Xd_0__inst_inst_add_8_47 ;
wire Xd_0__inst_inst_add_6_45_sumout ;
wire Xd_0__inst_inst_add_6_46 ;
wire Xd_0__inst_inst_add_6_47 ;
wire Xd_0__inst_inst_add_4_49_sumout ;
wire Xd_0__inst_inst_add_4_50 ;
wire Xd_0__inst_inst_add_4_51 ;
wire Xd_0__inst_inst_add_2_49_sumout ;
wire Xd_0__inst_inst_add_2_50 ;
wire Xd_0__inst_inst_add_2_51 ;
wire Xd_0__inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_add_0_50 ;
wire Xd_0__inst_inst_add_0_51 ;
wire Xd_0__inst_inst_add_8_49_sumout ;
wire Xd_0__inst_inst_add_8_50 ;
wire Xd_0__inst_inst_add_8_51 ;
wire Xd_0__inst_inst_add_6_49_sumout ;
wire Xd_0__inst_inst_add_6_50 ;
wire Xd_0__inst_inst_add_6_51 ;
wire Xd_0__inst_inst_add_4_53_sumout ;
wire Xd_0__inst_inst_add_2_53_sumout ;
wire Xd_0__inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_add_8_53_sumout ;
wire Xd_0__inst_inst_add_6_53_sumout ;
wire Xd_0__inst_mult_26_36 ;
wire Xd_0__inst_mult_26_37 ;
wire Xd_0__inst_mult_26_38 ;
wire Xd_0__inst_mult_28_36 ;
wire Xd_0__inst_mult_28_37 ;
wire Xd_0__inst_mult_28_38 ;
wire Xd_0__inst_mult_30_36 ;
wire Xd_0__inst_mult_30_37 ;
wire Xd_0__inst_mult_30_38 ;
wire Xd_0__inst_mult_20_44 ;
wire Xd_0__inst_mult_20_45 ;
wire Xd_0__inst_mult_22_36 ;
wire Xd_0__inst_mult_22_37 ;
wire Xd_0__inst_mult_22_38 ;
wire Xd_0__inst_mult_19_36 ;
wire Xd_0__inst_mult_19_37 ;
wire Xd_0__inst_mult_19_38 ;
wire Xd_0__inst_a1_15__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_23_44 ;
wire Xd_0__inst_mult_23_45 ;
wire Xd_0__inst_a1_15__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_mult_2_35 ;
wire Xd_0__inst_mult_2_36 ;
wire Xd_0__inst_mult_2_37 ;
wire Xd_0__inst_a1_8__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_26_40 ;
wire Xd_0__inst_mult_26_41 ;
wire Xd_0__inst_mult_26_42 ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_28_40 ;
wire Xd_0__inst_mult_28_41 ;
wire Xd_0__inst_mult_28_42 ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_30_40 ;
wire Xd_0__inst_mult_30_41 ;
wire Xd_0__inst_mult_30_42 ;
wire Xd_0__inst_i17_5_sumout ;
wire Xd_0__inst_i17_6 ;
wire Xd_0__inst_i17_7 ;
wire Xd_0__inst_a1_14__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_22_40 ;
wire Xd_0__inst_mult_22_41 ;
wire Xd_0__inst_mult_22_42 ;
wire Xd_0__inst_a1_11__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_19_40 ;
wire Xd_0__inst_mult_19_41 ;
wire Xd_0__inst_mult_19_42 ;
wire Xd_0__inst_i17_9_sumout ;
wire Xd_0__inst_i17_10 ;
wire Xd_0__inst_i17_11 ;
wire Xd_0__inst_a1_8__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_mult_0_35 ;
wire Xd_0__inst_mult_0_36 ;
wire Xd_0__inst_mult_0_37 ;
wire Xd_0__inst_mult_25_36 ;
wire Xd_0__inst_mult_25_37 ;
wire Xd_0__inst_mult_25_38 ;
wire Xd_0__inst_mult_24_47 ;
wire Xd_0__inst_mult_24_48 ;
wire Xd_0__inst_mult_24_49 ;
wire Xd_0__inst_mult_27_36 ;
wire Xd_0__inst_mult_27_37 ;
wire Xd_0__inst_mult_27_38 ;
wire Xd_0__inst_mult_26_43 ;
wire Xd_0__inst_mult_26_44 ;
wire Xd_0__inst_mult_26_45 ;
wire Xd_0__inst_mult_29_36 ;
wire Xd_0__inst_mult_29_37 ;
wire Xd_0__inst_mult_29_38 ;
wire Xd_0__inst_mult_28_43 ;
wire Xd_0__inst_mult_28_44 ;
wire Xd_0__inst_mult_28_45 ;
wire Xd_0__inst_mult_31_36 ;
wire Xd_0__inst_mult_31_37 ;
wire Xd_0__inst_mult_31_38 ;
wire Xd_0__inst_mult_20_47 ;
wire Xd_0__inst_mult_20_48 ;
wire Xd_0__inst_mult_20_49 ;
wire Xd_0__inst_mult_3_35 ;
wire Xd_0__inst_mult_3_36 ;
wire Xd_0__inst_mult_3_37 ;
wire Xd_0__inst_mult_1_35 ;
wire Xd_0__inst_mult_1_36 ;
wire Xd_0__inst_mult_1_37 ;
wire Xd_0__inst_mult_11_36 ;
wire Xd_0__inst_mult_11_37 ;
wire Xd_0__inst_mult_11_38 ;
wire Xd_0__inst_mult_30_43 ;
wire Xd_0__inst_mult_30_44 ;
wire Xd_0__inst_mult_30_45 ;
wire Xd_0__inst_mult_23_47 ;
wire Xd_0__inst_mult_23_48 ;
wire Xd_0__inst_mult_23_49 ;
wire Xd_0__inst_mult_22_43 ;
wire Xd_0__inst_mult_22_44 ;
wire Xd_0__inst_mult_22_45 ;
wire Xd_0__inst_mult_26_48 ;
wire Xd_0__inst_mult_26_49 ;
wire Xd_0__inst_mult_28_48 ;
wire Xd_0__inst_mult_28_49 ;
wire Xd_0__inst_mult_30_48 ;
wire Xd_0__inst_mult_30_49 ;
wire Xd_0__inst_mult_22_48 ;
wire Xd_0__inst_mult_22_49 ;
wire Xd_0__inst_mult_19_44 ;
wire Xd_0__inst_mult_19_45 ;
wire Xd_0__inst_mult_30_51 ;
wire Xd_0__inst_mult_30_52 ;
wire Xd_0__inst_mult_30_53 ;
wire Xd_0__inst_mult_31_40 ;
wire Xd_0__inst_mult_31_41 ;
wire Xd_0__inst_mult_31_42 ;
wire Xd_0__inst_mult_30_55 ;
wire Xd_0__inst_mult_30_56 ;
wire Xd_0__inst_mult_30_57 ;
wire Xd_0__inst_mult_31_43 ;
wire Xd_0__inst_mult_31_44 ;
wire Xd_0__inst_mult_31_45 ;
wire Xd_0__inst_mult_30_59 ;
wire Xd_0__inst_mult_30_60 ;
wire Xd_0__inst_mult_30_61 ;
wire Xd_0__inst_mult_31_47 ;
wire Xd_0__inst_mult_31_48 ;
wire Xd_0__inst_mult_31_49 ;
wire Xd_0__inst_mult_30_63 ;
wire Xd_0__inst_mult_30_64 ;
wire Xd_0__inst_mult_30_65 ;
wire Xd_0__inst_mult_31_51 ;
wire Xd_0__inst_mult_31_52 ;
wire Xd_0__inst_mult_31_53 ;
wire Xd_0__inst_mult_30_67 ;
wire Xd_0__inst_mult_30_68 ;
wire Xd_0__inst_mult_30_69 ;
wire Xd_0__inst_mult_31_55 ;
wire Xd_0__inst_mult_31_56 ;
wire Xd_0__inst_mult_31_57 ;
wire Xd_0__inst_mult_30_71 ;
wire Xd_0__inst_mult_30_72 ;
wire Xd_0__inst_mult_30_73 ;
wire Xd_0__inst_mult_31_59 ;
wire Xd_0__inst_mult_31_60 ;
wire Xd_0__inst_mult_31_61 ;
wire Xd_0__inst_mult_30_75 ;
wire Xd_0__inst_mult_31_63 ;
wire Xd_0__inst_mult_29_40 ;
wire Xd_0__inst_mult_29_41 ;
wire Xd_0__inst_mult_29_42 ;
wire Xd_0__inst_mult_31_67 ;
wire Xd_0__inst_mult_31_68 ;
wire Xd_0__inst_mult_31_69 ;
wire Xd_0__inst_mult_11_40 ;
wire Xd_0__inst_mult_11_41 ;
wire Xd_0__inst_mult_11_42 ;
wire Xd_0__inst_mult_25_40 ;
wire Xd_0__inst_mult_25_41 ;
wire Xd_0__inst_mult_25_42 ;
wire Xd_0__inst_mult_27_40 ;
wire Xd_0__inst_mult_27_41 ;
wire Xd_0__inst_mult_27_42 ;
wire Xd_0__inst_mult_30_79 ;
wire Xd_0__inst_mult_30_80 ;
wire Xd_0__inst_mult_30_81 ;
wire Xd_0__inst_mult_31_71 ;
wire Xd_0__inst_mult_31_72 ;
wire Xd_0__inst_mult_31_73 ;
wire Xd_0__inst_i17_13_sumout ;
wire Xd_0__inst_i17_14 ;
wire Xd_0__inst_i17_15 ;
wire Xd_0__inst_i17_17_sumout ;
wire Xd_0__inst_i17_18 ;
wire Xd_0__inst_i17_19 ;
wire Xd_0__inst_mult_30_83 ;
wire Xd_0__inst_mult_30_84 ;
wire Xd_0__inst_mult_30_85 ;
wire Xd_0__inst_mult_31_75 ;
wire Xd_0__inst_mult_31_76 ;
wire Xd_0__inst_mult_31_77 ;
wire Xd_0__inst_mult_30_87 ;
wire Xd_0__inst_mult_30_88 ;
wire Xd_0__inst_mult_30_89 ;
wire Xd_0__inst_mult_31_79 ;
wire Xd_0__inst_mult_31_80 ;
wire Xd_0__inst_mult_31_81 ;
wire Xd_0__inst_mult_16_35 ;
wire Xd_0__inst_mult_16_36 ;
wire Xd_0__inst_mult_16_37 ;
wire Xd_0__inst_mult_17_36 ;
wire Xd_0__inst_mult_17_37 ;
wire Xd_0__inst_mult_17_38 ;
wire Xd_0__inst_mult_14_35 ;
wire Xd_0__inst_mult_14_36 ;
wire Xd_0__inst_mult_14_37 ;
wire Xd_0__inst_mult_15_36 ;
wire Xd_0__inst_mult_15_37 ;
wire Xd_0__inst_mult_15_38 ;
wire Xd_0__inst_mult_12_35 ;
wire Xd_0__inst_mult_12_36 ;
wire Xd_0__inst_mult_12_37 ;
wire Xd_0__inst_mult_13_36 ;
wire Xd_0__inst_mult_13_37 ;
wire Xd_0__inst_mult_13_38 ;
wire Xd_0__inst_mult_10_35 ;
wire Xd_0__inst_mult_10_36 ;
wire Xd_0__inst_mult_10_37 ;
wire Xd_0__inst_mult_11_43 ;
wire Xd_0__inst_mult_11_44 ;
wire Xd_0__inst_mult_11_45 ;
wire Xd_0__inst_mult_8_35 ;
wire Xd_0__inst_mult_8_36 ;
wire Xd_0__inst_mult_8_37 ;
wire Xd_0__inst_mult_9_36 ;
wire Xd_0__inst_mult_9_37 ;
wire Xd_0__inst_mult_9_38 ;
wire Xd_0__inst_mult_6_34 ;
wire Xd_0__inst_mult_6_35 ;
wire Xd_0__inst_mult_6_36 ;
wire Xd_0__inst_mult_7_35 ;
wire Xd_0__inst_mult_7_36 ;
wire Xd_0__inst_mult_7_37 ;
wire Xd_0__inst_mult_4_34 ;
wire Xd_0__inst_mult_4_35 ;
wire Xd_0__inst_mult_4_36 ;
wire Xd_0__inst_mult_5_35 ;
wire Xd_0__inst_mult_5_36 ;
wire Xd_0__inst_mult_5_37 ;
wire Xd_0__inst_mult_2_39 ;
wire Xd_0__inst_mult_2_40 ;
wire Xd_0__inst_mult_2_41 ;
wire Xd_0__inst_mult_3_39 ;
wire Xd_0__inst_mult_3_40 ;
wire Xd_0__inst_mult_3_41 ;
wire Xd_0__inst_mult_0_39 ;
wire Xd_0__inst_mult_0_40 ;
wire Xd_0__inst_mult_0_41 ;
wire Xd_0__inst_mult_1_39 ;
wire Xd_0__inst_mult_1_40 ;
wire Xd_0__inst_mult_1_41 ;
wire Xd_0__inst_mult_28_51 ;
wire Xd_0__inst_mult_28_52 ;
wire Xd_0__inst_mult_28_53 ;
wire Xd_0__inst_mult_29_43 ;
wire Xd_0__inst_mult_29_44 ;
wire Xd_0__inst_mult_29_45 ;
wire Xd_0__inst_mult_26_51 ;
wire Xd_0__inst_mult_26_52 ;
wire Xd_0__inst_mult_26_53 ;
wire Xd_0__inst_mult_27_43 ;
wire Xd_0__inst_mult_27_44 ;
wire Xd_0__inst_mult_27_45 ;
wire Xd_0__inst_mult_24_51 ;
wire Xd_0__inst_mult_24_52 ;
wire Xd_0__inst_mult_24_53 ;
wire Xd_0__inst_mult_25_43 ;
wire Xd_0__inst_mult_25_44 ;
wire Xd_0__inst_mult_25_45 ;
wire Xd_0__inst_mult_22_51 ;
wire Xd_0__inst_mult_22_52 ;
wire Xd_0__inst_mult_22_53 ;
wire Xd_0__inst_mult_23_51 ;
wire Xd_0__inst_mult_23_52 ;
wire Xd_0__inst_mult_23_53 ;
wire Xd_0__inst_mult_20_51 ;
wire Xd_0__inst_mult_20_52 ;
wire Xd_0__inst_mult_20_53 ;
wire Xd_0__inst_mult_21_36 ;
wire Xd_0__inst_mult_21_37 ;
wire Xd_0__inst_mult_21_38 ;
wire Xd_0__inst_mult_18_35 ;
wire Xd_0__inst_mult_18_36 ;
wire Xd_0__inst_mult_18_37 ;
wire Xd_0__inst_mult_19_47 ;
wire Xd_0__inst_mult_19_48 ;
wire Xd_0__inst_mult_19_49 ;
wire Xd_0__inst_mult_30_92 ;
wire Xd_0__inst_mult_30_93 ;
wire Xd_0__inst_mult_31_84 ;
wire Xd_0__inst_mult_31_85 ;
wire Xd_0__inst_mult_16_39 ;
wire Xd_0__inst_mult_16_40 ;
wire Xd_0__inst_mult_16_41 ;
wire Xd_0__inst_mult_17_40 ;
wire Xd_0__inst_mult_17_41 ;
wire Xd_0__inst_mult_17_42 ;
wire Xd_0__inst_mult_14_39 ;
wire Xd_0__inst_mult_14_40 ;
wire Xd_0__inst_mult_14_41 ;
wire Xd_0__inst_mult_15_40 ;
wire Xd_0__inst_mult_15_41 ;
wire Xd_0__inst_mult_15_42 ;
wire Xd_0__inst_mult_12_39 ;
wire Xd_0__inst_mult_12_40 ;
wire Xd_0__inst_mult_12_41 ;
wire Xd_0__inst_mult_13_40 ;
wire Xd_0__inst_mult_13_41 ;
wire Xd_0__inst_mult_13_42 ;
wire Xd_0__inst_mult_10_39 ;
wire Xd_0__inst_mult_10_40 ;
wire Xd_0__inst_mult_10_41 ;
wire Xd_0__inst_mult_11_47 ;
wire Xd_0__inst_mult_11_48 ;
wire Xd_0__inst_mult_11_49 ;
wire Xd_0__inst_mult_8_39 ;
wire Xd_0__inst_mult_8_40 ;
wire Xd_0__inst_mult_8_41 ;
wire Xd_0__inst_mult_9_40 ;
wire Xd_0__inst_mult_9_41 ;
wire Xd_0__inst_mult_9_42 ;
wire Xd_0__inst_mult_6_38 ;
wire Xd_0__inst_mult_6_39 ;
wire Xd_0__inst_mult_6_40 ;
wire Xd_0__inst_mult_7_39 ;
wire Xd_0__inst_mult_7_40 ;
wire Xd_0__inst_mult_7_41 ;
wire Xd_0__inst_mult_4_38 ;
wire Xd_0__inst_mult_4_39 ;
wire Xd_0__inst_mult_4_40 ;
wire Xd_0__inst_mult_5_39 ;
wire Xd_0__inst_mult_5_40 ;
wire Xd_0__inst_mult_5_41 ;
wire Xd_0__inst_mult_2_42 ;
wire Xd_0__inst_mult_2_43 ;
wire Xd_0__inst_mult_2_44 ;
wire Xd_0__inst_mult_3_42 ;
wire Xd_0__inst_mult_3_43 ;
wire Xd_0__inst_mult_3_44 ;
wire Xd_0__inst_mult_0_42 ;
wire Xd_0__inst_mult_0_43 ;
wire Xd_0__inst_mult_0_44 ;
wire Xd_0__inst_mult_1_42 ;
wire Xd_0__inst_mult_1_43 ;
wire Xd_0__inst_mult_1_44 ;
wire Xd_0__inst_mult_28_55 ;
wire Xd_0__inst_mult_28_56 ;
wire Xd_0__inst_mult_28_57 ;
wire Xd_0__inst_mult_29_47 ;
wire Xd_0__inst_mult_29_48 ;
wire Xd_0__inst_mult_29_49 ;
wire Xd_0__inst_mult_26_55 ;
wire Xd_0__inst_mult_26_56 ;
wire Xd_0__inst_mult_26_57 ;
wire Xd_0__inst_mult_27_47 ;
wire Xd_0__inst_mult_27_48 ;
wire Xd_0__inst_mult_27_49 ;
wire Xd_0__inst_mult_24_55 ;
wire Xd_0__inst_mult_24_56 ;
wire Xd_0__inst_mult_24_57 ;
wire Xd_0__inst_mult_25_47 ;
wire Xd_0__inst_mult_25_48 ;
wire Xd_0__inst_mult_25_49 ;
wire Xd_0__inst_mult_22_55 ;
wire Xd_0__inst_mult_22_56 ;
wire Xd_0__inst_mult_22_57 ;
wire Xd_0__inst_mult_23_55 ;
wire Xd_0__inst_mult_23_56 ;
wire Xd_0__inst_mult_23_57 ;
wire Xd_0__inst_mult_20_55 ;
wire Xd_0__inst_mult_20_56 ;
wire Xd_0__inst_mult_20_57 ;
wire Xd_0__inst_mult_21_40 ;
wire Xd_0__inst_mult_21_41 ;
wire Xd_0__inst_mult_21_42 ;
wire Xd_0__inst_mult_18_39 ;
wire Xd_0__inst_mult_18_40 ;
wire Xd_0__inst_mult_18_41 ;
wire Xd_0__inst_mult_19_51 ;
wire Xd_0__inst_mult_19_52 ;
wire Xd_0__inst_mult_19_53 ;
wire Xd_0__inst_mult_16_42 ;
wire Xd_0__inst_mult_16_43 ;
wire Xd_0__inst_mult_16_44 ;
wire Xd_0__inst_mult_17_43 ;
wire Xd_0__inst_mult_17_44 ;
wire Xd_0__inst_mult_17_45 ;
wire Xd_0__inst_mult_14_42 ;
wire Xd_0__inst_mult_14_43 ;
wire Xd_0__inst_mult_14_44 ;
wire Xd_0__inst_mult_15_43 ;
wire Xd_0__inst_mult_15_44 ;
wire Xd_0__inst_mult_15_45 ;
wire Xd_0__inst_mult_12_42 ;
wire Xd_0__inst_mult_12_43 ;
wire Xd_0__inst_mult_12_44 ;
wire Xd_0__inst_mult_13_43 ;
wire Xd_0__inst_mult_13_44 ;
wire Xd_0__inst_mult_13_45 ;
wire Xd_0__inst_mult_10_42 ;
wire Xd_0__inst_mult_10_43 ;
wire Xd_0__inst_mult_10_44 ;
wire Xd_0__inst_mult_11_51 ;
wire Xd_0__inst_mult_11_52 ;
wire Xd_0__inst_mult_11_53 ;
wire Xd_0__inst_mult_8_42 ;
wire Xd_0__inst_mult_8_43 ;
wire Xd_0__inst_mult_8_44 ;
wire Xd_0__inst_mult_9_43 ;
wire Xd_0__inst_mult_9_44 ;
wire Xd_0__inst_mult_9_45 ;
wire Xd_0__inst_mult_6_41 ;
wire Xd_0__inst_mult_6_42 ;
wire Xd_0__inst_mult_6_43 ;
wire Xd_0__inst_mult_7_42 ;
wire Xd_0__inst_mult_7_43 ;
wire Xd_0__inst_mult_7_44 ;
wire Xd_0__inst_mult_4_41 ;
wire Xd_0__inst_mult_4_42 ;
wire Xd_0__inst_mult_4_43 ;
wire Xd_0__inst_mult_5_42 ;
wire Xd_0__inst_mult_5_43 ;
wire Xd_0__inst_mult_5_44 ;
wire Xd_0__inst_mult_2_46 ;
wire Xd_0__inst_mult_2_47 ;
wire Xd_0__inst_mult_2_48 ;
wire Xd_0__inst_mult_3_46 ;
wire Xd_0__inst_mult_3_47 ;
wire Xd_0__inst_mult_3_48 ;
wire Xd_0__inst_mult_0_46 ;
wire Xd_0__inst_mult_0_47 ;
wire Xd_0__inst_mult_0_48 ;
wire Xd_0__inst_mult_1_46 ;
wire Xd_0__inst_mult_1_47 ;
wire Xd_0__inst_mult_1_48 ;
wire Xd_0__inst_mult_28_59 ;
wire Xd_0__inst_mult_28_60 ;
wire Xd_0__inst_mult_28_61 ;
wire Xd_0__inst_mult_29_51 ;
wire Xd_0__inst_mult_29_52 ;
wire Xd_0__inst_mult_29_53 ;
wire Xd_0__inst_mult_26_59 ;
wire Xd_0__inst_mult_26_60 ;
wire Xd_0__inst_mult_26_61 ;
wire Xd_0__inst_mult_27_51 ;
wire Xd_0__inst_mult_27_52 ;
wire Xd_0__inst_mult_27_53 ;
wire Xd_0__inst_mult_24_59 ;
wire Xd_0__inst_mult_24_60 ;
wire Xd_0__inst_mult_24_61 ;
wire Xd_0__inst_mult_25_51 ;
wire Xd_0__inst_mult_25_52 ;
wire Xd_0__inst_mult_25_53 ;
wire Xd_0__inst_mult_22_59 ;
wire Xd_0__inst_mult_22_60 ;
wire Xd_0__inst_mult_22_61 ;
wire Xd_0__inst_mult_23_59 ;
wire Xd_0__inst_mult_23_60 ;
wire Xd_0__inst_mult_23_61 ;
wire Xd_0__inst_mult_20_59 ;
wire Xd_0__inst_mult_20_60 ;
wire Xd_0__inst_mult_20_61 ;
wire Xd_0__inst_mult_21_43 ;
wire Xd_0__inst_mult_21_44 ;
wire Xd_0__inst_mult_21_45 ;
wire Xd_0__inst_mult_18_42 ;
wire Xd_0__inst_mult_18_43 ;
wire Xd_0__inst_mult_18_44 ;
wire Xd_0__inst_mult_19_55 ;
wire Xd_0__inst_mult_19_56 ;
wire Xd_0__inst_mult_19_57 ;
wire Xd_0__inst_mult_16_46 ;
wire Xd_0__inst_mult_16_47 ;
wire Xd_0__inst_mult_16_48 ;
wire Xd_0__inst_mult_17_47 ;
wire Xd_0__inst_mult_17_48 ;
wire Xd_0__inst_mult_17_49 ;
wire Xd_0__inst_mult_14_46 ;
wire Xd_0__inst_mult_14_47 ;
wire Xd_0__inst_mult_14_48 ;
wire Xd_0__inst_mult_15_47 ;
wire Xd_0__inst_mult_15_48 ;
wire Xd_0__inst_mult_15_49 ;
wire Xd_0__inst_mult_12_46 ;
wire Xd_0__inst_mult_12_47 ;
wire Xd_0__inst_mult_12_48 ;
wire Xd_0__inst_mult_13_47 ;
wire Xd_0__inst_mult_13_48 ;
wire Xd_0__inst_mult_13_49 ;
wire Xd_0__inst_mult_10_46 ;
wire Xd_0__inst_mult_10_47 ;
wire Xd_0__inst_mult_10_48 ;
wire Xd_0__inst_mult_11_55 ;
wire Xd_0__inst_mult_11_56 ;
wire Xd_0__inst_mult_11_57 ;
wire Xd_0__inst_mult_8_46 ;
wire Xd_0__inst_mult_8_47 ;
wire Xd_0__inst_mult_8_48 ;
wire Xd_0__inst_mult_9_47 ;
wire Xd_0__inst_mult_9_48 ;
wire Xd_0__inst_mult_9_49 ;
wire Xd_0__inst_mult_6_45 ;
wire Xd_0__inst_mult_6_46 ;
wire Xd_0__inst_mult_6_47 ;
wire Xd_0__inst_mult_7_46 ;
wire Xd_0__inst_mult_7_47 ;
wire Xd_0__inst_mult_7_48 ;
wire Xd_0__inst_mult_4_45 ;
wire Xd_0__inst_mult_4_46 ;
wire Xd_0__inst_mult_4_47 ;
wire Xd_0__inst_mult_5_46 ;
wire Xd_0__inst_mult_5_47 ;
wire Xd_0__inst_mult_5_48 ;
wire Xd_0__inst_mult_2_50 ;
wire Xd_0__inst_mult_2_51 ;
wire Xd_0__inst_mult_2_52 ;
wire Xd_0__inst_mult_3_50 ;
wire Xd_0__inst_mult_3_51 ;
wire Xd_0__inst_mult_3_52 ;
wire Xd_0__inst_mult_0_50 ;
wire Xd_0__inst_mult_0_51 ;
wire Xd_0__inst_mult_0_52 ;
wire Xd_0__inst_mult_1_50 ;
wire Xd_0__inst_mult_1_51 ;
wire Xd_0__inst_mult_1_52 ;
wire Xd_0__inst_mult_28_63 ;
wire Xd_0__inst_mult_28_64 ;
wire Xd_0__inst_mult_28_65 ;
wire Xd_0__inst_mult_29_55 ;
wire Xd_0__inst_mult_29_56 ;
wire Xd_0__inst_mult_29_57 ;
wire Xd_0__inst_mult_26_63 ;
wire Xd_0__inst_mult_26_64 ;
wire Xd_0__inst_mult_26_65 ;
wire Xd_0__inst_mult_27_55 ;
wire Xd_0__inst_mult_27_56 ;
wire Xd_0__inst_mult_27_57 ;
wire Xd_0__inst_mult_24_63 ;
wire Xd_0__inst_mult_24_64 ;
wire Xd_0__inst_mult_24_65 ;
wire Xd_0__inst_mult_25_55 ;
wire Xd_0__inst_mult_25_56 ;
wire Xd_0__inst_mult_25_57 ;
wire Xd_0__inst_mult_22_63 ;
wire Xd_0__inst_mult_22_64 ;
wire Xd_0__inst_mult_22_65 ;
wire Xd_0__inst_mult_23_63 ;
wire Xd_0__inst_mult_23_64 ;
wire Xd_0__inst_mult_23_65 ;
wire Xd_0__inst_mult_20_63 ;
wire Xd_0__inst_mult_20_64 ;
wire Xd_0__inst_mult_20_65 ;
wire Xd_0__inst_mult_21_47 ;
wire Xd_0__inst_mult_21_48 ;
wire Xd_0__inst_mult_21_49 ;
wire Xd_0__inst_mult_18_46 ;
wire Xd_0__inst_mult_18_47 ;
wire Xd_0__inst_mult_18_48 ;
wire Xd_0__inst_mult_19_59 ;
wire Xd_0__inst_mult_19_60 ;
wire Xd_0__inst_mult_19_61 ;
wire Xd_0__inst_mult_16_50 ;
wire Xd_0__inst_mult_16_51 ;
wire Xd_0__inst_mult_16_52 ;
wire Xd_0__inst_mult_17_51 ;
wire Xd_0__inst_mult_17_52 ;
wire Xd_0__inst_mult_17_53 ;
wire Xd_0__inst_mult_14_50 ;
wire Xd_0__inst_mult_14_51 ;
wire Xd_0__inst_mult_14_52 ;
wire Xd_0__inst_mult_15_51 ;
wire Xd_0__inst_mult_15_52 ;
wire Xd_0__inst_mult_15_53 ;
wire Xd_0__inst_mult_12_50 ;
wire Xd_0__inst_mult_12_51 ;
wire Xd_0__inst_mult_12_52 ;
wire Xd_0__inst_mult_13_51 ;
wire Xd_0__inst_mult_13_52 ;
wire Xd_0__inst_mult_13_53 ;
wire Xd_0__inst_mult_10_50 ;
wire Xd_0__inst_mult_10_51 ;
wire Xd_0__inst_mult_10_52 ;
wire Xd_0__inst_mult_11_59 ;
wire Xd_0__inst_mult_11_60 ;
wire Xd_0__inst_mult_11_61 ;
wire Xd_0__inst_mult_8_50 ;
wire Xd_0__inst_mult_8_51 ;
wire Xd_0__inst_mult_8_52 ;
wire Xd_0__inst_mult_9_51 ;
wire Xd_0__inst_mult_9_52 ;
wire Xd_0__inst_mult_9_53 ;
wire Xd_0__inst_mult_6_49 ;
wire Xd_0__inst_mult_6_50 ;
wire Xd_0__inst_mult_6_51 ;
wire Xd_0__inst_mult_7_50 ;
wire Xd_0__inst_mult_7_51 ;
wire Xd_0__inst_mult_7_52 ;
wire Xd_0__inst_mult_4_49 ;
wire Xd_0__inst_mult_4_50 ;
wire Xd_0__inst_mult_4_51 ;
wire Xd_0__inst_mult_5_50 ;
wire Xd_0__inst_mult_5_51 ;
wire Xd_0__inst_mult_5_52 ;
wire Xd_0__inst_mult_2_54 ;
wire Xd_0__inst_mult_2_55 ;
wire Xd_0__inst_mult_2_56 ;
wire Xd_0__inst_mult_3_54 ;
wire Xd_0__inst_mult_3_55 ;
wire Xd_0__inst_mult_3_56 ;
wire Xd_0__inst_mult_0_54 ;
wire Xd_0__inst_mult_0_55 ;
wire Xd_0__inst_mult_0_56 ;
wire Xd_0__inst_mult_1_54 ;
wire Xd_0__inst_mult_1_55 ;
wire Xd_0__inst_mult_1_56 ;
wire Xd_0__inst_mult_28_67 ;
wire Xd_0__inst_mult_28_68 ;
wire Xd_0__inst_mult_28_69 ;
wire Xd_0__inst_mult_29_59 ;
wire Xd_0__inst_mult_29_60 ;
wire Xd_0__inst_mult_29_61 ;
wire Xd_0__inst_mult_26_67 ;
wire Xd_0__inst_mult_26_68 ;
wire Xd_0__inst_mult_26_69 ;
wire Xd_0__inst_mult_27_59 ;
wire Xd_0__inst_mult_27_60 ;
wire Xd_0__inst_mult_27_61 ;
wire Xd_0__inst_mult_24_67 ;
wire Xd_0__inst_mult_24_68 ;
wire Xd_0__inst_mult_24_69 ;
wire Xd_0__inst_mult_25_59 ;
wire Xd_0__inst_mult_25_60 ;
wire Xd_0__inst_mult_25_61 ;
wire Xd_0__inst_mult_22_67 ;
wire Xd_0__inst_mult_22_68 ;
wire Xd_0__inst_mult_22_69 ;
wire Xd_0__inst_mult_23_67 ;
wire Xd_0__inst_mult_23_68 ;
wire Xd_0__inst_mult_23_69 ;
wire Xd_0__inst_mult_20_67 ;
wire Xd_0__inst_mult_20_68 ;
wire Xd_0__inst_mult_20_69 ;
wire Xd_0__inst_mult_21_51 ;
wire Xd_0__inst_mult_21_52 ;
wire Xd_0__inst_mult_21_53 ;
wire Xd_0__inst_mult_18_50 ;
wire Xd_0__inst_mult_18_51 ;
wire Xd_0__inst_mult_18_52 ;
wire Xd_0__inst_mult_19_63 ;
wire Xd_0__inst_mult_19_64 ;
wire Xd_0__inst_mult_19_65 ;
wire Xd_0__inst_mult_16_54 ;
wire Xd_0__inst_mult_16_55 ;
wire Xd_0__inst_mult_16_56 ;
wire Xd_0__inst_mult_17_55 ;
wire Xd_0__inst_mult_17_56 ;
wire Xd_0__inst_mult_17_57 ;
wire Xd_0__inst_mult_14_54 ;
wire Xd_0__inst_mult_14_55 ;
wire Xd_0__inst_mult_14_56 ;
wire Xd_0__inst_mult_15_55 ;
wire Xd_0__inst_mult_15_56 ;
wire Xd_0__inst_mult_15_57 ;
wire Xd_0__inst_mult_12_54 ;
wire Xd_0__inst_mult_12_55 ;
wire Xd_0__inst_mult_12_56 ;
wire Xd_0__inst_mult_13_55 ;
wire Xd_0__inst_mult_13_56 ;
wire Xd_0__inst_mult_13_57 ;
wire Xd_0__inst_mult_10_54 ;
wire Xd_0__inst_mult_10_55 ;
wire Xd_0__inst_mult_10_56 ;
wire Xd_0__inst_mult_11_63 ;
wire Xd_0__inst_mult_11_64 ;
wire Xd_0__inst_mult_11_65 ;
wire Xd_0__inst_mult_8_54 ;
wire Xd_0__inst_mult_8_55 ;
wire Xd_0__inst_mult_8_56 ;
wire Xd_0__inst_mult_9_55 ;
wire Xd_0__inst_mult_9_56 ;
wire Xd_0__inst_mult_9_57 ;
wire Xd_0__inst_mult_6_53 ;
wire Xd_0__inst_mult_6_54 ;
wire Xd_0__inst_mult_6_55 ;
wire Xd_0__inst_mult_7_54 ;
wire Xd_0__inst_mult_7_55 ;
wire Xd_0__inst_mult_7_56 ;
wire Xd_0__inst_mult_4_53 ;
wire Xd_0__inst_mult_4_54 ;
wire Xd_0__inst_mult_4_55 ;
wire Xd_0__inst_mult_5_54 ;
wire Xd_0__inst_mult_5_55 ;
wire Xd_0__inst_mult_5_56 ;
wire Xd_0__inst_mult_2_58 ;
wire Xd_0__inst_mult_2_59 ;
wire Xd_0__inst_mult_2_60 ;
wire Xd_0__inst_mult_3_58 ;
wire Xd_0__inst_mult_3_59 ;
wire Xd_0__inst_mult_3_60 ;
wire Xd_0__inst_mult_0_58 ;
wire Xd_0__inst_mult_0_59 ;
wire Xd_0__inst_mult_0_60 ;
wire Xd_0__inst_mult_1_58 ;
wire Xd_0__inst_mult_1_59 ;
wire Xd_0__inst_mult_1_60 ;
wire Xd_0__inst_mult_28_71 ;
wire Xd_0__inst_mult_28_72 ;
wire Xd_0__inst_mult_28_73 ;
wire Xd_0__inst_mult_29_63 ;
wire Xd_0__inst_mult_29_64 ;
wire Xd_0__inst_mult_29_65 ;
wire Xd_0__inst_mult_26_71 ;
wire Xd_0__inst_mult_26_72 ;
wire Xd_0__inst_mult_26_73 ;
wire Xd_0__inst_mult_27_63 ;
wire Xd_0__inst_mult_27_64 ;
wire Xd_0__inst_mult_27_65 ;
wire Xd_0__inst_mult_24_71 ;
wire Xd_0__inst_mult_24_72 ;
wire Xd_0__inst_mult_24_73 ;
wire Xd_0__inst_mult_25_63 ;
wire Xd_0__inst_mult_25_64 ;
wire Xd_0__inst_mult_25_65 ;
wire Xd_0__inst_mult_22_71 ;
wire Xd_0__inst_mult_22_72 ;
wire Xd_0__inst_mult_22_73 ;
wire Xd_0__inst_mult_23_71 ;
wire Xd_0__inst_mult_23_72 ;
wire Xd_0__inst_mult_23_73 ;
wire Xd_0__inst_mult_20_71 ;
wire Xd_0__inst_mult_20_72 ;
wire Xd_0__inst_mult_20_73 ;
wire Xd_0__inst_mult_21_55 ;
wire Xd_0__inst_mult_21_56 ;
wire Xd_0__inst_mult_21_57 ;
wire Xd_0__inst_mult_18_54 ;
wire Xd_0__inst_mult_18_55 ;
wire Xd_0__inst_mult_18_56 ;
wire Xd_0__inst_mult_19_67 ;
wire Xd_0__inst_mult_19_68 ;
wire Xd_0__inst_mult_19_69 ;
wire Xd_0__inst_mult_17_59 ;
wire Xd_0__inst_mult_17_60 ;
wire Xd_0__inst_mult_17_61 ;
wire Xd_0__inst_mult_17_63 ;
wire Xd_0__inst_mult_15_59 ;
wire Xd_0__inst_mult_15_60 ;
wire Xd_0__inst_mult_15_61 ;
wire Xd_0__inst_mult_15_63 ;
wire Xd_0__inst_mult_13_59 ;
wire Xd_0__inst_mult_13_60 ;
wire Xd_0__inst_mult_13_61 ;
wire Xd_0__inst_mult_13_63 ;
wire Xd_0__inst_mult_21_59 ;
wire Xd_0__inst_mult_21_60 ;
wire Xd_0__inst_mult_21_61 ;
wire Xd_0__inst_mult_11_67 ;
wire Xd_0__inst_mult_9_59 ;
wire Xd_0__inst_mult_9_60 ;
wire Xd_0__inst_mult_9_61 ;
wire Xd_0__inst_mult_9_63 ;
wire Xd_0__inst_mult_7_58 ;
wire Xd_0__inst_mult_7_59 ;
wire Xd_0__inst_mult_7_60 ;
wire Xd_0__inst_mult_7_62 ;
wire Xd_0__inst_mult_5_58 ;
wire Xd_0__inst_mult_5_59 ;
wire Xd_0__inst_mult_5_60 ;
wire Xd_0__inst_mult_5_62 ;
wire Xd_0__inst_mult_2_62 ;
wire Xd_0__inst_mult_3_62 ;
wire Xd_0__inst_mult_0_62 ;
wire Xd_0__inst_mult_1_62 ;
wire Xd_0__inst_mult_28_75 ;
wire Xd_0__inst_mult_29_67 ;
wire Xd_0__inst_mult_26_75 ;
wire Xd_0__inst_mult_27_67 ;
wire Xd_0__inst_mult_24_75 ;
wire Xd_0__inst_mult_25_67 ;
wire Xd_0__inst_mult_22_75 ;
wire Xd_0__inst_mult_23_75 ;
wire Xd_0__inst_mult_20_75 ;
wire Xd_0__inst_mult_21_63 ;
wire Xd_0__inst_mult_19_71 ;
wire Xd_0__inst_mult_19_72 ;
wire Xd_0__inst_mult_19_73 ;
wire Xd_0__inst_mult_19_75 ;
wire Xd_0__inst_mult_16_58 ;
wire Xd_0__inst_mult_16_59 ;
wire Xd_0__inst_mult_16_60 ;
wire Xd_0__inst_mult_17_67 ;
wire Xd_0__inst_mult_17_68 ;
wire Xd_0__inst_mult_17_69 ;
wire Xd_0__inst_i17_21_sumout ;
wire Xd_0__inst_i17_22 ;
wire Xd_0__inst_i17_23 ;
wire Xd_0__inst_mult_14_58 ;
wire Xd_0__inst_mult_14_59 ;
wire Xd_0__inst_mult_14_60 ;
wire Xd_0__inst_mult_15_67 ;
wire Xd_0__inst_mult_15_68 ;
wire Xd_0__inst_mult_15_69 ;
wire Xd_0__inst_i17_25_sumout ;
wire Xd_0__inst_i17_26 ;
wire Xd_0__inst_i17_27 ;
wire Xd_0__inst_i17_29_sumout ;
wire Xd_0__inst_i17_30 ;
wire Xd_0__inst_i17_31 ;
wire Xd_0__inst_mult_12_58 ;
wire Xd_0__inst_mult_12_59 ;
wire Xd_0__inst_mult_12_60 ;
wire Xd_0__inst_mult_13_67 ;
wire Xd_0__inst_mult_13_68 ;
wire Xd_0__inst_mult_13_69 ;
wire Xd_0__inst_i17_33_sumout ;
wire Xd_0__inst_i17_34 ;
wire Xd_0__inst_i17_35 ;
wire Xd_0__inst_i17_37_sumout ;
wire Xd_0__inst_i17_38 ;
wire Xd_0__inst_i17_39 ;
wire Xd_0__inst_mult_29_71 ;
wire Xd_0__inst_mult_29_72 ;
wire Xd_0__inst_mult_29_73 ;
wire Xd_0__inst_mult_10_58 ;
wire Xd_0__inst_mult_10_59 ;
wire Xd_0__inst_mult_10_60 ;
wire Xd_0__inst_mult_11_71 ;
wire Xd_0__inst_mult_11_72 ;
wire Xd_0__inst_mult_11_73 ;
wire Xd_0__inst_i17_41_sumout ;
wire Xd_0__inst_i17_42 ;
wire Xd_0__inst_i17_43 ;
wire Xd_0__inst_mult_8_58 ;
wire Xd_0__inst_mult_8_59 ;
wire Xd_0__inst_mult_8_60 ;
wire Xd_0__inst_mult_9_67 ;
wire Xd_0__inst_mult_9_68 ;
wire Xd_0__inst_mult_9_69 ;
wire Xd_0__inst_i17_45_sumout ;
wire Xd_0__inst_i17_46 ;
wire Xd_0__inst_i17_47 ;
wire Xd_0__inst_i17_49_sumout ;
wire Xd_0__inst_i17_50 ;
wire Xd_0__inst_i17_51 ;
wire Xd_0__inst_mult_6_57 ;
wire Xd_0__inst_mult_6_58 ;
wire Xd_0__inst_mult_6_59 ;
wire Xd_0__inst_mult_7_66 ;
wire Xd_0__inst_mult_7_67 ;
wire Xd_0__inst_mult_7_68 ;
wire Xd_0__inst_i17_53_sumout ;
wire Xd_0__inst_i17_54 ;
wire Xd_0__inst_i17_55 ;
wire Xd_0__inst_i17_57_sumout ;
wire Xd_0__inst_i17_58 ;
wire Xd_0__inst_i17_59 ;
wire Xd_0__inst_mult_31_87 ;
wire Xd_0__inst_mult_31_88 ;
wire Xd_0__inst_mult_31_89 ;
wire Xd_0__inst_mult_4_57 ;
wire Xd_0__inst_mult_4_58 ;
wire Xd_0__inst_mult_4_59 ;
wire Xd_0__inst_mult_5_66 ;
wire Xd_0__inst_mult_5_67 ;
wire Xd_0__inst_mult_5_68 ;
wire Xd_0__inst_i17_61_sumout ;
wire Xd_0__inst_i17_62 ;
wire Xd_0__inst_i17_63 ;
wire Xd_0__inst_i17_65_sumout ;
wire Xd_0__inst_i17_66 ;
wire Xd_0__inst_i17_67 ;
wire Xd_0__inst_mult_2_66 ;
wire Xd_0__inst_mult_2_67 ;
wire Xd_0__inst_mult_2_68 ;
wire Xd_0__inst_mult_3_66 ;
wire Xd_0__inst_mult_3_67 ;
wire Xd_0__inst_mult_3_68 ;
wire Xd_0__inst_i17_69_sumout ;
wire Xd_0__inst_i17_70 ;
wire Xd_0__inst_i17_71 ;
wire Xd_0__inst_i17_73_sumout ;
wire Xd_0__inst_i17_74 ;
wire Xd_0__inst_i17_75 ;
wire Xd_0__inst_mult_0_66 ;
wire Xd_0__inst_mult_0_67 ;
wire Xd_0__inst_mult_0_68 ;
wire Xd_0__inst_mult_1_66 ;
wire Xd_0__inst_mult_1_67 ;
wire Xd_0__inst_mult_1_68 ;
wire Xd_0__inst_i17_77_sumout ;
wire Xd_0__inst_i17_78 ;
wire Xd_0__inst_i17_79 ;
wire Xd_0__inst_i17_81_sumout ;
wire Xd_0__inst_i17_82 ;
wire Xd_0__inst_i17_83 ;
wire Xd_0__inst_mult_11_75 ;
wire Xd_0__inst_mult_11_76 ;
wire Xd_0__inst_mult_11_77 ;
wire Xd_0__inst_mult_28_79 ;
wire Xd_0__inst_mult_28_80 ;
wire Xd_0__inst_mult_28_81 ;
wire Xd_0__inst_mult_29_75 ;
wire Xd_0__inst_mult_29_76 ;
wire Xd_0__inst_mult_29_77 ;
wire Xd_0__inst_i17_85_sumout ;
wire Xd_0__inst_i17_86 ;
wire Xd_0__inst_i17_87 ;
wire Xd_0__inst_i17_89_sumout ;
wire Xd_0__inst_i17_90 ;
wire Xd_0__inst_i17_91 ;
wire Xd_0__inst_mult_26_79 ;
wire Xd_0__inst_mult_26_80 ;
wire Xd_0__inst_mult_26_81 ;
wire Xd_0__inst_mult_27_71 ;
wire Xd_0__inst_mult_27_72 ;
wire Xd_0__inst_mult_27_73 ;
wire Xd_0__inst_i17_93_sumout ;
wire Xd_0__inst_i17_94 ;
wire Xd_0__inst_i17_95 ;
wire Xd_0__inst_mult_24_79 ;
wire Xd_0__inst_mult_24_80 ;
wire Xd_0__inst_mult_24_81 ;
wire Xd_0__inst_mult_25_71 ;
wire Xd_0__inst_mult_25_72 ;
wire Xd_0__inst_mult_25_73 ;
wire Xd_0__inst_i17_97_sumout ;
wire Xd_0__inst_i17_98 ;
wire Xd_0__inst_i17_99 ;
wire Xd_0__inst_i17_101_sumout ;
wire Xd_0__inst_i17_102 ;
wire Xd_0__inst_i17_103 ;
wire Xd_0__inst_mult_25_75 ;
wire Xd_0__inst_mult_25_76 ;
wire Xd_0__inst_mult_25_77 ;
wire Xd_0__inst_mult_22_79 ;
wire Xd_0__inst_mult_22_80 ;
wire Xd_0__inst_mult_22_81 ;
wire Xd_0__inst_mult_23_79 ;
wire Xd_0__inst_mult_23_80 ;
wire Xd_0__inst_mult_23_81 ;
wire Xd_0__inst_i17_105_sumout ;
wire Xd_0__inst_i17_106 ;
wire Xd_0__inst_i17_107 ;
wire Xd_0__inst_i17_109_sumout ;
wire Xd_0__inst_i17_110 ;
wire Xd_0__inst_i17_111 ;
wire Xd_0__inst_mult_20_79 ;
wire Xd_0__inst_mult_20_80 ;
wire Xd_0__inst_mult_20_81 ;
wire Xd_0__inst_mult_21_67 ;
wire Xd_0__inst_mult_21_68 ;
wire Xd_0__inst_mult_21_69 ;
wire Xd_0__inst_i17_113_sumout ;
wire Xd_0__inst_i17_114 ;
wire Xd_0__inst_i17_115 ;
wire Xd_0__inst_i17_117_sumout ;
wire Xd_0__inst_i17_118 ;
wire Xd_0__inst_i17_119 ;
wire Xd_0__inst_mult_18_58 ;
wire Xd_0__inst_mult_18_59 ;
wire Xd_0__inst_mult_18_60 ;
wire Xd_0__inst_mult_19_79 ;
wire Xd_0__inst_mult_19_80 ;
wire Xd_0__inst_mult_19_81 ;
wire Xd_0__inst_i17_121_sumout ;
wire Xd_0__inst_i17_122 ;
wire Xd_0__inst_i17_123 ;
wire Xd_0__inst_i17_125_sumout ;
wire Xd_0__inst_i17_126 ;
wire Xd_0__inst_i17_127 ;
wire Xd_0__inst_mult_27_75 ;
wire Xd_0__inst_mult_27_76 ;
wire Xd_0__inst_mult_27_77 ;
wire Xd_0__inst_mult_30_95 ;
wire Xd_0__inst_mult_30_96 ;
wire Xd_0__inst_mult_30_97 ;
wire Xd_0__inst_mult_16_62 ;
wire Xd_0__inst_mult_16_63 ;
wire Xd_0__inst_mult_16_64 ;
wire Xd_0__inst_mult_17_71 ;
wire Xd_0__inst_mult_17_72 ;
wire Xd_0__inst_mult_17_73 ;
wire Xd_0__inst_mult_14_62 ;
wire Xd_0__inst_mult_14_63 ;
wire Xd_0__inst_mult_14_64 ;
wire Xd_0__inst_mult_15_71 ;
wire Xd_0__inst_mult_15_72 ;
wire Xd_0__inst_mult_15_73 ;
wire Xd_0__inst_mult_12_62 ;
wire Xd_0__inst_mult_12_63 ;
wire Xd_0__inst_mult_12_64 ;
wire Xd_0__inst_mult_13_71 ;
wire Xd_0__inst_mult_13_72 ;
wire Xd_0__inst_mult_13_73 ;
wire Xd_0__inst_mult_10_62 ;
wire Xd_0__inst_mult_10_63 ;
wire Xd_0__inst_mult_10_64 ;
wire Xd_0__inst_mult_11_79 ;
wire Xd_0__inst_mult_11_80 ;
wire Xd_0__inst_mult_11_81 ;
wire Xd_0__inst_mult_8_62 ;
wire Xd_0__inst_mult_8_63 ;
wire Xd_0__inst_mult_8_64 ;
wire Xd_0__inst_mult_9_71 ;
wire Xd_0__inst_mult_9_72 ;
wire Xd_0__inst_mult_9_73 ;
wire Xd_0__inst_mult_6_61 ;
wire Xd_0__inst_mult_6_62 ;
wire Xd_0__inst_mult_6_63 ;
wire Xd_0__inst_mult_7_70 ;
wire Xd_0__inst_mult_7_71 ;
wire Xd_0__inst_mult_7_72 ;
wire Xd_0__inst_mult_4_61 ;
wire Xd_0__inst_mult_4_62 ;
wire Xd_0__inst_mult_4_63 ;
wire Xd_0__inst_mult_5_70 ;
wire Xd_0__inst_mult_5_71 ;
wire Xd_0__inst_mult_5_72 ;
wire Xd_0__inst_mult_2_70 ;
wire Xd_0__inst_mult_2_71 ;
wire Xd_0__inst_mult_2_72 ;
wire Xd_0__inst_mult_3_70 ;
wire Xd_0__inst_mult_3_71 ;
wire Xd_0__inst_mult_3_72 ;
wire Xd_0__inst_mult_0_70 ;
wire Xd_0__inst_mult_0_71 ;
wire Xd_0__inst_mult_0_72 ;
wire Xd_0__inst_mult_1_70 ;
wire Xd_0__inst_mult_1_71 ;
wire Xd_0__inst_mult_1_72 ;
wire Xd_0__inst_mult_28_83 ;
wire Xd_0__inst_mult_28_84 ;
wire Xd_0__inst_mult_28_85 ;
wire Xd_0__inst_mult_29_79 ;
wire Xd_0__inst_mult_29_80 ;
wire Xd_0__inst_mult_29_81 ;
wire Xd_0__inst_mult_26_83 ;
wire Xd_0__inst_mult_26_84 ;
wire Xd_0__inst_mult_26_85 ;
wire Xd_0__inst_mult_27_79 ;
wire Xd_0__inst_mult_27_80 ;
wire Xd_0__inst_mult_27_81 ;
wire Xd_0__inst_mult_24_83 ;
wire Xd_0__inst_mult_24_84 ;
wire Xd_0__inst_mult_24_85 ;
wire Xd_0__inst_mult_25_79 ;
wire Xd_0__inst_mult_25_80 ;
wire Xd_0__inst_mult_25_81 ;
wire Xd_0__inst_mult_22_83 ;
wire Xd_0__inst_mult_22_84 ;
wire Xd_0__inst_mult_22_85 ;
wire Xd_0__inst_mult_23_83 ;
wire Xd_0__inst_mult_23_84 ;
wire Xd_0__inst_mult_23_85 ;
wire Xd_0__inst_mult_20_83 ;
wire Xd_0__inst_mult_20_84 ;
wire Xd_0__inst_mult_20_85 ;
wire Xd_0__inst_mult_21_71 ;
wire Xd_0__inst_mult_21_72 ;
wire Xd_0__inst_mult_21_73 ;
wire Xd_0__inst_mult_18_62 ;
wire Xd_0__inst_mult_18_63 ;
wire Xd_0__inst_mult_18_64 ;
wire Xd_0__inst_mult_19_83 ;
wire Xd_0__inst_mult_19_84 ;
wire Xd_0__inst_mult_19_85 ;
wire Xd_0__inst_mult_16_66 ;
wire Xd_0__inst_mult_16_67 ;
wire Xd_0__inst_mult_16_68 ;
wire Xd_0__inst_mult_17_75 ;
wire Xd_0__inst_mult_17_76 ;
wire Xd_0__inst_mult_17_77 ;
wire Xd_0__inst_mult_14_66 ;
wire Xd_0__inst_mult_14_67 ;
wire Xd_0__inst_mult_14_68 ;
wire Xd_0__inst_mult_15_75 ;
wire Xd_0__inst_mult_15_76 ;
wire Xd_0__inst_mult_15_77 ;
wire Xd_0__inst_mult_12_66 ;
wire Xd_0__inst_mult_12_67 ;
wire Xd_0__inst_mult_12_68 ;
wire Xd_0__inst_mult_13_75 ;
wire Xd_0__inst_mult_13_76 ;
wire Xd_0__inst_mult_13_77 ;
wire Xd_0__inst_mult_10_66 ;
wire Xd_0__inst_mult_10_67 ;
wire Xd_0__inst_mult_10_68 ;
wire Xd_0__inst_mult_11_83 ;
wire Xd_0__inst_mult_11_84 ;
wire Xd_0__inst_mult_11_85 ;
wire Xd_0__inst_mult_8_66 ;
wire Xd_0__inst_mult_8_67 ;
wire Xd_0__inst_mult_8_68 ;
wire Xd_0__inst_mult_9_75 ;
wire Xd_0__inst_mult_9_76 ;
wire Xd_0__inst_mult_9_77 ;
wire Xd_0__inst_mult_6_65 ;
wire Xd_0__inst_mult_6_66 ;
wire Xd_0__inst_mult_6_67 ;
wire Xd_0__inst_mult_7_74 ;
wire Xd_0__inst_mult_7_75 ;
wire Xd_0__inst_mult_7_76 ;
wire Xd_0__inst_mult_4_65 ;
wire Xd_0__inst_mult_4_66 ;
wire Xd_0__inst_mult_4_67 ;
wire Xd_0__inst_mult_5_74 ;
wire Xd_0__inst_mult_5_75 ;
wire Xd_0__inst_mult_5_76 ;
wire Xd_0__inst_mult_2_74 ;
wire Xd_0__inst_mult_2_75 ;
wire Xd_0__inst_mult_2_76 ;
wire Xd_0__inst_mult_3_74 ;
wire Xd_0__inst_mult_3_75 ;
wire Xd_0__inst_mult_3_76 ;
wire Xd_0__inst_mult_0_74 ;
wire Xd_0__inst_mult_0_75 ;
wire Xd_0__inst_mult_0_76 ;
wire Xd_0__inst_mult_1_74 ;
wire Xd_0__inst_mult_1_75 ;
wire Xd_0__inst_mult_1_76 ;
wire Xd_0__inst_mult_28_87 ;
wire Xd_0__inst_mult_28_88 ;
wire Xd_0__inst_mult_28_89 ;
wire Xd_0__inst_mult_29_83 ;
wire Xd_0__inst_mult_29_84 ;
wire Xd_0__inst_mult_29_85 ;
wire Xd_0__inst_mult_26_87 ;
wire Xd_0__inst_mult_26_88 ;
wire Xd_0__inst_mult_26_89 ;
wire Xd_0__inst_mult_27_83 ;
wire Xd_0__inst_mult_27_84 ;
wire Xd_0__inst_mult_27_85 ;
wire Xd_0__inst_mult_24_87 ;
wire Xd_0__inst_mult_24_88 ;
wire Xd_0__inst_mult_24_89 ;
wire Xd_0__inst_mult_25_83 ;
wire Xd_0__inst_mult_25_84 ;
wire Xd_0__inst_mult_25_85 ;
wire Xd_0__inst_mult_22_87 ;
wire Xd_0__inst_mult_22_88 ;
wire Xd_0__inst_mult_22_89 ;
wire Xd_0__inst_mult_23_87 ;
wire Xd_0__inst_mult_23_88 ;
wire Xd_0__inst_mult_23_89 ;
wire Xd_0__inst_mult_20_87 ;
wire Xd_0__inst_mult_20_88 ;
wire Xd_0__inst_mult_20_89 ;
wire Xd_0__inst_mult_21_75 ;
wire Xd_0__inst_mult_21_76 ;
wire Xd_0__inst_mult_21_77 ;
wire Xd_0__inst_mult_18_66 ;
wire Xd_0__inst_mult_18_67 ;
wire Xd_0__inst_mult_18_68 ;
wire Xd_0__inst_mult_19_87 ;
wire Xd_0__inst_mult_19_88 ;
wire Xd_0__inst_mult_19_89 ;
wire Xd_0__inst_mult_16_71 ;
wire Xd_0__inst_mult_16_72 ;
wire Xd_0__inst_mult_17_80 ;
wire Xd_0__inst_mult_17_81 ;
wire Xd_0__inst_mult_14_71 ;
wire Xd_0__inst_mult_14_72 ;
wire Xd_0__inst_mult_15_80 ;
wire Xd_0__inst_mult_15_81 ;
wire Xd_0__inst_mult_12_71 ;
wire Xd_0__inst_mult_12_72 ;
wire Xd_0__inst_mult_13_80 ;
wire Xd_0__inst_mult_13_81 ;
wire Xd_0__inst_mult_10_71 ;
wire Xd_0__inst_mult_10_72 ;
wire Xd_0__inst_mult_11_88 ;
wire Xd_0__inst_mult_11_89 ;
wire Xd_0__inst_mult_8_71 ;
wire Xd_0__inst_mult_8_72 ;
wire Xd_0__inst_mult_9_80 ;
wire Xd_0__inst_mult_9_81 ;
wire Xd_0__inst_mult_6_70 ;
wire Xd_0__inst_mult_6_71 ;
wire Xd_0__inst_mult_7_79 ;
wire Xd_0__inst_mult_7_80 ;
wire Xd_0__inst_mult_4_70 ;
wire Xd_0__inst_mult_4_71 ;
wire Xd_0__inst_mult_5_79 ;
wire Xd_0__inst_mult_5_80 ;
wire Xd_0__inst_mult_2_79 ;
wire Xd_0__inst_mult_2_80 ;
wire Xd_0__inst_mult_3_79 ;
wire Xd_0__inst_mult_3_80 ;
wire Xd_0__inst_mult_0_79 ;
wire Xd_0__inst_mult_0_80 ;
wire Xd_0__inst_mult_1_79 ;
wire Xd_0__inst_mult_1_80 ;
wire Xd_0__inst_mult_28_92 ;
wire Xd_0__inst_mult_28_93 ;
wire Xd_0__inst_mult_29_88 ;
wire Xd_0__inst_mult_29_89 ;
wire Xd_0__inst_mult_26_92 ;
wire Xd_0__inst_mult_26_93 ;
wire Xd_0__inst_mult_27_88 ;
wire Xd_0__inst_mult_27_89 ;
wire Xd_0__inst_mult_24_92 ;
wire Xd_0__inst_mult_24_93 ;
wire Xd_0__inst_mult_25_88 ;
wire Xd_0__inst_mult_25_89 ;
wire Xd_0__inst_mult_22_92 ;
wire Xd_0__inst_mult_22_93 ;
wire Xd_0__inst_mult_23_92 ;
wire Xd_0__inst_mult_23_93 ;
wire Xd_0__inst_mult_20_92 ;
wire Xd_0__inst_mult_20_93 ;
wire Xd_0__inst_mult_21_80 ;
wire Xd_0__inst_mult_21_81 ;
wire Xd_0__inst_mult_18_71 ;
wire Xd_0__inst_mult_18_72 ;
wire Xd_0__inst_mult_19_92 ;
wire Xd_0__inst_mult_19_93 ;
wire Xd_0__inst_mult_30_99 ;
wire Xd_0__inst_mult_30_100 ;
wire Xd_0__inst_mult_30_101 ;
wire Xd_0__inst_mult_31_91 ;
wire Xd_0__inst_mult_31_92 ;
wire Xd_0__inst_mult_31_93 ;
wire Xd_0__inst_mult_30_103 ;
wire Xd_0__inst_mult_30_104 ;
wire Xd_0__inst_mult_30_105 ;
wire Xd_0__inst_mult_31_95 ;
wire Xd_0__inst_mult_31_96 ;
wire Xd_0__inst_mult_31_97 ;
wire Xd_0__inst_mult_30_107 ;
wire Xd_0__inst_mult_30_108 ;
wire Xd_0__inst_mult_30_109 ;
wire Xd_0__inst_mult_31_99 ;
wire Xd_0__inst_mult_31_100 ;
wire Xd_0__inst_mult_31_101 ;
wire Xd_0__inst_mult_30_111 ;
wire Xd_0__inst_mult_30_112 ;
wire Xd_0__inst_mult_30_113 ;
wire Xd_0__inst_mult_31_103 ;
wire Xd_0__inst_mult_31_104 ;
wire Xd_0__inst_mult_31_105 ;
wire Xd_0__inst_mult_30_115 ;
wire Xd_0__inst_mult_30_116 ;
wire Xd_0__inst_mult_30_117 ;
wire Xd_0__inst_mult_31_107 ;
wire Xd_0__inst_mult_31_108 ;
wire Xd_0__inst_mult_31_109 ;
wire Xd_0__inst_mult_31_111 ;
wire Xd_0__inst_mult_22_95 ;
wire Xd_0__inst_mult_22_96 ;
wire Xd_0__inst_mult_22_97 ;
wire Xd_0__inst_mult_15_83 ;
wire Xd_0__inst_mult_15_84 ;
wire Xd_0__inst_mult_15_85 ;
wire Xd_0__inst_mult_29_91 ;
wire Xd_0__inst_mult_29_92 ;
wire Xd_0__inst_mult_29_93 ;
wire Xd_0__inst_mult_29_96 ;
wire Xd_0__inst_mult_29_97 ;
wire Xd_0__inst_mult_11_91 ;
wire Xd_0__inst_mult_11_92 ;
wire Xd_0__inst_mult_11_93 ;
wire Xd_0__inst_mult_9_83 ;
wire Xd_0__inst_mult_9_84 ;
wire Xd_0__inst_mult_9_85 ;
wire Xd_0__inst_mult_31_116 ;
wire Xd_0__inst_mult_31_117 ;
wire Xd_0__inst_mult_8_74 ;
wire Xd_0__inst_mult_8_75 ;
wire Xd_0__inst_mult_8_76 ;
wire Xd_0__inst_mult_7_82 ;
wire Xd_0__inst_mult_7_83 ;
wire Xd_0__inst_mult_7_84 ;
wire Xd_0__inst_mult_2_82 ;
wire Xd_0__inst_mult_2_83 ;
wire Xd_0__inst_mult_2_84 ;
wire Xd_0__inst_mult_0_82 ;
wire Xd_0__inst_mult_0_83 ;
wire Xd_0__inst_mult_0_84 ;
wire Xd_0__inst_mult_11_96 ;
wire Xd_0__inst_mult_11_97 ;
wire Xd_0__inst_mult_21_83 ;
wire Xd_0__inst_mult_21_84 ;
wire Xd_0__inst_mult_21_85 ;
wire Xd_0__inst_mult_26_95 ;
wire Xd_0__inst_mult_26_96 ;
wire Xd_0__inst_mult_26_97 ;
wire Xd_0__inst_mult_24_95 ;
wire Xd_0__inst_mult_24_96 ;
wire Xd_0__inst_mult_24_97 ;
wire Xd_0__inst_mult_25_92 ;
wire Xd_0__inst_mult_25_93 ;
wire Xd_0__inst_mult_19_95 ;
wire Xd_0__inst_mult_19_96 ;
wire Xd_0__inst_mult_19_97 ;
wire Xd_0__inst_mult_17_83 ;
wire Xd_0__inst_mult_17_84 ;
wire Xd_0__inst_mult_17_85 ;
wire Xd_0__inst_mult_12_74 ;
wire Xd_0__inst_mult_12_75 ;
wire Xd_0__inst_mult_12_76 ;
wire Xd_0__inst_mult_27_92 ;
wire Xd_0__inst_mult_27_93 ;
wire Xd_0__inst_mult_16_74 ;
wire Xd_0__inst_mult_16_75 ;
wire Xd_0__inst_mult_16_76 ;
wire Xd_0__inst_mult_16_78 ;
wire Xd_0__inst_mult_16_79 ;
wire Xd_0__inst_mult_16_80 ;
wire Xd_0__inst_mult_17_87 ;
wire Xd_0__inst_mult_17_88 ;
wire Xd_0__inst_mult_17_89 ;
wire Xd_0__inst_mult_14_74 ;
wire Xd_0__inst_mult_14_75 ;
wire Xd_0__inst_mult_14_76 ;
wire Xd_0__inst_mult_14_78 ;
wire Xd_0__inst_mult_14_79 ;
wire Xd_0__inst_mult_14_80 ;
wire Xd_0__inst_mult_15_87 ;
wire Xd_0__inst_mult_15_88 ;
wire Xd_0__inst_mult_15_89 ;
wire Xd_0__inst_mult_12_78 ;
wire Xd_0__inst_mult_12_79 ;
wire Xd_0__inst_mult_12_80 ;
wire Xd_0__inst_mult_12_82 ;
wire Xd_0__inst_mult_12_83 ;
wire Xd_0__inst_mult_12_84 ;
wire Xd_0__inst_mult_13_83 ;
wire Xd_0__inst_mult_13_84 ;
wire Xd_0__inst_mult_13_85 ;
wire Xd_0__inst_mult_10_74 ;
wire Xd_0__inst_mult_10_75 ;
wire Xd_0__inst_mult_10_76 ;
wire Xd_0__inst_mult_10_78 ;
wire Xd_0__inst_mult_10_79 ;
wire Xd_0__inst_mult_10_80 ;
wire Xd_0__inst_mult_11_99 ;
wire Xd_0__inst_mult_11_100 ;
wire Xd_0__inst_mult_11_101 ;
wire Xd_0__inst_mult_8_78 ;
wire Xd_0__inst_mult_8_79 ;
wire Xd_0__inst_mult_8_80 ;
wire Xd_0__inst_mult_8_82 ;
wire Xd_0__inst_mult_8_83 ;
wire Xd_0__inst_mult_8_84 ;
wire Xd_0__inst_mult_9_87 ;
wire Xd_0__inst_mult_9_88 ;
wire Xd_0__inst_mult_9_89 ;
wire Xd_0__inst_mult_6_73 ;
wire Xd_0__inst_mult_6_74 ;
wire Xd_0__inst_mult_6_75 ;
wire Xd_0__inst_mult_6_77 ;
wire Xd_0__inst_mult_6_78 ;
wire Xd_0__inst_mult_6_79 ;
wire Xd_0__inst_mult_7_86 ;
wire Xd_0__inst_mult_7_87 ;
wire Xd_0__inst_mult_7_88 ;
wire Xd_0__inst_mult_4_73 ;
wire Xd_0__inst_mult_4_74 ;
wire Xd_0__inst_mult_4_75 ;
wire Xd_0__inst_mult_4_77 ;
wire Xd_0__inst_mult_4_78 ;
wire Xd_0__inst_mult_4_79 ;
wire Xd_0__inst_mult_5_82 ;
wire Xd_0__inst_mult_5_83 ;
wire Xd_0__inst_mult_5_84 ;
wire Xd_0__inst_mult_2_86 ;
wire Xd_0__inst_mult_2_87 ;
wire Xd_0__inst_mult_2_88 ;
wire Xd_0__inst_mult_3_82 ;
wire Xd_0__inst_mult_3_83 ;
wire Xd_0__inst_mult_3_84 ;
wire Xd_0__inst_mult_0_86 ;
wire Xd_0__inst_mult_0_87 ;
wire Xd_0__inst_mult_0_88 ;
wire Xd_0__inst_mult_1_82 ;
wire Xd_0__inst_mult_1_83 ;
wire Xd_0__inst_mult_1_84 ;
wire Xd_0__inst_mult_28_95 ;
wire Xd_0__inst_mult_28_96 ;
wire Xd_0__inst_mult_28_97 ;
wire Xd_0__inst_mult_29_99 ;
wire Xd_0__inst_mult_29_100 ;
wire Xd_0__inst_mult_29_101 ;
wire Xd_0__inst_mult_26_99 ;
wire Xd_0__inst_mult_26_100 ;
wire Xd_0__inst_mult_26_101 ;
wire Xd_0__inst_mult_27_95 ;
wire Xd_0__inst_mult_27_96 ;
wire Xd_0__inst_mult_27_97 ;
wire Xd_0__inst_mult_24_99 ;
wire Xd_0__inst_mult_24_100 ;
wire Xd_0__inst_mult_24_101 ;
wire Xd_0__inst_mult_25_95 ;
wire Xd_0__inst_mult_25_96 ;
wire Xd_0__inst_mult_25_97 ;
wire Xd_0__inst_mult_22_99 ;
wire Xd_0__inst_mult_22_100 ;
wire Xd_0__inst_mult_22_101 ;
wire Xd_0__inst_mult_23_95 ;
wire Xd_0__inst_mult_23_96 ;
wire Xd_0__inst_mult_23_97 ;
wire Xd_0__inst_mult_20_95 ;
wire Xd_0__inst_mult_20_96 ;
wire Xd_0__inst_mult_20_97 ;
wire Xd_0__inst_mult_21_87 ;
wire Xd_0__inst_mult_21_88 ;
wire Xd_0__inst_mult_21_89 ;
wire Xd_0__inst_mult_18_74 ;
wire Xd_0__inst_mult_18_75 ;
wire Xd_0__inst_mult_18_76 ;
wire Xd_0__inst_mult_18_78 ;
wire Xd_0__inst_mult_18_79 ;
wire Xd_0__inst_mult_18_80 ;
wire Xd_0__inst_mult_19_99 ;
wire Xd_0__inst_mult_19_100 ;
wire Xd_0__inst_mult_19_101 ;
wire Xd_0__inst_mult_16_82 ;
wire Xd_0__inst_mult_16_83 ;
wire Xd_0__inst_mult_16_84 ;
wire Xd_0__inst_mult_16_86 ;
wire Xd_0__inst_mult_16_87 ;
wire Xd_0__inst_mult_16_88 ;
wire Xd_0__inst_mult_17_91 ;
wire Xd_0__inst_mult_17_92 ;
wire Xd_0__inst_mult_17_93 ;
wire Xd_0__inst_mult_17_95 ;
wire Xd_0__inst_mult_17_96 ;
wire Xd_0__inst_mult_17_97 ;
wire Xd_0__inst_mult_14_82 ;
wire Xd_0__inst_mult_14_83 ;
wire Xd_0__inst_mult_14_84 ;
wire Xd_0__inst_mult_14_86 ;
wire Xd_0__inst_mult_14_87 ;
wire Xd_0__inst_mult_14_88 ;
wire Xd_0__inst_mult_15_91 ;
wire Xd_0__inst_mult_15_92 ;
wire Xd_0__inst_mult_15_93 ;
wire Xd_0__inst_mult_15_95 ;
wire Xd_0__inst_mult_15_96 ;
wire Xd_0__inst_mult_15_97 ;
wire Xd_0__inst_mult_12_86 ;
wire Xd_0__inst_mult_12_87 ;
wire Xd_0__inst_mult_12_88 ;
wire Xd_0__inst_mult_12_90 ;
wire Xd_0__inst_mult_12_91 ;
wire Xd_0__inst_mult_12_92 ;
wire Xd_0__inst_mult_13_87 ;
wire Xd_0__inst_mult_13_88 ;
wire Xd_0__inst_mult_13_89 ;
wire Xd_0__inst_mult_13_91 ;
wire Xd_0__inst_mult_13_92 ;
wire Xd_0__inst_mult_13_93 ;
wire Xd_0__inst_mult_10_82 ;
wire Xd_0__inst_mult_10_83 ;
wire Xd_0__inst_mult_10_84 ;
wire Xd_0__inst_mult_10_86 ;
wire Xd_0__inst_mult_10_87 ;
wire Xd_0__inst_mult_10_88 ;
wire Xd_0__inst_mult_11_103 ;
wire Xd_0__inst_mult_11_104 ;
wire Xd_0__inst_mult_11_105 ;
wire Xd_0__inst_mult_8_86 ;
wire Xd_0__inst_mult_8_87 ;
wire Xd_0__inst_mult_8_88 ;
wire Xd_0__inst_mult_8_90 ;
wire Xd_0__inst_mult_8_91 ;
wire Xd_0__inst_mult_8_92 ;
wire Xd_0__inst_mult_9_91 ;
wire Xd_0__inst_mult_9_92 ;
wire Xd_0__inst_mult_9_93 ;
wire Xd_0__inst_mult_9_95 ;
wire Xd_0__inst_mult_9_96 ;
wire Xd_0__inst_mult_9_97 ;
wire Xd_0__inst_mult_6_81 ;
wire Xd_0__inst_mult_6_82 ;
wire Xd_0__inst_mult_6_83 ;
wire Xd_0__inst_mult_6_85 ;
wire Xd_0__inst_mult_6_86 ;
wire Xd_0__inst_mult_6_87 ;
wire Xd_0__inst_mult_7_90 ;
wire Xd_0__inst_mult_7_91 ;
wire Xd_0__inst_mult_7_92 ;
wire Xd_0__inst_mult_7_94 ;
wire Xd_0__inst_mult_7_95 ;
wire Xd_0__inst_mult_7_96 ;
wire Xd_0__inst_mult_4_81 ;
wire Xd_0__inst_mult_4_82 ;
wire Xd_0__inst_mult_4_83 ;
wire Xd_0__inst_mult_4_85 ;
wire Xd_0__inst_mult_4_86 ;
wire Xd_0__inst_mult_4_87 ;
wire Xd_0__inst_mult_5_86 ;
wire Xd_0__inst_mult_5_87 ;
wire Xd_0__inst_mult_5_88 ;
wire Xd_0__inst_mult_5_90 ;
wire Xd_0__inst_mult_5_91 ;
wire Xd_0__inst_mult_5_92 ;
wire Xd_0__inst_mult_2_90 ;
wire Xd_0__inst_mult_2_91 ;
wire Xd_0__inst_mult_2_92 ;
wire Xd_0__inst_mult_2_94 ;
wire Xd_0__inst_mult_2_95 ;
wire Xd_0__inst_mult_2_96 ;
wire Xd_0__inst_mult_3_86 ;
wire Xd_0__inst_mult_3_87 ;
wire Xd_0__inst_mult_3_88 ;
wire Xd_0__inst_mult_3_90 ;
wire Xd_0__inst_mult_3_91 ;
wire Xd_0__inst_mult_3_92 ;
wire Xd_0__inst_mult_0_90 ;
wire Xd_0__inst_mult_0_91 ;
wire Xd_0__inst_mult_0_92 ;
wire Xd_0__inst_mult_0_94 ;
wire Xd_0__inst_mult_0_95 ;
wire Xd_0__inst_mult_0_96 ;
wire Xd_0__inst_mult_1_86 ;
wire Xd_0__inst_mult_1_87 ;
wire Xd_0__inst_mult_1_88 ;
wire Xd_0__inst_mult_1_90 ;
wire Xd_0__inst_mult_1_91 ;
wire Xd_0__inst_mult_1_92 ;
wire Xd_0__inst_mult_28_99 ;
wire Xd_0__inst_mult_28_100 ;
wire Xd_0__inst_mult_28_101 ;
wire Xd_0__inst_mult_29_103 ;
wire Xd_0__inst_mult_29_104 ;
wire Xd_0__inst_mult_29_105 ;
wire Xd_0__inst_mult_26_103 ;
wire Xd_0__inst_mult_26_104 ;
wire Xd_0__inst_mult_26_105 ;
wire Xd_0__inst_mult_27_99 ;
wire Xd_0__inst_mult_27_100 ;
wire Xd_0__inst_mult_27_101 ;
wire Xd_0__inst_mult_24_103 ;
wire Xd_0__inst_mult_24_104 ;
wire Xd_0__inst_mult_24_105 ;
wire Xd_0__inst_mult_25_99 ;
wire Xd_0__inst_mult_25_100 ;
wire Xd_0__inst_mult_25_101 ;
wire Xd_0__inst_mult_22_103 ;
wire Xd_0__inst_mult_22_104 ;
wire Xd_0__inst_mult_22_105 ;
wire Xd_0__inst_mult_23_99 ;
wire Xd_0__inst_mult_23_100 ;
wire Xd_0__inst_mult_23_101 ;
wire Xd_0__inst_mult_20_99 ;
wire Xd_0__inst_mult_20_100 ;
wire Xd_0__inst_mult_20_101 ;
wire Xd_0__inst_mult_21_91 ;
wire Xd_0__inst_mult_21_92 ;
wire Xd_0__inst_mult_21_93 ;
wire Xd_0__inst_mult_21_95 ;
wire Xd_0__inst_mult_21_96 ;
wire Xd_0__inst_mult_21_97 ;
wire Xd_0__inst_mult_18_82 ;
wire Xd_0__inst_mult_18_83 ;
wire Xd_0__inst_mult_18_84 ;
wire Xd_0__inst_mult_18_86 ;
wire Xd_0__inst_mult_18_87 ;
wire Xd_0__inst_mult_18_88 ;
wire Xd_0__inst_mult_19_103 ;
wire Xd_0__inst_mult_19_104 ;
wire Xd_0__inst_mult_19_105 ;
wire Xd_0__inst_mult_16_90 ;
wire Xd_0__inst_mult_16_91 ;
wire Xd_0__inst_mult_16_92 ;
wire Xd_0__inst_mult_16_94 ;
wire Xd_0__inst_mult_16_95 ;
wire Xd_0__inst_mult_16_96 ;
wire Xd_0__inst_mult_17_99 ;
wire Xd_0__inst_mult_17_100 ;
wire Xd_0__inst_mult_17_101 ;
wire Xd_0__inst_mult_17_103 ;
wire Xd_0__inst_mult_17_104 ;
wire Xd_0__inst_mult_17_105 ;
wire Xd_0__inst_mult_14_90 ;
wire Xd_0__inst_mult_14_91 ;
wire Xd_0__inst_mult_14_92 ;
wire Xd_0__inst_mult_14_94 ;
wire Xd_0__inst_mult_14_95 ;
wire Xd_0__inst_mult_14_96 ;
wire Xd_0__inst_mult_15_99 ;
wire Xd_0__inst_mult_15_100 ;
wire Xd_0__inst_mult_15_101 ;
wire Xd_0__inst_mult_15_103 ;
wire Xd_0__inst_mult_12_94 ;
wire Xd_0__inst_mult_12_95 ;
wire Xd_0__inst_mult_12_96 ;
wire Xd_0__inst_mult_12_98 ;
wire Xd_0__inst_mult_12_99 ;
wire Xd_0__inst_mult_12_100 ;
wire Xd_0__inst_mult_13_95 ;
wire Xd_0__inst_mult_13_96 ;
wire Xd_0__inst_mult_13_97 ;
wire Xd_0__inst_mult_13_99 ;
wire Xd_0__inst_mult_13_100 ;
wire Xd_0__inst_mult_13_101 ;
wire Xd_0__inst_mult_10_90 ;
wire Xd_0__inst_mult_10_91 ;
wire Xd_0__inst_mult_10_92 ;
wire Xd_0__inst_mult_10_94 ;
wire Xd_0__inst_mult_10_95 ;
wire Xd_0__inst_mult_10_96 ;
wire Xd_0__inst_mult_11_107 ;
wire Xd_0__inst_mult_11_108 ;
wire Xd_0__inst_mult_11_109 ;
wire Xd_0__inst_mult_8_94 ;
wire Xd_0__inst_mult_8_95 ;
wire Xd_0__inst_mult_8_96 ;
wire Xd_0__inst_mult_8_98 ;
wire Xd_0__inst_mult_8_99 ;
wire Xd_0__inst_mult_8_100 ;
wire Xd_0__inst_mult_9_99 ;
wire Xd_0__inst_mult_9_100 ;
wire Xd_0__inst_mult_9_101 ;
wire Xd_0__inst_mult_9_103 ;
wire Xd_0__inst_mult_6_89 ;
wire Xd_0__inst_mult_6_90 ;
wire Xd_0__inst_mult_6_91 ;
wire Xd_0__inst_mult_7_98 ;
wire Xd_0__inst_mult_7_99 ;
wire Xd_0__inst_mult_7_100 ;
wire Xd_0__inst_mult_4_89 ;
wire Xd_0__inst_mult_4_90 ;
wire Xd_0__inst_mult_4_91 ;
wire Xd_0__inst_mult_5_94 ;
wire Xd_0__inst_mult_5_95 ;
wire Xd_0__inst_mult_5_96 ;
wire Xd_0__inst_mult_2_98 ;
wire Xd_0__inst_mult_2_99 ;
wire Xd_0__inst_mult_2_100 ;
wire Xd_0__inst_mult_3_94 ;
wire Xd_0__inst_mult_3_95 ;
wire Xd_0__inst_mult_3_96 ;
wire Xd_0__inst_mult_0_98 ;
wire Xd_0__inst_mult_0_99 ;
wire Xd_0__inst_mult_0_100 ;
wire Xd_0__inst_mult_1_94 ;
wire Xd_0__inst_mult_1_95 ;
wire Xd_0__inst_mult_1_96 ;
wire Xd_0__inst_mult_28_103 ;
wire Xd_0__inst_mult_28_104 ;
wire Xd_0__inst_mult_28_105 ;
wire Xd_0__inst_mult_29_107 ;
wire Xd_0__inst_mult_29_108 ;
wire Xd_0__inst_mult_29_109 ;
wire Xd_0__inst_mult_26_107 ;
wire Xd_0__inst_mult_26_108 ;
wire Xd_0__inst_mult_26_109 ;
wire Xd_0__inst_mult_27_103 ;
wire Xd_0__inst_mult_27_104 ;
wire Xd_0__inst_mult_27_105 ;
wire Xd_0__inst_mult_24_107 ;
wire Xd_0__inst_mult_24_108 ;
wire Xd_0__inst_mult_24_109 ;
wire Xd_0__inst_mult_25_103 ;
wire Xd_0__inst_mult_25_104 ;
wire Xd_0__inst_mult_25_105 ;
wire Xd_0__inst_mult_22_107 ;
wire Xd_0__inst_mult_22_108 ;
wire Xd_0__inst_mult_22_109 ;
wire Xd_0__inst_mult_23_103 ;
wire Xd_0__inst_mult_23_104 ;
wire Xd_0__inst_mult_23_105 ;
wire Xd_0__inst_mult_20_103 ;
wire Xd_0__inst_mult_20_104 ;
wire Xd_0__inst_mult_20_105 ;
wire Xd_0__inst_mult_21_99 ;
wire Xd_0__inst_mult_21_100 ;
wire Xd_0__inst_mult_21_101 ;
wire Xd_0__inst_mult_21_103 ;
wire Xd_0__inst_mult_21_104 ;
wire Xd_0__inst_mult_21_105 ;
wire Xd_0__inst_mult_18_90 ;
wire Xd_0__inst_mult_18_91 ;
wire Xd_0__inst_mult_18_92 ;
wire Xd_0__inst_mult_18_94 ;
wire Xd_0__inst_mult_18_95 ;
wire Xd_0__inst_mult_18_96 ;
wire Xd_0__inst_mult_19_107 ;
wire Xd_0__inst_mult_19_108 ;
wire Xd_0__inst_mult_19_109 ;
wire Xd_0__inst_mult_16_98 ;
wire Xd_0__inst_mult_16_99 ;
wire Xd_0__inst_mult_16_100 ;
wire Xd_0__inst_mult_17_107 ;
wire Xd_0__inst_mult_17_108 ;
wire Xd_0__inst_mult_17_109 ;
wire Xd_0__inst_mult_14_98 ;
wire Xd_0__inst_mult_14_99 ;
wire Xd_0__inst_mult_14_100 ;
wire Xd_0__inst_mult_15_107 ;
wire Xd_0__inst_mult_15_108 ;
wire Xd_0__inst_mult_15_109 ;
wire Xd_0__inst_mult_12_102 ;
wire Xd_0__inst_mult_12_103 ;
wire Xd_0__inst_mult_12_104 ;
wire Xd_0__inst_mult_13_103 ;
wire Xd_0__inst_mult_13_104 ;
wire Xd_0__inst_mult_13_105 ;
wire Xd_0__inst_mult_10_98 ;
wire Xd_0__inst_mult_10_99 ;
wire Xd_0__inst_mult_10_100 ;
wire Xd_0__inst_mult_11_111 ;
wire Xd_0__inst_mult_11_112 ;
wire Xd_0__inst_mult_11_113 ;
wire Xd_0__inst_mult_8_102 ;
wire Xd_0__inst_mult_8_103 ;
wire Xd_0__inst_mult_8_104 ;
wire Xd_0__inst_mult_9_107 ;
wire Xd_0__inst_mult_9_108 ;
wire Xd_0__inst_mult_9_109 ;
wire Xd_0__inst_mult_6_93 ;
wire Xd_0__inst_mult_6_94 ;
wire Xd_0__inst_mult_6_95 ;
wire Xd_0__inst_mult_7_102 ;
wire Xd_0__inst_mult_7_103 ;
wire Xd_0__inst_mult_7_104 ;
wire Xd_0__inst_mult_4_93 ;
wire Xd_0__inst_mult_4_94 ;
wire Xd_0__inst_mult_4_95 ;
wire Xd_0__inst_mult_5_98 ;
wire Xd_0__inst_mult_5_99 ;
wire Xd_0__inst_mult_5_100 ;
wire Xd_0__inst_mult_2_102 ;
wire Xd_0__inst_mult_2_103 ;
wire Xd_0__inst_mult_2_104 ;
wire Xd_0__inst_mult_3_98 ;
wire Xd_0__inst_mult_3_99 ;
wire Xd_0__inst_mult_3_100 ;
wire Xd_0__inst_mult_0_102 ;
wire Xd_0__inst_mult_0_103 ;
wire Xd_0__inst_mult_0_104 ;
wire Xd_0__inst_mult_1_98 ;
wire Xd_0__inst_mult_1_99 ;
wire Xd_0__inst_mult_1_100 ;
wire Xd_0__inst_mult_28_107 ;
wire Xd_0__inst_mult_28_108 ;
wire Xd_0__inst_mult_28_109 ;
wire Xd_0__inst_mult_29_111 ;
wire Xd_0__inst_mult_29_112 ;
wire Xd_0__inst_mult_29_113 ;
wire Xd_0__inst_mult_26_111 ;
wire Xd_0__inst_mult_26_112 ;
wire Xd_0__inst_mult_26_113 ;
wire Xd_0__inst_mult_27_107 ;
wire Xd_0__inst_mult_27_108 ;
wire Xd_0__inst_mult_27_109 ;
wire Xd_0__inst_mult_24_111 ;
wire Xd_0__inst_mult_24_112 ;
wire Xd_0__inst_mult_24_113 ;
wire Xd_0__inst_mult_25_107 ;
wire Xd_0__inst_mult_25_108 ;
wire Xd_0__inst_mult_25_109 ;
wire Xd_0__inst_mult_22_111 ;
wire Xd_0__inst_mult_22_112 ;
wire Xd_0__inst_mult_22_113 ;
wire Xd_0__inst_mult_23_107 ;
wire Xd_0__inst_mult_23_108 ;
wire Xd_0__inst_mult_23_109 ;
wire Xd_0__inst_mult_20_107 ;
wire Xd_0__inst_mult_20_108 ;
wire Xd_0__inst_mult_20_109 ;
wire Xd_0__inst_mult_21_107 ;
wire Xd_0__inst_mult_21_108 ;
wire Xd_0__inst_mult_21_109 ;
wire Xd_0__inst_mult_18_98 ;
wire Xd_0__inst_mult_18_99 ;
wire Xd_0__inst_mult_18_100 ;
wire Xd_0__inst_mult_19_111 ;
wire Xd_0__inst_mult_19_112 ;
wire Xd_0__inst_mult_19_113 ;
wire Xd_0__inst_mult_16_102 ;
wire Xd_0__inst_mult_16_103 ;
wire Xd_0__inst_mult_16_104 ;
wire Xd_0__inst_mult_17_111 ;
wire Xd_0__inst_mult_17_112 ;
wire Xd_0__inst_mult_17_113 ;
wire Xd_0__inst_mult_14_102 ;
wire Xd_0__inst_mult_14_103 ;
wire Xd_0__inst_mult_14_104 ;
wire Xd_0__inst_mult_15_111 ;
wire Xd_0__inst_mult_15_112 ;
wire Xd_0__inst_mult_15_113 ;
wire Xd_0__inst_mult_12_106 ;
wire Xd_0__inst_mult_12_107 ;
wire Xd_0__inst_mult_12_108 ;
wire Xd_0__inst_mult_13_107 ;
wire Xd_0__inst_mult_13_108 ;
wire Xd_0__inst_mult_13_109 ;
wire Xd_0__inst_mult_10_102 ;
wire Xd_0__inst_mult_10_103 ;
wire Xd_0__inst_mult_10_104 ;
wire Xd_0__inst_mult_11_115 ;
wire Xd_0__inst_mult_11_116 ;
wire Xd_0__inst_mult_11_117 ;
wire Xd_0__inst_mult_8_106 ;
wire Xd_0__inst_mult_8_107 ;
wire Xd_0__inst_mult_8_108 ;
wire Xd_0__inst_mult_9_111 ;
wire Xd_0__inst_mult_9_112 ;
wire Xd_0__inst_mult_9_113 ;
wire Xd_0__inst_mult_6_97 ;
wire Xd_0__inst_mult_6_98 ;
wire Xd_0__inst_mult_6_99 ;
wire Xd_0__inst_mult_7_106 ;
wire Xd_0__inst_mult_7_107 ;
wire Xd_0__inst_mult_7_108 ;
wire Xd_0__inst_mult_4_97 ;
wire Xd_0__inst_mult_4_98 ;
wire Xd_0__inst_mult_4_99 ;
wire Xd_0__inst_mult_5_102 ;
wire Xd_0__inst_mult_5_103 ;
wire Xd_0__inst_mult_5_104 ;
wire Xd_0__inst_mult_2_106 ;
wire Xd_0__inst_mult_2_107 ;
wire Xd_0__inst_mult_2_108 ;
wire Xd_0__inst_mult_3_102 ;
wire Xd_0__inst_mult_3_103 ;
wire Xd_0__inst_mult_3_104 ;
wire Xd_0__inst_mult_0_106 ;
wire Xd_0__inst_mult_0_107 ;
wire Xd_0__inst_mult_0_108 ;
wire Xd_0__inst_mult_1_102 ;
wire Xd_0__inst_mult_1_103 ;
wire Xd_0__inst_mult_1_104 ;
wire Xd_0__inst_mult_28_111 ;
wire Xd_0__inst_mult_28_112 ;
wire Xd_0__inst_mult_28_113 ;
wire Xd_0__inst_mult_29_115 ;
wire Xd_0__inst_mult_29_116 ;
wire Xd_0__inst_mult_29_117 ;
wire Xd_0__inst_mult_26_115 ;
wire Xd_0__inst_mult_26_116 ;
wire Xd_0__inst_mult_26_117 ;
wire Xd_0__inst_mult_27_111 ;
wire Xd_0__inst_mult_27_112 ;
wire Xd_0__inst_mult_27_113 ;
wire Xd_0__inst_mult_24_115 ;
wire Xd_0__inst_mult_24_116 ;
wire Xd_0__inst_mult_24_117 ;
wire Xd_0__inst_mult_25_111 ;
wire Xd_0__inst_mult_25_112 ;
wire Xd_0__inst_mult_25_113 ;
wire Xd_0__inst_mult_22_115 ;
wire Xd_0__inst_mult_22_116 ;
wire Xd_0__inst_mult_22_117 ;
wire Xd_0__inst_mult_23_111 ;
wire Xd_0__inst_mult_23_112 ;
wire Xd_0__inst_mult_23_113 ;
wire Xd_0__inst_mult_20_111 ;
wire Xd_0__inst_mult_20_112 ;
wire Xd_0__inst_mult_20_113 ;
wire Xd_0__inst_mult_21_111 ;
wire Xd_0__inst_mult_21_112 ;
wire Xd_0__inst_mult_21_113 ;
wire Xd_0__inst_mult_18_102 ;
wire Xd_0__inst_mult_18_103 ;
wire Xd_0__inst_mult_18_104 ;
wire Xd_0__inst_mult_19_115 ;
wire Xd_0__inst_mult_19_116 ;
wire Xd_0__inst_mult_19_117 ;
wire Xd_0__inst_mult_16_106 ;
wire Xd_0__inst_mult_14_106 ;
wire Xd_0__inst_mult_13_111 ;
wire Xd_0__inst_mult_10_106 ;
wire Xd_0__inst_mult_6_101 ;
wire Xd_0__inst_mult_4_101 ;
wire Xd_0__inst_mult_5_106 ;
wire Xd_0__inst_mult_3_106 ;
wire Xd_0__inst_mult_1_106 ;
wire Xd_0__inst_mult_28_115 ;
wire Xd_0__inst_mult_27_115 ;
wire Xd_0__inst_mult_25_115 ;
wire Xd_0__inst_mult_23_115 ;
wire Xd_0__inst_mult_20_115 ;
wire Xd_0__inst_mult_18_106 ;
wire Xd_0__inst_mult_16_111 ;
wire Xd_0__inst_mult_16_112 ;
wire Xd_0__inst_mult_17_116 ;
wire Xd_0__inst_mult_17_117 ;
wire Xd_0__inst_mult_14_111 ;
wire Xd_0__inst_mult_14_112 ;
wire Xd_0__inst_mult_15_116 ;
wire Xd_0__inst_mult_15_117 ;
wire Xd_0__inst_mult_12_111 ;
wire Xd_0__inst_mult_12_112 ;
wire Xd_0__inst_mult_13_116 ;
wire Xd_0__inst_mult_13_117 ;
wire Xd_0__inst_mult_10_111 ;
wire Xd_0__inst_mult_10_112 ;
wire Xd_0__inst_mult_8_111 ;
wire Xd_0__inst_mult_8_112 ;
wire Xd_0__inst_mult_9_116 ;
wire Xd_0__inst_mult_9_117 ;
wire Xd_0__inst_mult_6_106 ;
wire Xd_0__inst_mult_6_107 ;
wire Xd_0__inst_mult_7_111 ;
wire Xd_0__inst_mult_7_112 ;
wire Xd_0__inst_mult_4_106 ;
wire Xd_0__inst_mult_4_107 ;
wire Xd_0__inst_mult_5_111 ;
wire Xd_0__inst_mult_5_112 ;
wire Xd_0__inst_mult_2_111 ;
wire Xd_0__inst_mult_2_112 ;
wire Xd_0__inst_mult_3_111 ;
wire Xd_0__inst_mult_3_112 ;
wire Xd_0__inst_mult_0_111 ;
wire Xd_0__inst_mult_0_112 ;
wire Xd_0__inst_mult_1_111 ;
wire Xd_0__inst_mult_1_112 ;
wire Xd_0__inst_mult_21_116 ;
wire Xd_0__inst_mult_21_117 ;
wire Xd_0__inst_mult_18_111 ;
wire Xd_0__inst_mult_18_112 ;
wire Xd_0__inst_inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_2__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_4__0__q ;
wire Xd_0__inst_inst_first_level_3__0__q ;
wire Xd_0__inst_inst_first_level_5__0__q ;
wire Xd_0__inst_inst_first_level_2__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_4__1__q ;
wire Xd_0__inst_inst_first_level_3__1__q ;
wire Xd_0__inst_inst_first_level_5__1__q ;
wire Xd_0__inst_inst_first_level_2__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_4__2__q ;
wire Xd_0__inst_inst_first_level_3__2__q ;
wire Xd_0__inst_inst_first_level_5__2__q ;
wire Xd_0__inst_inst_first_level_2__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_4__3__q ;
wire Xd_0__inst_inst_first_level_3__3__q ;
wire Xd_0__inst_inst_first_level_5__3__q ;
wire Xd_0__inst_inst_first_level_2__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_4__4__q ;
wire Xd_0__inst_inst_first_level_3__4__q ;
wire Xd_0__inst_inst_first_level_5__4__q ;
wire Xd_0__inst_inst_first_level_2__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_4__5__q ;
wire Xd_0__inst_inst_first_level_3__5__q ;
wire Xd_0__inst_inst_first_level_5__5__q ;
wire Xd_0__inst_inst_first_level_2__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_4__6__q ;
wire Xd_0__inst_inst_first_level_3__6__q ;
wire Xd_0__inst_inst_first_level_5__6__q ;
wire Xd_0__inst_inst_first_level_2__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_4__7__q ;
wire Xd_0__inst_inst_first_level_3__7__q ;
wire Xd_0__inst_inst_first_level_5__7__q ;
wire Xd_0__inst_inst_first_level_2__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_4__8__q ;
wire Xd_0__inst_inst_first_level_3__8__q ;
wire Xd_0__inst_inst_first_level_5__8__q ;
wire Xd_0__inst_inst_first_level_2__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_4__9__q ;
wire Xd_0__inst_inst_first_level_3__9__q ;
wire Xd_0__inst_inst_first_level_5__9__q ;
wire Xd_0__inst_inst_first_level_2__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_4__10__q ;
wire Xd_0__inst_inst_first_level_3__10__q ;
wire Xd_0__inst_inst_first_level_5__10__q ;
wire Xd_0__inst_inst_first_level_2__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_4__11__q ;
wire Xd_0__inst_inst_first_level_3__11__q ;
wire Xd_0__inst_inst_first_level_5__13__q ;
wire Xd_0__inst_inst_first_level_2__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_4__12__q ;
wire Xd_0__inst_inst_first_level_3__12__q ;
wire Xd_0__inst_inst_first_level_2__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_4__13__q ;
wire Xd_0__inst_inst_first_level_3__13__q ;
wire Xd_0__inst_r_sum1_15__0__q ;
wire Xd_0__inst_r_sum1_15__1__q ;
wire Xd_0__inst_r_sum1_15__2__q ;
wire Xd_0__inst_r_sum1_15__3__q ;
wire Xd_0__inst_r_sum1_15__4__q ;
wire Xd_0__inst_r_sum1_15__5__q ;
wire Xd_0__inst_r_sum1_15__6__q ;
wire Xd_0__inst_r_sum1_15__7__q ;
wire Xd_0__inst_r_sum1_15__8__q ;
wire Xd_0__inst_r_sum1_15__9__q ;
wire Xd_0__inst_r_sum1_15__10__q ;
wire Xd_0__inst_r_sum1_15__11__q ;
wire Xd_0__inst_r_sum1_8__0__q ;
wire Xd_0__inst_r_sum1_7__0__q ;
wire Xd_0__inst_r_sum1_6__0__q ;
wire Xd_0__inst_r_sum1_5__0__q ;
wire Xd_0__inst_r_sum1_4__0__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_14__0__q ;
wire Xd_0__inst_r_sum1_13__0__q ;
wire Xd_0__inst_r_sum1_12__0__q ;
wire Xd_0__inst_r_sum1_11__0__q ;
wire Xd_0__inst_r_sum1_10__0__q ;
wire Xd_0__inst_r_sum1_9__0__q ;
wire Xd_0__inst_r_sum1_8__1__q ;
wire Xd_0__inst_r_sum1_7__1__q ;
wire Xd_0__inst_r_sum1_6__1__q ;
wire Xd_0__inst_r_sum1_5__1__q ;
wire Xd_0__inst_r_sum1_4__1__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_14__1__q ;
wire Xd_0__inst_r_sum1_13__1__q ;
wire Xd_0__inst_r_sum1_12__1__q ;
wire Xd_0__inst_r_sum1_11__1__q ;
wire Xd_0__inst_r_sum1_10__1__q ;
wire Xd_0__inst_r_sum1_9__1__q ;
wire Xd_0__inst_r_sum1_8__2__q ;
wire Xd_0__inst_r_sum1_7__2__q ;
wire Xd_0__inst_r_sum1_6__2__q ;
wire Xd_0__inst_r_sum1_5__2__q ;
wire Xd_0__inst_r_sum1_4__2__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_14__2__q ;
wire Xd_0__inst_r_sum1_13__2__q ;
wire Xd_0__inst_r_sum1_12__2__q ;
wire Xd_0__inst_r_sum1_11__2__q ;
wire Xd_0__inst_r_sum1_10__2__q ;
wire Xd_0__inst_r_sum1_9__2__q ;
wire Xd_0__inst_r_sum1_8__3__q ;
wire Xd_0__inst_r_sum1_7__3__q ;
wire Xd_0__inst_r_sum1_6__3__q ;
wire Xd_0__inst_r_sum1_5__3__q ;
wire Xd_0__inst_r_sum1_4__3__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_14__3__q ;
wire Xd_0__inst_r_sum1_13__3__q ;
wire Xd_0__inst_r_sum1_12__3__q ;
wire Xd_0__inst_r_sum1_11__3__q ;
wire Xd_0__inst_r_sum1_10__3__q ;
wire Xd_0__inst_r_sum1_9__3__q ;
wire Xd_0__inst_r_sum1_8__4__q ;
wire Xd_0__inst_r_sum1_7__4__q ;
wire Xd_0__inst_r_sum1_6__4__q ;
wire Xd_0__inst_r_sum1_5__4__q ;
wire Xd_0__inst_r_sum1_4__4__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_14__4__q ;
wire Xd_0__inst_r_sum1_13__4__q ;
wire Xd_0__inst_r_sum1_12__4__q ;
wire Xd_0__inst_r_sum1_11__4__q ;
wire Xd_0__inst_r_sum1_10__4__q ;
wire Xd_0__inst_r_sum1_9__4__q ;
wire Xd_0__inst_r_sum1_8__5__q ;
wire Xd_0__inst_r_sum1_7__5__q ;
wire Xd_0__inst_r_sum1_6__5__q ;
wire Xd_0__inst_r_sum1_5__5__q ;
wire Xd_0__inst_r_sum1_4__5__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_14__5__q ;
wire Xd_0__inst_r_sum1_13__5__q ;
wire Xd_0__inst_r_sum1_12__5__q ;
wire Xd_0__inst_r_sum1_11__5__q ;
wire Xd_0__inst_r_sum1_10__5__q ;
wire Xd_0__inst_r_sum1_9__5__q ;
wire Xd_0__inst_r_sum1_8__6__q ;
wire Xd_0__inst_r_sum1_7__6__q ;
wire Xd_0__inst_r_sum1_6__6__q ;
wire Xd_0__inst_r_sum1_5__6__q ;
wire Xd_0__inst_r_sum1_4__6__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_14__6__q ;
wire Xd_0__inst_r_sum1_13__6__q ;
wire Xd_0__inst_r_sum1_12__6__q ;
wire Xd_0__inst_r_sum1_11__6__q ;
wire Xd_0__inst_r_sum1_10__6__q ;
wire Xd_0__inst_r_sum1_9__6__q ;
wire Xd_0__inst_r_sum1_8__7__q ;
wire Xd_0__inst_r_sum1_7__7__q ;
wire Xd_0__inst_r_sum1_6__7__q ;
wire Xd_0__inst_r_sum1_5__7__q ;
wire Xd_0__inst_r_sum1_4__7__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_14__7__q ;
wire Xd_0__inst_r_sum1_13__7__q ;
wire Xd_0__inst_r_sum1_12__7__q ;
wire Xd_0__inst_r_sum1_11__7__q ;
wire Xd_0__inst_r_sum1_10__7__q ;
wire Xd_0__inst_r_sum1_9__7__q ;
wire Xd_0__inst_r_sum1_8__8__q ;
wire Xd_0__inst_r_sum1_7__8__q ;
wire Xd_0__inst_r_sum1_6__8__q ;
wire Xd_0__inst_r_sum1_5__8__q ;
wire Xd_0__inst_r_sum1_4__8__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_14__8__q ;
wire Xd_0__inst_r_sum1_13__8__q ;
wire Xd_0__inst_r_sum1_12__8__q ;
wire Xd_0__inst_r_sum1_11__8__q ;
wire Xd_0__inst_r_sum1_10__8__q ;
wire Xd_0__inst_r_sum1_9__8__q ;
wire Xd_0__inst_r_sum1_8__9__q ;
wire Xd_0__inst_r_sum1_7__9__q ;
wire Xd_0__inst_r_sum1_6__9__q ;
wire Xd_0__inst_r_sum1_5__9__q ;
wire Xd_0__inst_r_sum1_4__9__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_14__9__q ;
wire Xd_0__inst_r_sum1_13__9__q ;
wire Xd_0__inst_r_sum1_12__9__q ;
wire Xd_0__inst_r_sum1_11__9__q ;
wire Xd_0__inst_r_sum1_10__9__q ;
wire Xd_0__inst_r_sum1_9__9__q ;
wire Xd_0__inst_r_sum1_8__10__q ;
wire Xd_0__inst_r_sum1_7__10__q ;
wire Xd_0__inst_r_sum1_6__10__q ;
wire Xd_0__inst_r_sum1_5__10__q ;
wire Xd_0__inst_r_sum1_4__10__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_14__10__q ;
wire Xd_0__inst_r_sum1_13__10__q ;
wire Xd_0__inst_r_sum1_12__10__q ;
wire Xd_0__inst_r_sum1_11__10__q ;
wire Xd_0__inst_r_sum1_10__10__q ;
wire Xd_0__inst_r_sum1_9__10__q ;
wire Xd_0__inst_r_sum1_8__11__q ;
wire Xd_0__inst_r_sum1_7__11__q ;
wire Xd_0__inst_r_sum1_6__11__q ;
wire Xd_0__inst_r_sum1_5__11__q ;
wire Xd_0__inst_r_sum1_4__11__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_14__11__q ;
wire Xd_0__inst_r_sum1_13__11__q ;
wire Xd_0__inst_r_sum1_12__11__q ;
wire Xd_0__inst_r_sum1_11__11__q ;
wire Xd_0__inst_r_sum1_10__11__q ;
wire Xd_0__inst_r_sum1_9__11__q ;
wire Xd_0__inst_product_30__0__q ;
wire Xd_0__inst_product_31__0__q ;
wire Xd_0__inst_product_30__1__q ;
wire Xd_0__inst_product_31__1__q ;
wire Xd_0__inst_product_30__2__q ;
wire Xd_0__inst_product_31__2__q ;
wire Xd_0__inst_product_30__3__q ;
wire Xd_0__inst_product_31__3__q ;
wire Xd_0__inst_product_30__4__q ;
wire Xd_0__inst_product_31__4__q ;
wire Xd_0__inst_product_30__5__q ;
wire Xd_0__inst_product_31__5__q ;
wire Xd_0__inst_product_30__6__q ;
wire Xd_0__inst_product_31__6__q ;
wire Xd_0__inst_product_30__7__q ;
wire Xd_0__inst_product_31__7__q ;
wire Xd_0__inst_product_30__8__q ;
wire Xd_0__inst_product_31__8__q ;
wire Xd_0__inst_product_30__9__q ;
wire Xd_0__inst_product_31__9__q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_product_16__0__q ;
wire Xd_0__inst_product_17__0__q ;
wire Xd_0__inst_product_14__0__q ;
wire Xd_0__inst_product_15__0__q ;
wire Xd_0__inst_product_12__0__q ;
wire Xd_0__inst_product_13__0__q ;
wire Xd_0__inst_product_10__0__q ;
wire Xd_0__inst_product_11__0__q ;
wire Xd_0__inst_product_8__0__q ;
wire Xd_0__inst_product_9__0__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product_28__0__q ;
wire Xd_0__inst_product_29__0__q ;
wire Xd_0__inst_product_26__0__q ;
wire Xd_0__inst_product_27__0__q ;
wire Xd_0__inst_product_24__0__q ;
wire Xd_0__inst_product_25__0__q ;
wire Xd_0__inst_product_22__0__q ;
wire Xd_0__inst_product_23__0__q ;
wire Xd_0__inst_product_20__0__q ;
wire Xd_0__inst_product_21__0__q ;
wire Xd_0__inst_product_18__0__q ;
wire Xd_0__inst_product_19__0__q ;
wire Xd_0__inst_product1_30__0__q ;
wire Xd_0__inst_product1_31__0__q ;
wire Xd_0__inst_product_16__1__q ;
wire Xd_0__inst_product_17__1__q ;
wire Xd_0__inst_product_14__1__q ;
wire Xd_0__inst_product_15__1__q ;
wire Xd_0__inst_product_12__1__q ;
wire Xd_0__inst_product_13__1__q ;
wire Xd_0__inst_product_10__1__q ;
wire Xd_0__inst_product_11__1__q ;
wire Xd_0__inst_product_8__1__q ;
wire Xd_0__inst_product_9__1__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product_28__1__q ;
wire Xd_0__inst_product_29__1__q ;
wire Xd_0__inst_product_26__1__q ;
wire Xd_0__inst_product_27__1__q ;
wire Xd_0__inst_product_24__1__q ;
wire Xd_0__inst_product_25__1__q ;
wire Xd_0__inst_product_22__1__q ;
wire Xd_0__inst_product_23__1__q ;
wire Xd_0__inst_product_20__1__q ;
wire Xd_0__inst_product_21__1__q ;
wire Xd_0__inst_product_18__1__q ;
wire Xd_0__inst_product_19__1__q ;
wire Xd_0__inst_product1_30__1__q ;
wire Xd_0__inst_product1_31__1__q ;
wire Xd_0__inst_product_16__2__q ;
wire Xd_0__inst_product_17__2__q ;
wire Xd_0__inst_product_14__2__q ;
wire Xd_0__inst_product_15__2__q ;
wire Xd_0__inst_product_12__2__q ;
wire Xd_0__inst_product_13__2__q ;
wire Xd_0__inst_product_10__2__q ;
wire Xd_0__inst_product_11__2__q ;
wire Xd_0__inst_product_8__2__q ;
wire Xd_0__inst_product_9__2__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product_28__2__q ;
wire Xd_0__inst_product_29__2__q ;
wire Xd_0__inst_product_26__2__q ;
wire Xd_0__inst_product_27__2__q ;
wire Xd_0__inst_product_24__2__q ;
wire Xd_0__inst_product_25__2__q ;
wire Xd_0__inst_product_22__2__q ;
wire Xd_0__inst_product_23__2__q ;
wire Xd_0__inst_product_20__2__q ;
wire Xd_0__inst_product_21__2__q ;
wire Xd_0__inst_product_18__2__q ;
wire Xd_0__inst_product_19__2__q ;
wire Xd_0__inst_product1_30__2__q ;
wire Xd_0__inst_product1_31__2__q ;
wire Xd_0__inst_product_16__3__q ;
wire Xd_0__inst_product_17__3__q ;
wire Xd_0__inst_product_14__3__q ;
wire Xd_0__inst_product_15__3__q ;
wire Xd_0__inst_product_12__3__q ;
wire Xd_0__inst_product_13__3__q ;
wire Xd_0__inst_product_10__3__q ;
wire Xd_0__inst_product_11__3__q ;
wire Xd_0__inst_product_8__3__q ;
wire Xd_0__inst_product_9__3__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product_28__3__q ;
wire Xd_0__inst_product_29__3__q ;
wire Xd_0__inst_product_26__3__q ;
wire Xd_0__inst_product_27__3__q ;
wire Xd_0__inst_product_24__3__q ;
wire Xd_0__inst_product_25__3__q ;
wire Xd_0__inst_product_22__3__q ;
wire Xd_0__inst_product_23__3__q ;
wire Xd_0__inst_product_20__3__q ;
wire Xd_0__inst_product_21__3__q ;
wire Xd_0__inst_product_18__3__q ;
wire Xd_0__inst_product_19__3__q ;
wire Xd_0__inst_product_16__4__q ;
wire Xd_0__inst_product_17__4__q ;
wire Xd_0__inst_product_14__4__q ;
wire Xd_0__inst_product_15__4__q ;
wire Xd_0__inst_product_12__4__q ;
wire Xd_0__inst_product_13__4__q ;
wire Xd_0__inst_product_10__4__q ;
wire Xd_0__inst_product_11__4__q ;
wire Xd_0__inst_product_8__4__q ;
wire Xd_0__inst_product_9__4__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product_28__4__q ;
wire Xd_0__inst_product_29__4__q ;
wire Xd_0__inst_product_26__4__q ;
wire Xd_0__inst_product_27__4__q ;
wire Xd_0__inst_product_24__4__q ;
wire Xd_0__inst_product_25__4__q ;
wire Xd_0__inst_product_22__4__q ;
wire Xd_0__inst_product_23__4__q ;
wire Xd_0__inst_product_20__4__q ;
wire Xd_0__inst_product_21__4__q ;
wire Xd_0__inst_product_18__4__q ;
wire Xd_0__inst_product_19__4__q ;
wire Xd_0__inst_product_16__5__q ;
wire Xd_0__inst_product_17__5__q ;
wire Xd_0__inst_product_14__5__q ;
wire Xd_0__inst_product_15__5__q ;
wire Xd_0__inst_product_12__5__q ;
wire Xd_0__inst_product_13__5__q ;
wire Xd_0__inst_product_10__5__q ;
wire Xd_0__inst_product_11__5__q ;
wire Xd_0__inst_product_8__5__q ;
wire Xd_0__inst_product_9__5__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_28__5__q ;
wire Xd_0__inst_product_29__5__q ;
wire Xd_0__inst_product_26__5__q ;
wire Xd_0__inst_product_27__5__q ;
wire Xd_0__inst_product_24__5__q ;
wire Xd_0__inst_product_25__5__q ;
wire Xd_0__inst_product_22__5__q ;
wire Xd_0__inst_product_23__5__q ;
wire Xd_0__inst_product_20__5__q ;
wire Xd_0__inst_product_21__5__q ;
wire Xd_0__inst_product_18__5__q ;
wire Xd_0__inst_product_19__5__q ;
wire Xd_0__inst_product_16__6__q ;
wire Xd_0__inst_product_17__6__q ;
wire Xd_0__inst_product_14__6__q ;
wire Xd_0__inst_product_15__6__q ;
wire Xd_0__inst_product_12__6__q ;
wire Xd_0__inst_product_13__6__q ;
wire Xd_0__inst_product_10__6__q ;
wire Xd_0__inst_product_11__6__q ;
wire Xd_0__inst_product_8__6__q ;
wire Xd_0__inst_product_9__6__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_28__6__q ;
wire Xd_0__inst_product_29__6__q ;
wire Xd_0__inst_product_26__6__q ;
wire Xd_0__inst_product_27__6__q ;
wire Xd_0__inst_product_24__6__q ;
wire Xd_0__inst_product_25__6__q ;
wire Xd_0__inst_product_22__6__q ;
wire Xd_0__inst_product_23__6__q ;
wire Xd_0__inst_product_20__6__q ;
wire Xd_0__inst_product_21__6__q ;
wire Xd_0__inst_product_18__6__q ;
wire Xd_0__inst_product_19__6__q ;
wire Xd_0__inst_product_16__7__q ;
wire Xd_0__inst_product_17__7__q ;
wire Xd_0__inst_product_14__7__q ;
wire Xd_0__inst_product_15__7__q ;
wire Xd_0__inst_product_12__7__q ;
wire Xd_0__inst_product_13__7__q ;
wire Xd_0__inst_product_10__7__q ;
wire Xd_0__inst_product_11__7__q ;
wire Xd_0__inst_product_8__7__q ;
wire Xd_0__inst_product_9__7__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_28__7__q ;
wire Xd_0__inst_product_29__7__q ;
wire Xd_0__inst_product_26__7__q ;
wire Xd_0__inst_product_27__7__q ;
wire Xd_0__inst_product_24__7__q ;
wire Xd_0__inst_product_25__7__q ;
wire Xd_0__inst_product_22__7__q ;
wire Xd_0__inst_product_23__7__q ;
wire Xd_0__inst_product_20__7__q ;
wire Xd_0__inst_product_21__7__q ;
wire Xd_0__inst_product_18__7__q ;
wire Xd_0__inst_product_19__7__q ;
wire Xd_0__inst_product_16__8__q ;
wire Xd_0__inst_product_17__8__q ;
wire Xd_0__inst_product_14__8__q ;
wire Xd_0__inst_product_15__8__q ;
wire Xd_0__inst_product_12__8__q ;
wire Xd_0__inst_product_13__8__q ;
wire Xd_0__inst_product_10__8__q ;
wire Xd_0__inst_product_11__8__q ;
wire Xd_0__inst_product_8__8__q ;
wire Xd_0__inst_product_9__8__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_28__8__q ;
wire Xd_0__inst_product_29__8__q ;
wire Xd_0__inst_product_26__8__q ;
wire Xd_0__inst_product_27__8__q ;
wire Xd_0__inst_product_24__8__q ;
wire Xd_0__inst_product_25__8__q ;
wire Xd_0__inst_product_22__8__q ;
wire Xd_0__inst_product_23__8__q ;
wire Xd_0__inst_product_20__8__q ;
wire Xd_0__inst_product_21__8__q ;
wire Xd_0__inst_product_18__8__q ;
wire Xd_0__inst_product_19__8__q ;
wire Xd_0__inst_product_16__9__q ;
wire Xd_0__inst_product_17__9__q ;
wire Xd_0__inst_product_14__9__q ;
wire Xd_0__inst_product_15__9__q ;
wire Xd_0__inst_product_12__9__q ;
wire Xd_0__inst_product_13__9__q ;
wire Xd_0__inst_product_10__9__q ;
wire Xd_0__inst_product_11__9__q ;
wire Xd_0__inst_product_8__9__q ;
wire Xd_0__inst_product_9__9__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_28__9__q ;
wire Xd_0__inst_product_29__9__q ;
wire Xd_0__inst_product_26__9__q ;
wire Xd_0__inst_product_27__9__q ;
wire Xd_0__inst_product_24__9__q ;
wire Xd_0__inst_product_25__9__q ;
wire Xd_0__inst_product_22__9__q ;
wire Xd_0__inst_product_23__9__q ;
wire Xd_0__inst_product_20__9__q ;
wire Xd_0__inst_product_21__9__q ;
wire Xd_0__inst_product_18__9__q ;
wire Xd_0__inst_product_19__9__q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_25_0_q ;
wire Xd_0__inst_mult_25_1_q ;
wire Xd_0__inst_mult_24_0_q ;
wire Xd_0__inst_mult_24_1_q ;
wire Xd_0__inst_mult_27_0_q ;
wire Xd_0__inst_mult_27_1_q ;
wire Xd_0__inst_mult_26_0_q ;
wire Xd_0__inst_mult_26_1_q ;
wire Xd_0__inst_mult_29_0_q ;
wire Xd_0__inst_mult_29_1_q ;
wire Xd_0__inst_mult_28_0_q ;
wire Xd_0__inst_mult_28_1_q ;
wire Xd_0__inst_mult_31_0_q ;
wire Xd_0__inst_mult_31_1_q ;
wire Xd_0__inst_mult_20_0_q ;
wire Xd_0__inst_mult_20_1_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_1_0_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_11_0_q ;
wire Xd_0__inst_mult_11_1_q ;
wire Xd_0__inst_mult_30_0_q ;
wire Xd_0__inst_mult_30_1_q ;
wire Xd_0__inst_mult_23_0_q ;
wire Xd_0__inst_mult_23_1_q ;
wire Xd_0__inst_mult_22_0_q ;
wire Xd_0__inst_mult_22_1_q ;
wire Xd_0__inst_product1_16__0__q ;
wire Xd_0__inst_product1_17__0__q ;
wire Xd_0__inst_product1_14__0__q ;
wire Xd_0__inst_product1_15__0__q ;
wire Xd_0__inst_product1_12__0__q ;
wire Xd_0__inst_product1_13__0__q ;
wire Xd_0__inst_product1_10__0__q ;
wire Xd_0__inst_product1_11__0__q ;
wire Xd_0__inst_product1_8__0__q ;
wire Xd_0__inst_product1_9__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_28__0__q ;
wire Xd_0__inst_product1_29__0__q ;
wire Xd_0__inst_product1_26__0__q ;
wire Xd_0__inst_product1_27__0__q ;
wire Xd_0__inst_product1_24__0__q ;
wire Xd_0__inst_product1_25__0__q ;
wire Xd_0__inst_product1_22__0__q ;
wire Xd_0__inst_product1_23__0__q ;
wire Xd_0__inst_product1_20__0__q ;
wire Xd_0__inst_product1_21__0__q ;
wire Xd_0__inst_product1_18__0__q ;
wire Xd_0__inst_product1_19__0__q ;
wire Xd_0__inst_product1_16__1__q ;
wire Xd_0__inst_product1_17__1__q ;
wire Xd_0__inst_product1_14__1__q ;
wire Xd_0__inst_product1_15__1__q ;
wire Xd_0__inst_product1_12__1__q ;
wire Xd_0__inst_product1_13__1__q ;
wire Xd_0__inst_product1_10__1__q ;
wire Xd_0__inst_product1_11__1__q ;
wire Xd_0__inst_product1_8__1__q ;
wire Xd_0__inst_product1_9__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_28__1__q ;
wire Xd_0__inst_product1_29__1__q ;
wire Xd_0__inst_product1_26__1__q ;
wire Xd_0__inst_product1_27__1__q ;
wire Xd_0__inst_product1_24__1__q ;
wire Xd_0__inst_product1_25__1__q ;
wire Xd_0__inst_product1_22__1__q ;
wire Xd_0__inst_product1_23__1__q ;
wire Xd_0__inst_product1_20__1__q ;
wire Xd_0__inst_product1_21__1__q ;
wire Xd_0__inst_product1_18__1__q ;
wire Xd_0__inst_product1_19__1__q ;
wire Xd_0__inst_product1_16__2__q ;
wire Xd_0__inst_product1_17__2__q ;
wire Xd_0__inst_product1_14__2__q ;
wire Xd_0__inst_product1_15__2__q ;
wire Xd_0__inst_product1_12__2__q ;
wire Xd_0__inst_product1_13__2__q ;
wire Xd_0__inst_product1_10__2__q ;
wire Xd_0__inst_product1_11__2__q ;
wire Xd_0__inst_product1_8__2__q ;
wire Xd_0__inst_product1_9__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_product1_28__2__q ;
wire Xd_0__inst_product1_29__2__q ;
wire Xd_0__inst_product1_26__2__q ;
wire Xd_0__inst_product1_27__2__q ;
wire Xd_0__inst_product1_24__2__q ;
wire Xd_0__inst_product1_25__2__q ;
wire Xd_0__inst_product1_22__2__q ;
wire Xd_0__inst_product1_23__2__q ;
wire Xd_0__inst_product1_20__2__q ;
wire Xd_0__inst_product1_21__2__q ;
wire Xd_0__inst_product1_18__2__q ;
wire Xd_0__inst_product1_19__2__q ;
wire Xd_0__inst_mult_30_4_q ;
wire Xd_0__inst_mult_30_2_q ;
wire Xd_0__inst_mult_30_5_q ;
wire Xd_0__inst_mult_31_4_q ;
wire Xd_0__inst_mult_31_2_q ;
wire Xd_0__inst_mult_31_5_q ;
wire Xd_0__inst_mult_30_6_q ;
wire Xd_0__inst_mult_30_7_q ;
wire Xd_0__inst_mult_31_6_q ;
wire Xd_0__inst_mult_31_7_q ;
wire Xd_0__inst_mult_30_8_q ;
wire Xd_0__inst_mult_30_9_q ;
wire Xd_0__inst_mult_30_10_q ;
wire Xd_0__inst_mult_31_8_q ;
wire Xd_0__inst_mult_31_9_q ;
wire Xd_0__inst_mult_31_10_q ;
wire Xd_0__inst_mult_30_11_q ;
wire Xd_0__inst_mult_30_12_q ;
wire Xd_0__inst_mult_31_11_q ;
wire Xd_0__inst_mult_31_12_q ;
wire Xd_0__inst_mult_30_13_q ;
wire Xd_0__inst_mult_31_13_q ;
wire Xd_0__inst_mult_30_14_q ;
wire Xd_0__inst_mult_30_15_q ;
wire Xd_0__inst_mult_31_14_q ;
wire Xd_0__inst_mult_31_15_q ;
wire Xd_0__inst_mult_16_4_q ;
wire Xd_0__inst_mult_16_2_q ;
wire Xd_0__inst_mult_16_5_q ;
wire Xd_0__inst_mult_17_4_q ;
wire Xd_0__inst_mult_17_2_q ;
wire Xd_0__inst_mult_17_5_q ;
wire Xd_0__inst_mult_14_4_q ;
wire Xd_0__inst_mult_14_2_q ;
wire Xd_0__inst_mult_14_5_q ;
wire Xd_0__inst_mult_15_4_q ;
wire Xd_0__inst_mult_15_2_q ;
wire Xd_0__inst_mult_15_5_q ;
wire Xd_0__inst_mult_12_4_q ;
wire Xd_0__inst_mult_12_2_q ;
wire Xd_0__inst_mult_12_5_q ;
wire Xd_0__inst_mult_13_4_q ;
wire Xd_0__inst_mult_13_2_q ;
wire Xd_0__inst_mult_13_5_q ;
wire Xd_0__inst_mult_10_4_q ;
wire Xd_0__inst_mult_10_2_q ;
wire Xd_0__inst_mult_10_5_q ;
wire Xd_0__inst_mult_11_4_q ;
wire Xd_0__inst_mult_11_2_q ;
wire Xd_0__inst_mult_11_5_q ;
wire Xd_0__inst_mult_8_4_q ;
wire Xd_0__inst_mult_8_2_q ;
wire Xd_0__inst_mult_8_5_q ;
wire Xd_0__inst_mult_9_4_q ;
wire Xd_0__inst_mult_9_2_q ;
wire Xd_0__inst_mult_9_5_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_28_4_q ;
wire Xd_0__inst_mult_28_2_q ;
wire Xd_0__inst_mult_28_5_q ;
wire Xd_0__inst_mult_29_4_q ;
wire Xd_0__inst_mult_29_2_q ;
wire Xd_0__inst_mult_29_5_q ;
wire Xd_0__inst_mult_26_4_q ;
wire Xd_0__inst_mult_26_2_q ;
wire Xd_0__inst_mult_26_5_q ;
wire Xd_0__inst_mult_27_4_q ;
wire Xd_0__inst_mult_27_2_q ;
wire Xd_0__inst_mult_27_5_q ;
wire Xd_0__inst_mult_24_4_q ;
wire Xd_0__inst_mult_24_2_q ;
wire Xd_0__inst_mult_24_5_q ;
wire Xd_0__inst_mult_25_4_q ;
wire Xd_0__inst_mult_25_2_q ;
wire Xd_0__inst_mult_25_5_q ;
wire Xd_0__inst_mult_22_4_q ;
wire Xd_0__inst_mult_22_2_q ;
wire Xd_0__inst_mult_22_5_q ;
wire Xd_0__inst_mult_23_4_q ;
wire Xd_0__inst_mult_23_2_q ;
wire Xd_0__inst_mult_23_5_q ;
wire Xd_0__inst_mult_20_4_q ;
wire Xd_0__inst_mult_20_2_q ;
wire Xd_0__inst_mult_20_5_q ;
wire Xd_0__inst_mult_21_4_q ;
wire Xd_0__inst_mult_21_2_q ;
wire Xd_0__inst_mult_21_5_q ;
wire Xd_0__inst_mult_18_4_q ;
wire Xd_0__inst_mult_18_2_q ;
wire Xd_0__inst_mult_18_5_q ;
wire Xd_0__inst_mult_19_4_q ;
wire Xd_0__inst_mult_19_2_q ;
wire Xd_0__inst_mult_19_5_q ;
wire Xd_0__inst_mult_30_3_q ;
wire Xd_0__inst_mult_31_3_q ;
wire Xd_0__inst_mult_16_6_q ;
wire Xd_0__inst_mult_16_7_q ;
wire Xd_0__inst_mult_17_6_q ;
wire Xd_0__inst_mult_17_7_q ;
wire Xd_0__inst_mult_14_6_q ;
wire Xd_0__inst_mult_14_7_q ;
wire Xd_0__inst_mult_15_6_q ;
wire Xd_0__inst_mult_15_7_q ;
wire Xd_0__inst_mult_12_6_q ;
wire Xd_0__inst_mult_12_7_q ;
wire Xd_0__inst_mult_13_6_q ;
wire Xd_0__inst_mult_13_7_q ;
wire Xd_0__inst_mult_10_6_q ;
wire Xd_0__inst_mult_10_7_q ;
wire Xd_0__inst_mult_11_6_q ;
wire Xd_0__inst_mult_11_7_q ;
wire Xd_0__inst_mult_8_6_q ;
wire Xd_0__inst_mult_8_7_q ;
wire Xd_0__inst_mult_9_6_q ;
wire Xd_0__inst_mult_9_7_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_28_6_q ;
wire Xd_0__inst_mult_28_7_q ;
wire Xd_0__inst_mult_29_6_q ;
wire Xd_0__inst_mult_29_7_q ;
wire Xd_0__inst_mult_26_6_q ;
wire Xd_0__inst_mult_26_7_q ;
wire Xd_0__inst_mult_27_6_q ;
wire Xd_0__inst_mult_27_7_q ;
wire Xd_0__inst_mult_24_6_q ;
wire Xd_0__inst_mult_24_7_q ;
wire Xd_0__inst_mult_25_6_q ;
wire Xd_0__inst_mult_25_7_q ;
wire Xd_0__inst_mult_22_6_q ;
wire Xd_0__inst_mult_22_7_q ;
wire Xd_0__inst_mult_23_6_q ;
wire Xd_0__inst_mult_23_7_q ;
wire Xd_0__inst_mult_20_6_q ;
wire Xd_0__inst_mult_20_7_q ;
wire Xd_0__inst_mult_21_6_q ;
wire Xd_0__inst_mult_21_7_q ;
wire Xd_0__inst_mult_18_6_q ;
wire Xd_0__inst_mult_18_7_q ;
wire Xd_0__inst_mult_19_6_q ;
wire Xd_0__inst_mult_19_7_q ;
wire Xd_0__inst_mult_16_8_q ;
wire Xd_0__inst_mult_16_9_q ;
wire Xd_0__inst_mult_16_10_q ;
wire Xd_0__inst_mult_17_8_q ;
wire Xd_0__inst_mult_17_9_q ;
wire Xd_0__inst_mult_17_10_q ;
wire Xd_0__inst_mult_14_8_q ;
wire Xd_0__inst_mult_14_9_q ;
wire Xd_0__inst_mult_14_10_q ;
wire Xd_0__inst_mult_15_8_q ;
wire Xd_0__inst_mult_15_9_q ;
wire Xd_0__inst_mult_15_10_q ;
wire Xd_0__inst_mult_12_8_q ;
wire Xd_0__inst_mult_12_9_q ;
wire Xd_0__inst_mult_12_10_q ;
wire Xd_0__inst_mult_13_8_q ;
wire Xd_0__inst_mult_13_9_q ;
wire Xd_0__inst_mult_13_10_q ;
wire Xd_0__inst_mult_10_8_q ;
wire Xd_0__inst_mult_10_9_q ;
wire Xd_0__inst_mult_10_10_q ;
wire Xd_0__inst_mult_11_8_q ;
wire Xd_0__inst_mult_11_9_q ;
wire Xd_0__inst_mult_11_10_q ;
wire Xd_0__inst_mult_8_8_q ;
wire Xd_0__inst_mult_8_9_q ;
wire Xd_0__inst_mult_8_10_q ;
wire Xd_0__inst_mult_9_8_q ;
wire Xd_0__inst_mult_9_9_q ;
wire Xd_0__inst_mult_9_10_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_28_8_q ;
wire Xd_0__inst_mult_28_9_q ;
wire Xd_0__inst_mult_28_10_q ;
wire Xd_0__inst_mult_29_8_q ;
wire Xd_0__inst_mult_29_9_q ;
wire Xd_0__inst_mult_29_10_q ;
wire Xd_0__inst_mult_26_8_q ;
wire Xd_0__inst_mult_26_9_q ;
wire Xd_0__inst_mult_26_10_q ;
wire Xd_0__inst_mult_27_8_q ;
wire Xd_0__inst_mult_27_9_q ;
wire Xd_0__inst_mult_27_10_q ;
wire Xd_0__inst_mult_24_8_q ;
wire Xd_0__inst_mult_24_9_q ;
wire Xd_0__inst_mult_24_10_q ;
wire Xd_0__inst_mult_25_8_q ;
wire Xd_0__inst_mult_25_9_q ;
wire Xd_0__inst_mult_25_10_q ;
wire Xd_0__inst_mult_22_8_q ;
wire Xd_0__inst_mult_22_9_q ;
wire Xd_0__inst_mult_22_10_q ;
wire Xd_0__inst_mult_23_8_q ;
wire Xd_0__inst_mult_23_9_q ;
wire Xd_0__inst_mult_23_10_q ;
wire Xd_0__inst_mult_20_8_q ;
wire Xd_0__inst_mult_20_9_q ;
wire Xd_0__inst_mult_20_10_q ;
wire Xd_0__inst_mult_21_8_q ;
wire Xd_0__inst_mult_21_9_q ;
wire Xd_0__inst_mult_21_10_q ;
wire Xd_0__inst_mult_18_8_q ;
wire Xd_0__inst_mult_18_9_q ;
wire Xd_0__inst_mult_18_10_q ;
wire Xd_0__inst_mult_19_8_q ;
wire Xd_0__inst_mult_19_9_q ;
wire Xd_0__inst_mult_19_10_q ;
wire Xd_0__inst_mult_16_11_q ;
wire Xd_0__inst_mult_16_12_q ;
wire Xd_0__inst_mult_17_11_q ;
wire Xd_0__inst_mult_17_12_q ;
wire Xd_0__inst_mult_14_11_q ;
wire Xd_0__inst_mult_14_12_q ;
wire Xd_0__inst_mult_15_11_q ;
wire Xd_0__inst_mult_15_12_q ;
wire Xd_0__inst_mult_12_11_q ;
wire Xd_0__inst_mult_12_12_q ;
wire Xd_0__inst_mult_13_11_q ;
wire Xd_0__inst_mult_13_12_q ;
wire Xd_0__inst_mult_10_11_q ;
wire Xd_0__inst_mult_10_12_q ;
wire Xd_0__inst_mult_11_11_q ;
wire Xd_0__inst_mult_11_12_q ;
wire Xd_0__inst_mult_8_11_q ;
wire Xd_0__inst_mult_8_12_q ;
wire Xd_0__inst_mult_9_11_q ;
wire Xd_0__inst_mult_9_12_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_28_11_q ;
wire Xd_0__inst_mult_28_12_q ;
wire Xd_0__inst_mult_29_11_q ;
wire Xd_0__inst_mult_29_12_q ;
wire Xd_0__inst_mult_26_11_q ;
wire Xd_0__inst_mult_26_12_q ;
wire Xd_0__inst_mult_27_11_q ;
wire Xd_0__inst_mult_27_12_q ;
wire Xd_0__inst_mult_24_11_q ;
wire Xd_0__inst_mult_24_12_q ;
wire Xd_0__inst_mult_25_11_q ;
wire Xd_0__inst_mult_25_12_q ;
wire Xd_0__inst_mult_22_11_q ;
wire Xd_0__inst_mult_22_12_q ;
wire Xd_0__inst_mult_23_11_q ;
wire Xd_0__inst_mult_23_12_q ;
wire Xd_0__inst_mult_20_11_q ;
wire Xd_0__inst_mult_20_12_q ;
wire Xd_0__inst_mult_21_11_q ;
wire Xd_0__inst_mult_21_12_q ;
wire Xd_0__inst_mult_18_11_q ;
wire Xd_0__inst_mult_18_12_q ;
wire Xd_0__inst_mult_19_11_q ;
wire Xd_0__inst_mult_19_12_q ;
wire Xd_0__inst_mult_16_0_q ;
wire Xd_0__inst_mult_16_13_q ;
wire Xd_0__inst_mult_17_0_q ;
wire Xd_0__inst_mult_17_13_q ;
wire Xd_0__inst_mult_14_0_q ;
wire Xd_0__inst_mult_14_13_q ;
wire Xd_0__inst_mult_15_0_q ;
wire Xd_0__inst_mult_15_13_q ;
wire Xd_0__inst_mult_12_0_q ;
wire Xd_0__inst_mult_12_13_q ;
wire Xd_0__inst_mult_13_0_q ;
wire Xd_0__inst_mult_13_13_q ;
wire Xd_0__inst_mult_10_0_q ;
wire Xd_0__inst_mult_10_13_q ;
wire Xd_0__inst_mult_11_13_q ;
wire Xd_0__inst_mult_8_0_q ;
wire Xd_0__inst_mult_8_13_q ;
wire Xd_0__inst_mult_9_0_q ;
wire Xd_0__inst_mult_9_13_q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_28_13_q ;
wire Xd_0__inst_mult_29_13_q ;
wire Xd_0__inst_mult_26_13_q ;
wire Xd_0__inst_mult_27_13_q ;
wire Xd_0__inst_mult_24_13_q ;
wire Xd_0__inst_mult_25_13_q ;
wire Xd_0__inst_mult_22_13_q ;
wire Xd_0__inst_mult_23_13_q ;
wire Xd_0__inst_mult_20_13_q ;
wire Xd_0__inst_mult_21_0_q ;
wire Xd_0__inst_mult_21_13_q ;
wire Xd_0__inst_mult_18_0_q ;
wire Xd_0__inst_mult_18_13_q ;
wire Xd_0__inst_mult_19_0_q ;
wire Xd_0__inst_mult_19_13_q ;
wire Xd_0__inst_mult_16_14_q ;
wire Xd_0__inst_mult_16_15_q ;
wire Xd_0__inst_mult_17_14_q ;
wire Xd_0__inst_mult_17_15_q ;
wire Xd_0__inst_mult_14_14_q ;
wire Xd_0__inst_mult_14_15_q ;
wire Xd_0__inst_mult_15_14_q ;
wire Xd_0__inst_mult_15_15_q ;
wire Xd_0__inst_mult_12_14_q ;
wire Xd_0__inst_mult_12_15_q ;
wire Xd_0__inst_mult_13_14_q ;
wire Xd_0__inst_mult_13_15_q ;
wire Xd_0__inst_mult_10_14_q ;
wire Xd_0__inst_mult_10_15_q ;
wire Xd_0__inst_mult_11_14_q ;
wire Xd_0__inst_mult_11_15_q ;
wire Xd_0__inst_mult_8_14_q ;
wire Xd_0__inst_mult_8_15_q ;
wire Xd_0__inst_mult_9_14_q ;
wire Xd_0__inst_mult_9_15_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_28_14_q ;
wire Xd_0__inst_mult_28_15_q ;
wire Xd_0__inst_mult_29_14_q ;
wire Xd_0__inst_mult_29_15_q ;
wire Xd_0__inst_mult_26_14_q ;
wire Xd_0__inst_mult_26_15_q ;
wire Xd_0__inst_mult_27_14_q ;
wire Xd_0__inst_mult_27_15_q ;
wire Xd_0__inst_mult_24_14_q ;
wire Xd_0__inst_mult_24_15_q ;
wire Xd_0__inst_mult_25_14_q ;
wire Xd_0__inst_mult_25_15_q ;
wire Xd_0__inst_mult_22_14_q ;
wire Xd_0__inst_mult_22_15_q ;
wire Xd_0__inst_mult_23_14_q ;
wire Xd_0__inst_mult_23_15_q ;
wire Xd_0__inst_mult_20_14_q ;
wire Xd_0__inst_mult_20_15_q ;
wire Xd_0__inst_mult_21_14_q ;
wire Xd_0__inst_mult_21_15_q ;
wire Xd_0__inst_mult_18_14_q ;
wire Xd_0__inst_mult_18_15_q ;
wire Xd_0__inst_mult_19_14_q ;
wire Xd_0__inst_mult_19_15_q ;
wire Xd_0__inst_mult_17_1_q ;
wire Xd_0__inst_mult_15_1_q ;
wire Xd_0__inst_mult_13_1_q ;
wire Xd_0__inst_mult_21_1_q ;
wire Xd_0__inst_mult_9_1_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_19_1_q ;
wire Xd_0__inst_mult_16_1_q ;
wire Xd_0__inst_mult_16_3_q ;
wire Xd_0__inst_mult_17_3_q ;
wire Xd_0__inst_mult_14_1_q ;
wire Xd_0__inst_mult_14_3_q ;
wire Xd_0__inst_mult_15_3_q ;
wire Xd_0__inst_mult_12_1_q ;
wire Xd_0__inst_mult_12_3_q ;
wire Xd_0__inst_mult_13_3_q ;
wire Xd_0__inst_mult_10_1_q ;
wire Xd_0__inst_mult_10_3_q ;
wire Xd_0__inst_mult_11_3_q ;
wire Xd_0__inst_mult_8_1_q ;
wire Xd_0__inst_mult_8_3_q ;
wire Xd_0__inst_mult_9_3_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_28_3_q ;
wire Xd_0__inst_mult_29_3_q ;
wire Xd_0__inst_mult_26_3_q ;
wire Xd_0__inst_mult_27_3_q ;
wire Xd_0__inst_mult_24_3_q ;
wire Xd_0__inst_mult_25_3_q ;
wire Xd_0__inst_mult_22_3_q ;
wire Xd_0__inst_mult_23_3_q ;
wire Xd_0__inst_mult_20_3_q ;
wire Xd_0__inst_mult_21_3_q ;
wire Xd_0__inst_mult_18_1_q ;
wire Xd_0__inst_mult_18_3_q ;
wire Xd_0__inst_mult_19_3_q ;
wire [0:31] Xd_0__inst_sign1 ;
wire [0:31] Xd_0__inst_sign ;
wire [15:0] Xd_0__inst_inst_inst_inst_dout ;
wire [11:0] Xd_0__inst_a1_9__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_10__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_11__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_12__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_13__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_14__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_6__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_7__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_8__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_15__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_4__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_5__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_3__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_2__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_1__adder1_inst_dout ;
wire [11:0] Xd_0__inst_a1_0__adder1_inst_dout ;


twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__0__q  $ (!Xd_0__inst_inst_inst_first_level_1__0__q ) ) + ( Xd_0__inst_mult_24_38  ) + ( Xd_0__inst_mult_24_37  ))
// Xd_0__inst_inst_inst_inst_add_0_2  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__0__q  $ (!Xd_0__inst_inst_inst_first_level_1__0__q ) ) + ( Xd_0__inst_mult_24_38  ) + ( Xd_0__inst_mult_24_37  ))
// Xd_0__inst_inst_inst_inst_add_0_3  = SHARE((Xd_0__inst_inst_inst_first_level_0__0__q  & Xd_0__inst_inst_inst_first_level_1__0__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__0__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_37 ),
	.sharein(Xd_0__inst_mult_24_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__1__q  $ (!Xd_0__inst_inst_inst_first_level_1__1__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_inst_add_0_6  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__1__q  $ (!Xd_0__inst_inst_inst_first_level_1__1__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_inst_add_0_7  = SHARE((Xd_0__inst_inst_inst_first_level_0__1__q  & Xd_0__inst_inst_inst_first_level_1__1__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__1__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__2__q  $ (!Xd_0__inst_inst_inst_first_level_1__2__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_inst_add_0_10  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__2__q  $ (!Xd_0__inst_inst_inst_first_level_1__2__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_inst_add_0_11  = SHARE((Xd_0__inst_inst_inst_first_level_0__2__q  & Xd_0__inst_inst_inst_first_level_1__2__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__2__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__3__q  $ (!Xd_0__inst_inst_inst_first_level_1__3__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_inst_add_0_14  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__3__q  $ (!Xd_0__inst_inst_inst_first_level_1__3__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_inst_add_0_15  = SHARE((Xd_0__inst_inst_inst_first_level_0__3__q  & Xd_0__inst_inst_inst_first_level_1__3__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__3__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__4__q  $ (!Xd_0__inst_inst_inst_first_level_1__4__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_inst_add_0_18  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__4__q  $ (!Xd_0__inst_inst_inst_first_level_1__4__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_inst_add_0_19  = SHARE((Xd_0__inst_inst_inst_first_level_0__4__q  & Xd_0__inst_inst_inst_first_level_1__4__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__4__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__5__q  $ (!Xd_0__inst_inst_inst_first_level_1__5__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_inst_add_0_22  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__5__q  $ (!Xd_0__inst_inst_inst_first_level_1__5__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_inst_add_0_23  = SHARE((Xd_0__inst_inst_inst_first_level_0__5__q  & Xd_0__inst_inst_inst_first_level_1__5__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__5__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__6__q  $ (!Xd_0__inst_inst_inst_first_level_1__6__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_inst_add_0_26  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__6__q  $ (!Xd_0__inst_inst_inst_first_level_1__6__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_inst_add_0_27  = SHARE((Xd_0__inst_inst_inst_first_level_0__6__q  & Xd_0__inst_inst_inst_first_level_1__6__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__6__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__7__q  $ (!Xd_0__inst_inst_inst_first_level_1__7__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_inst_add_0_30  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__7__q  $ (!Xd_0__inst_inst_inst_first_level_1__7__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_inst_add_0_31  = SHARE((Xd_0__inst_inst_inst_first_level_0__7__q  & Xd_0__inst_inst_inst_first_level_1__7__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__7__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__8__q  $ (!Xd_0__inst_inst_inst_first_level_1__8__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_inst_add_0_34  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__8__q  $ (!Xd_0__inst_inst_inst_first_level_1__8__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_inst_add_0_35  = SHARE((Xd_0__inst_inst_inst_first_level_0__8__q  & Xd_0__inst_inst_inst_first_level_1__8__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__8__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__9__q  $ (!Xd_0__inst_inst_inst_first_level_1__9__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_inst_add_0_38  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__9__q  $ (!Xd_0__inst_inst_inst_first_level_1__9__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_inst_add_0_39  = SHARE((Xd_0__inst_inst_inst_first_level_0__9__q  & Xd_0__inst_inst_inst_first_level_1__9__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__9__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__10__q  $ (!Xd_0__inst_inst_inst_first_level_1__10__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_inst_add_0_42  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__10__q  $ (!Xd_0__inst_inst_inst_first_level_1__10__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_inst_add_0_43  = SHARE((Xd_0__inst_inst_inst_first_level_0__10__q  & Xd_0__inst_inst_inst_first_level_1__10__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__10__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__11__q  $ (!Xd_0__inst_inst_inst_first_level_1__11__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_inst_add_0_46  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__11__q  $ (!Xd_0__inst_inst_inst_first_level_1__11__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_inst_add_0_47  = SHARE((Xd_0__inst_inst_inst_first_level_0__11__q  & Xd_0__inst_inst_inst_first_level_1__11__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__11__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__12__q  $ (!Xd_0__inst_inst_inst_first_level_1__12__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_inst_add_0_50  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__12__q  $ (!Xd_0__inst_inst_inst_first_level_1__12__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_inst_add_0_51  = SHARE((Xd_0__inst_inst_inst_first_level_0__12__q  & Xd_0__inst_inst_inst_first_level_1__12__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__12__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__13__q  $ (!Xd_0__inst_inst_inst_first_level_1__13__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_inst_add_0_54  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__13__q  $ (!Xd_0__inst_inst_inst_first_level_1__13__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_inst_add_0_55  = SHARE((Xd_0__inst_inst_inst_first_level_0__13__q  & Xd_0__inst_inst_inst_first_level_1__13__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__13__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__14__q  $ (!Xd_0__inst_inst_inst_first_level_1__14__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_inst_add_0_58  = CARRY(( !Xd_0__inst_inst_inst_first_level_0__14__q  $ (!Xd_0__inst_inst_inst_first_level_1__14__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_inst_add_0_59  = SHARE((Xd_0__inst_inst_inst_first_level_0__14__q  & Xd_0__inst_inst_inst_first_level_1__14__q ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__14__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000000000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_inst_inst_first_level_0__15__q  $ (!Xd_0__inst_inst_inst_first_level_1__15__q ) ) + ( Xd_0__inst_inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_inst_add_0_58  ))

	.dataa(!Xd_0__inst_inst_inst_first_level_0__15__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_inst_first_level_1__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_35 (
// Equation(s):
// Xd_0__inst_mult_24_36  = SUM(( GND ) + ( Xd_0__inst_mult_24_42  ) + ( Xd_0__inst_mult_24_41  ))
// Xd_0__inst_mult_24_37  = CARRY(( GND ) + ( Xd_0__inst_mult_24_42  ) + ( Xd_0__inst_mult_24_41  ))
// Xd_0__inst_mult_24_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_41 ),
	.sharein(Xd_0__inst_mult_24_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_36 ),
	.cout(Xd_0__inst_mult_24_37 ),
	.shareout(Xd_0__inst_mult_24_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_mult_20_38  ) + ( Xd_0__inst_mult_20_37  ))
// Xd_0__inst_inst_inst_add_0_2  = CARRY(( !Xd_0__inst_inst_first_level_2__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q  $ (Xd_0__inst_inst_first_level_0__0__q )) ) + ( Xd_0__inst_mult_20_38  ) + ( Xd_0__inst_mult_20_37  ))
// Xd_0__inst_inst_inst_add_0_3  = SHARE((!Xd_0__inst_inst_first_level_2__0__q  & (Xd_0__inst_inst_first_level_1__0__q  & Xd_0__inst_inst_first_level_0__0__q )) # (Xd_0__inst_inst_first_level_2__0__q  & ((Xd_0__inst_inst_first_level_0__0__q ) # 
// (Xd_0__inst_inst_first_level_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__0__q ),
	.datac(!Xd_0__inst_inst_first_level_1__0__q ),
	.datad(!Xd_0__inst_inst_first_level_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_37 ),
	.sharein(Xd_0__inst_mult_20_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_1 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__0__q  $ (!Xd_0__inst_inst_first_level_3__0__q  $ (Xd_0__inst_inst_first_level_5__0__q )) ) + ( Xd_0__inst_mult_23_38  ) + ( Xd_0__inst_mult_23_37  ))
// Xd_0__inst_inst_inst_add_3_2  = CARRY(( !Xd_0__inst_inst_first_level_4__0__q  $ (!Xd_0__inst_inst_first_level_3__0__q  $ (Xd_0__inst_inst_first_level_5__0__q )) ) + ( Xd_0__inst_mult_23_38  ) + ( Xd_0__inst_mult_23_37  ))
// Xd_0__inst_inst_inst_add_3_3  = SHARE((!Xd_0__inst_inst_first_level_4__0__q  & (Xd_0__inst_inst_first_level_3__0__q  & Xd_0__inst_inst_first_level_5__0__q )) # (Xd_0__inst_inst_first_level_4__0__q  & ((Xd_0__inst_inst_first_level_5__0__q ) # 
// (Xd_0__inst_inst_first_level_3__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__0__q ),
	.datac(!Xd_0__inst_inst_first_level_3__0__q ),
	.datad(!Xd_0__inst_inst_first_level_5__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_37 ),
	.sharein(Xd_0__inst_mult_23_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_2 ),
	.shareout(Xd_0__inst_inst_inst_add_3_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24 (
// Equation(s):
// Xd_0__inst_mult_24_40  = SUM(( (!din_a[148] & (((din_a[147] & din_b[145])))) # (din_a[148] & (!din_b[144] $ (((!din_a[147]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_24_45  ) + ( Xd_0__inst_mult_24_44  ))
// Xd_0__inst_mult_24_41  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[145])))) # (din_a[148] & (!din_b[144] $ (((!din_a[147]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_24_45  ) + ( Xd_0__inst_mult_24_44  ))
// Xd_0__inst_mult_24_42  = SHARE((din_a[148] & (din_b[144] & (din_a[147] & din_b[145]))))

	.dataa(!din_a[148]),
	.datab(!din_b[144]),
	.datac(!din_a[147]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_44 ),
	.sharein(Xd_0__inst_mult_24_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_40 ),
	.cout(Xd_0__inst_mult_24_41 ),
	.shareout(Xd_0__inst_mult_24_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_6  = CARRY(( !Xd_0__inst_inst_first_level_2__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q  $ (Xd_0__inst_inst_first_level_0__1__q )) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_7  = SHARE((!Xd_0__inst_inst_first_level_2__1__q  & (Xd_0__inst_inst_first_level_1__1__q  & Xd_0__inst_inst_first_level_0__1__q )) # (Xd_0__inst_inst_first_level_2__1__q  & ((Xd_0__inst_inst_first_level_0__1__q ) # 
// (Xd_0__inst_inst_first_level_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__1__q ),
	.datac(!Xd_0__inst_inst_first_level_1__1__q ),
	.datad(!Xd_0__inst_inst_first_level_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_5 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__1__q  $ (!Xd_0__inst_inst_first_level_3__1__q  $ (Xd_0__inst_inst_first_level_5__1__q )) ) + ( Xd_0__inst_inst_inst_add_3_3  ) + ( Xd_0__inst_inst_inst_add_3_2  ))
// Xd_0__inst_inst_inst_add_3_6  = CARRY(( !Xd_0__inst_inst_first_level_4__1__q  $ (!Xd_0__inst_inst_first_level_3__1__q  $ (Xd_0__inst_inst_first_level_5__1__q )) ) + ( Xd_0__inst_inst_inst_add_3_3  ) + ( Xd_0__inst_inst_inst_add_3_2  ))
// Xd_0__inst_inst_inst_add_3_7  = SHARE((!Xd_0__inst_inst_first_level_4__1__q  & (Xd_0__inst_inst_first_level_3__1__q  & Xd_0__inst_inst_first_level_5__1__q )) # (Xd_0__inst_inst_first_level_4__1__q  & ((Xd_0__inst_inst_first_level_5__1__q ) # 
// (Xd_0__inst_inst_first_level_3__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__1__q ),
	.datac(!Xd_0__inst_inst_first_level_3__1__q ),
	.datad(!Xd_0__inst_inst_first_level_5__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_2 ),
	.sharein(Xd_0__inst_inst_inst_add_3_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_5_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_6 ),
	.shareout(Xd_0__inst_inst_inst_add_3_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_10  = CARRY(( !Xd_0__inst_inst_first_level_2__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q  $ (Xd_0__inst_inst_first_level_0__2__q )) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_11  = SHARE((!Xd_0__inst_inst_first_level_2__2__q  & (Xd_0__inst_inst_first_level_1__2__q  & Xd_0__inst_inst_first_level_0__2__q )) # (Xd_0__inst_inst_first_level_2__2__q  & ((Xd_0__inst_inst_first_level_0__2__q ) # 
// (Xd_0__inst_inst_first_level_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__2__q ),
	.datac(!Xd_0__inst_inst_first_level_1__2__q ),
	.datad(!Xd_0__inst_inst_first_level_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_9 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__2__q  $ (!Xd_0__inst_inst_first_level_3__2__q  $ (Xd_0__inst_inst_first_level_5__2__q )) ) + ( Xd_0__inst_inst_inst_add_3_7  ) + ( Xd_0__inst_inst_inst_add_3_6  ))
// Xd_0__inst_inst_inst_add_3_10  = CARRY(( !Xd_0__inst_inst_first_level_4__2__q  $ (!Xd_0__inst_inst_first_level_3__2__q  $ (Xd_0__inst_inst_first_level_5__2__q )) ) + ( Xd_0__inst_inst_inst_add_3_7  ) + ( Xd_0__inst_inst_inst_add_3_6  ))
// Xd_0__inst_inst_inst_add_3_11  = SHARE((!Xd_0__inst_inst_first_level_4__2__q  & (Xd_0__inst_inst_first_level_3__2__q  & Xd_0__inst_inst_first_level_5__2__q )) # (Xd_0__inst_inst_first_level_4__2__q  & ((Xd_0__inst_inst_first_level_5__2__q ) # 
// (Xd_0__inst_inst_first_level_3__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__2__q ),
	.datac(!Xd_0__inst_inst_first_level_3__2__q ),
	.datad(!Xd_0__inst_inst_first_level_5__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_6 ),
	.sharein(Xd_0__inst_inst_inst_add_3_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_9_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_10 ),
	.shareout(Xd_0__inst_inst_inst_add_3_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_14  = CARRY(( !Xd_0__inst_inst_first_level_2__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q  $ (Xd_0__inst_inst_first_level_0__3__q )) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_15  = SHARE((!Xd_0__inst_inst_first_level_2__3__q  & (Xd_0__inst_inst_first_level_1__3__q  & Xd_0__inst_inst_first_level_0__3__q )) # (Xd_0__inst_inst_first_level_2__3__q  & ((Xd_0__inst_inst_first_level_0__3__q ) # 
// (Xd_0__inst_inst_first_level_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__3__q ),
	.datac(!Xd_0__inst_inst_first_level_1__3__q ),
	.datad(!Xd_0__inst_inst_first_level_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_13 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__3__q  $ (!Xd_0__inst_inst_first_level_3__3__q  $ (Xd_0__inst_inst_first_level_5__3__q )) ) + ( Xd_0__inst_inst_inst_add_3_11  ) + ( Xd_0__inst_inst_inst_add_3_10  ))
// Xd_0__inst_inst_inst_add_3_14  = CARRY(( !Xd_0__inst_inst_first_level_4__3__q  $ (!Xd_0__inst_inst_first_level_3__3__q  $ (Xd_0__inst_inst_first_level_5__3__q )) ) + ( Xd_0__inst_inst_inst_add_3_11  ) + ( Xd_0__inst_inst_inst_add_3_10  ))
// Xd_0__inst_inst_inst_add_3_15  = SHARE((!Xd_0__inst_inst_first_level_4__3__q  & (Xd_0__inst_inst_first_level_3__3__q  & Xd_0__inst_inst_first_level_5__3__q )) # (Xd_0__inst_inst_first_level_4__3__q  & ((Xd_0__inst_inst_first_level_5__3__q ) # 
// (Xd_0__inst_inst_first_level_3__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__3__q ),
	.datac(!Xd_0__inst_inst_first_level_3__3__q ),
	.datad(!Xd_0__inst_inst_first_level_5__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_10 ),
	.sharein(Xd_0__inst_inst_inst_add_3_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_13_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_14 ),
	.shareout(Xd_0__inst_inst_inst_add_3_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_18  = CARRY(( !Xd_0__inst_inst_first_level_2__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q  $ (Xd_0__inst_inst_first_level_0__4__q )) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_19  = SHARE((!Xd_0__inst_inst_first_level_2__4__q  & (Xd_0__inst_inst_first_level_1__4__q  & Xd_0__inst_inst_first_level_0__4__q )) # (Xd_0__inst_inst_first_level_2__4__q  & ((Xd_0__inst_inst_first_level_0__4__q ) # 
// (Xd_0__inst_inst_first_level_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__4__q ),
	.datac(!Xd_0__inst_inst_first_level_1__4__q ),
	.datad(!Xd_0__inst_inst_first_level_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_17 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__4__q  $ (!Xd_0__inst_inst_first_level_3__4__q  $ (Xd_0__inst_inst_first_level_5__4__q )) ) + ( Xd_0__inst_inst_inst_add_3_15  ) + ( Xd_0__inst_inst_inst_add_3_14  ))
// Xd_0__inst_inst_inst_add_3_18  = CARRY(( !Xd_0__inst_inst_first_level_4__4__q  $ (!Xd_0__inst_inst_first_level_3__4__q  $ (Xd_0__inst_inst_first_level_5__4__q )) ) + ( Xd_0__inst_inst_inst_add_3_15  ) + ( Xd_0__inst_inst_inst_add_3_14  ))
// Xd_0__inst_inst_inst_add_3_19  = SHARE((!Xd_0__inst_inst_first_level_4__4__q  & (Xd_0__inst_inst_first_level_3__4__q  & Xd_0__inst_inst_first_level_5__4__q )) # (Xd_0__inst_inst_first_level_4__4__q  & ((Xd_0__inst_inst_first_level_5__4__q ) # 
// (Xd_0__inst_inst_first_level_3__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__4__q ),
	.datac(!Xd_0__inst_inst_first_level_3__4__q ),
	.datad(!Xd_0__inst_inst_first_level_5__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_14 ),
	.sharein(Xd_0__inst_inst_inst_add_3_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_17_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_18 ),
	.shareout(Xd_0__inst_inst_inst_add_3_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_22  = CARRY(( !Xd_0__inst_inst_first_level_2__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q  $ (Xd_0__inst_inst_first_level_0__5__q )) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_23  = SHARE((!Xd_0__inst_inst_first_level_2__5__q  & (Xd_0__inst_inst_first_level_1__5__q  & Xd_0__inst_inst_first_level_0__5__q )) # (Xd_0__inst_inst_first_level_2__5__q  & ((Xd_0__inst_inst_first_level_0__5__q ) # 
// (Xd_0__inst_inst_first_level_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__5__q ),
	.datac(!Xd_0__inst_inst_first_level_1__5__q ),
	.datad(!Xd_0__inst_inst_first_level_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_21 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__5__q  $ (!Xd_0__inst_inst_first_level_3__5__q  $ (Xd_0__inst_inst_first_level_5__5__q )) ) + ( Xd_0__inst_inst_inst_add_3_19  ) + ( Xd_0__inst_inst_inst_add_3_18  ))
// Xd_0__inst_inst_inst_add_3_22  = CARRY(( !Xd_0__inst_inst_first_level_4__5__q  $ (!Xd_0__inst_inst_first_level_3__5__q  $ (Xd_0__inst_inst_first_level_5__5__q )) ) + ( Xd_0__inst_inst_inst_add_3_19  ) + ( Xd_0__inst_inst_inst_add_3_18  ))
// Xd_0__inst_inst_inst_add_3_23  = SHARE((!Xd_0__inst_inst_first_level_4__5__q  & (Xd_0__inst_inst_first_level_3__5__q  & Xd_0__inst_inst_first_level_5__5__q )) # (Xd_0__inst_inst_first_level_4__5__q  & ((Xd_0__inst_inst_first_level_5__5__q ) # 
// (Xd_0__inst_inst_first_level_3__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__5__q ),
	.datac(!Xd_0__inst_inst_first_level_3__5__q ),
	.datad(!Xd_0__inst_inst_first_level_5__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_18 ),
	.sharein(Xd_0__inst_inst_inst_add_3_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_22 ),
	.shareout(Xd_0__inst_inst_inst_add_3_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_26  = CARRY(( !Xd_0__inst_inst_first_level_2__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q  $ (Xd_0__inst_inst_first_level_0__6__q )) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_27  = SHARE((!Xd_0__inst_inst_first_level_2__6__q  & (Xd_0__inst_inst_first_level_1__6__q  & Xd_0__inst_inst_first_level_0__6__q )) # (Xd_0__inst_inst_first_level_2__6__q  & ((Xd_0__inst_inst_first_level_0__6__q ) # 
// (Xd_0__inst_inst_first_level_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__6__q ),
	.datac(!Xd_0__inst_inst_first_level_1__6__q ),
	.datad(!Xd_0__inst_inst_first_level_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_25 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__6__q  $ (!Xd_0__inst_inst_first_level_3__6__q  $ (Xd_0__inst_inst_first_level_5__6__q )) ) + ( Xd_0__inst_inst_inst_add_3_23  ) + ( Xd_0__inst_inst_inst_add_3_22  ))
// Xd_0__inst_inst_inst_add_3_26  = CARRY(( !Xd_0__inst_inst_first_level_4__6__q  $ (!Xd_0__inst_inst_first_level_3__6__q  $ (Xd_0__inst_inst_first_level_5__6__q )) ) + ( Xd_0__inst_inst_inst_add_3_23  ) + ( Xd_0__inst_inst_inst_add_3_22  ))
// Xd_0__inst_inst_inst_add_3_27  = SHARE((!Xd_0__inst_inst_first_level_4__6__q  & (Xd_0__inst_inst_first_level_3__6__q  & Xd_0__inst_inst_first_level_5__6__q )) # (Xd_0__inst_inst_first_level_4__6__q  & ((Xd_0__inst_inst_first_level_5__6__q ) # 
// (Xd_0__inst_inst_first_level_3__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__6__q ),
	.datac(!Xd_0__inst_inst_first_level_3__6__q ),
	.datad(!Xd_0__inst_inst_first_level_5__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_22 ),
	.sharein(Xd_0__inst_inst_inst_add_3_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_25_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_26 ),
	.shareout(Xd_0__inst_inst_inst_add_3_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_30  = CARRY(( !Xd_0__inst_inst_first_level_2__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q  $ (Xd_0__inst_inst_first_level_0__7__q )) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_31  = SHARE((!Xd_0__inst_inst_first_level_2__7__q  & (Xd_0__inst_inst_first_level_1__7__q  & Xd_0__inst_inst_first_level_0__7__q )) # (Xd_0__inst_inst_first_level_2__7__q  & ((Xd_0__inst_inst_first_level_0__7__q ) # 
// (Xd_0__inst_inst_first_level_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__7__q ),
	.datac(!Xd_0__inst_inst_first_level_1__7__q ),
	.datad(!Xd_0__inst_inst_first_level_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_29 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__7__q  $ (!Xd_0__inst_inst_first_level_3__7__q  $ (Xd_0__inst_inst_first_level_5__7__q )) ) + ( Xd_0__inst_inst_inst_add_3_27  ) + ( Xd_0__inst_inst_inst_add_3_26  ))
// Xd_0__inst_inst_inst_add_3_30  = CARRY(( !Xd_0__inst_inst_first_level_4__7__q  $ (!Xd_0__inst_inst_first_level_3__7__q  $ (Xd_0__inst_inst_first_level_5__7__q )) ) + ( Xd_0__inst_inst_inst_add_3_27  ) + ( Xd_0__inst_inst_inst_add_3_26  ))
// Xd_0__inst_inst_inst_add_3_31  = SHARE((!Xd_0__inst_inst_first_level_4__7__q  & (Xd_0__inst_inst_first_level_3__7__q  & Xd_0__inst_inst_first_level_5__7__q )) # (Xd_0__inst_inst_first_level_4__7__q  & ((Xd_0__inst_inst_first_level_5__7__q ) # 
// (Xd_0__inst_inst_first_level_3__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__7__q ),
	.datac(!Xd_0__inst_inst_first_level_3__7__q ),
	.datad(!Xd_0__inst_inst_first_level_5__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_26 ),
	.sharein(Xd_0__inst_inst_inst_add_3_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_29_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_30 ),
	.shareout(Xd_0__inst_inst_inst_add_3_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_34  = CARRY(( !Xd_0__inst_inst_first_level_2__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q  $ (Xd_0__inst_inst_first_level_0__8__q )) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_35  = SHARE((!Xd_0__inst_inst_first_level_2__8__q  & (Xd_0__inst_inst_first_level_1__8__q  & Xd_0__inst_inst_first_level_0__8__q )) # (Xd_0__inst_inst_first_level_2__8__q  & ((Xd_0__inst_inst_first_level_0__8__q ) # 
// (Xd_0__inst_inst_first_level_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__8__q ),
	.datac(!Xd_0__inst_inst_first_level_1__8__q ),
	.datad(!Xd_0__inst_inst_first_level_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_33 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__8__q  $ (!Xd_0__inst_inst_first_level_3__8__q  $ (Xd_0__inst_inst_first_level_5__8__q )) ) + ( Xd_0__inst_inst_inst_add_3_31  ) + ( Xd_0__inst_inst_inst_add_3_30  ))
// Xd_0__inst_inst_inst_add_3_34  = CARRY(( !Xd_0__inst_inst_first_level_4__8__q  $ (!Xd_0__inst_inst_first_level_3__8__q  $ (Xd_0__inst_inst_first_level_5__8__q )) ) + ( Xd_0__inst_inst_inst_add_3_31  ) + ( Xd_0__inst_inst_inst_add_3_30  ))
// Xd_0__inst_inst_inst_add_3_35  = SHARE((!Xd_0__inst_inst_first_level_4__8__q  & (Xd_0__inst_inst_first_level_3__8__q  & Xd_0__inst_inst_first_level_5__8__q )) # (Xd_0__inst_inst_first_level_4__8__q  & ((Xd_0__inst_inst_first_level_5__8__q ) # 
// (Xd_0__inst_inst_first_level_3__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__8__q ),
	.datac(!Xd_0__inst_inst_first_level_3__8__q ),
	.datad(!Xd_0__inst_inst_first_level_5__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_30 ),
	.sharein(Xd_0__inst_inst_inst_add_3_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_33_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_34 ),
	.shareout(Xd_0__inst_inst_inst_add_3_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_38  = CARRY(( !Xd_0__inst_inst_first_level_2__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q  $ (Xd_0__inst_inst_first_level_0__9__q )) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_39  = SHARE((!Xd_0__inst_inst_first_level_2__9__q  & (Xd_0__inst_inst_first_level_1__9__q  & Xd_0__inst_inst_first_level_0__9__q )) # (Xd_0__inst_inst_first_level_2__9__q  & ((Xd_0__inst_inst_first_level_0__9__q ) # 
// (Xd_0__inst_inst_first_level_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__9__q ),
	.datac(!Xd_0__inst_inst_first_level_1__9__q ),
	.datad(!Xd_0__inst_inst_first_level_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_37 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__9__q  $ (!Xd_0__inst_inst_first_level_3__9__q  $ (Xd_0__inst_inst_first_level_5__9__q )) ) + ( Xd_0__inst_inst_inst_add_3_35  ) + ( Xd_0__inst_inst_inst_add_3_34  ))
// Xd_0__inst_inst_inst_add_3_38  = CARRY(( !Xd_0__inst_inst_first_level_4__9__q  $ (!Xd_0__inst_inst_first_level_3__9__q  $ (Xd_0__inst_inst_first_level_5__9__q )) ) + ( Xd_0__inst_inst_inst_add_3_35  ) + ( Xd_0__inst_inst_inst_add_3_34  ))
// Xd_0__inst_inst_inst_add_3_39  = SHARE((!Xd_0__inst_inst_first_level_4__9__q  & (Xd_0__inst_inst_first_level_3__9__q  & Xd_0__inst_inst_first_level_5__9__q )) # (Xd_0__inst_inst_first_level_4__9__q  & ((Xd_0__inst_inst_first_level_5__9__q ) # 
// (Xd_0__inst_inst_first_level_3__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__9__q ),
	.datac(!Xd_0__inst_inst_first_level_3__9__q ),
	.datad(!Xd_0__inst_inst_first_level_5__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_34 ),
	.sharein(Xd_0__inst_inst_inst_add_3_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_37_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_38 ),
	.shareout(Xd_0__inst_inst_inst_add_3_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_42  = CARRY(( !Xd_0__inst_inst_first_level_2__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q  $ (Xd_0__inst_inst_first_level_0__10__q )) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_43  = SHARE((!Xd_0__inst_inst_first_level_2__10__q  & (Xd_0__inst_inst_first_level_1__10__q  & Xd_0__inst_inst_first_level_0__10__q )) # (Xd_0__inst_inst_first_level_2__10__q  & ((Xd_0__inst_inst_first_level_0__10__q ) # 
// (Xd_0__inst_inst_first_level_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__10__q ),
	.datac(!Xd_0__inst_inst_first_level_1__10__q ),
	.datad(!Xd_0__inst_inst_first_level_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_41 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__10__q  $ (!Xd_0__inst_inst_first_level_3__10__q  $ (Xd_0__inst_inst_first_level_5__10__q )) ) + ( Xd_0__inst_inst_inst_add_3_39  ) + ( Xd_0__inst_inst_inst_add_3_38  ))
// Xd_0__inst_inst_inst_add_3_42  = CARRY(( !Xd_0__inst_inst_first_level_4__10__q  $ (!Xd_0__inst_inst_first_level_3__10__q  $ (Xd_0__inst_inst_first_level_5__10__q )) ) + ( Xd_0__inst_inst_inst_add_3_39  ) + ( Xd_0__inst_inst_inst_add_3_38  ))
// Xd_0__inst_inst_inst_add_3_43  = SHARE((!Xd_0__inst_inst_first_level_4__10__q  & (Xd_0__inst_inst_first_level_3__10__q  & Xd_0__inst_inst_first_level_5__10__q )) # (Xd_0__inst_inst_first_level_4__10__q  & ((Xd_0__inst_inst_first_level_5__10__q ) # 
// (Xd_0__inst_inst_first_level_3__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__10__q ),
	.datac(!Xd_0__inst_inst_first_level_3__10__q ),
	.datad(!Xd_0__inst_inst_first_level_5__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_38 ),
	.sharein(Xd_0__inst_inst_inst_add_3_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_42 ),
	.shareout(Xd_0__inst_inst_inst_add_3_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_46  = CARRY(( !Xd_0__inst_inst_first_level_2__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q  $ (Xd_0__inst_inst_first_level_0__11__q )) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_47  = SHARE((!Xd_0__inst_inst_first_level_2__11__q  & (Xd_0__inst_inst_first_level_1__11__q  & Xd_0__inst_inst_first_level_0__11__q )) # (Xd_0__inst_inst_first_level_2__11__q  & ((Xd_0__inst_inst_first_level_0__11__q ) # 
// (Xd_0__inst_inst_first_level_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__11__q ),
	.datac(!Xd_0__inst_inst_first_level_1__11__q ),
	.datad(!Xd_0__inst_inst_first_level_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_45 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__11__q  $ (!Xd_0__inst_inst_first_level_3__11__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_43  ) + ( Xd_0__inst_inst_inst_add_3_42  ))
// Xd_0__inst_inst_inst_add_3_46  = CARRY(( !Xd_0__inst_inst_first_level_4__11__q  $ (!Xd_0__inst_inst_first_level_3__11__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_43  ) + ( Xd_0__inst_inst_inst_add_3_42  ))
// Xd_0__inst_inst_inst_add_3_47  = SHARE((!Xd_0__inst_inst_first_level_4__11__q  & (Xd_0__inst_inst_first_level_3__11__q  & Xd_0__inst_inst_first_level_5__13__q )) # (Xd_0__inst_inst_first_level_4__11__q  & ((Xd_0__inst_inst_first_level_5__13__q ) # 
// (Xd_0__inst_inst_first_level_3__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__11__q ),
	.datac(!Xd_0__inst_inst_first_level_3__11__q ),
	.datad(!Xd_0__inst_inst_first_level_5__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_42 ),
	.sharein(Xd_0__inst_inst_inst_add_3_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_45_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_46 ),
	.shareout(Xd_0__inst_inst_inst_add_3_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_50  = CARRY(( !Xd_0__inst_inst_first_level_2__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q  $ (Xd_0__inst_inst_first_level_0__12__q )) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_51  = SHARE((!Xd_0__inst_inst_first_level_2__12__q  & (Xd_0__inst_inst_first_level_1__12__q  & Xd_0__inst_inst_first_level_0__12__q )) # (Xd_0__inst_inst_first_level_2__12__q  & ((Xd_0__inst_inst_first_level_0__12__q ) # 
// (Xd_0__inst_inst_first_level_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__12__q ),
	.datac(!Xd_0__inst_inst_first_level_1__12__q ),
	.datad(!Xd_0__inst_inst_first_level_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_49 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__12__q  $ (!Xd_0__inst_inst_first_level_3__12__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_47  ) + ( Xd_0__inst_inst_inst_add_3_46  ))
// Xd_0__inst_inst_inst_add_3_50  = CARRY(( !Xd_0__inst_inst_first_level_4__12__q  $ (!Xd_0__inst_inst_first_level_3__12__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_47  ) + ( Xd_0__inst_inst_inst_add_3_46  ))
// Xd_0__inst_inst_inst_add_3_51  = SHARE((!Xd_0__inst_inst_first_level_4__12__q  & (Xd_0__inst_inst_first_level_3__12__q  & Xd_0__inst_inst_first_level_5__13__q )) # (Xd_0__inst_inst_first_level_4__12__q  & ((Xd_0__inst_inst_first_level_5__13__q ) # 
// (Xd_0__inst_inst_first_level_3__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__12__q ),
	.datac(!Xd_0__inst_inst_first_level_3__12__q ),
	.datad(!Xd_0__inst_inst_first_level_5__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_46 ),
	.sharein(Xd_0__inst_inst_inst_add_3_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_49_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_50 ),
	.shareout(Xd_0__inst_inst_inst_add_3_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_54  = CARRY(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_55  = SHARE((!Xd_0__inst_inst_first_level_2__13__q  & (Xd_0__inst_inst_first_level_1__13__q  & Xd_0__inst_inst_first_level_0__13__q )) # (Xd_0__inst_inst_first_level_2__13__q  & ((Xd_0__inst_inst_first_level_0__13__q ) # 
// (Xd_0__inst_inst_first_level_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__13__q ),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_53 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_51  ) + ( Xd_0__inst_inst_inst_add_3_50  ))
// Xd_0__inst_inst_inst_add_3_54  = CARRY(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_51  ) + ( Xd_0__inst_inst_inst_add_3_50  ))
// Xd_0__inst_inst_inst_add_3_55  = SHARE((!Xd_0__inst_inst_first_level_4__13__q  & (Xd_0__inst_inst_first_level_3__13__q  & Xd_0__inst_inst_first_level_5__13__q )) # (Xd_0__inst_inst_first_level_4__13__q  & ((Xd_0__inst_inst_first_level_5__13__q ) # 
// (Xd_0__inst_inst_first_level_3__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__13__q ),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_5__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_50 ),
	.sharein(Xd_0__inst_inst_inst_add_3_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_53_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_54 ),
	.shareout(Xd_0__inst_inst_inst_add_3_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_58  = CARRY(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_59  = SHARE((!Xd_0__inst_inst_first_level_2__13__q  & (Xd_0__inst_inst_first_level_1__13__q  & Xd_0__inst_inst_first_level_0__13__q )) # (Xd_0__inst_inst_first_level_2__13__q  & ((Xd_0__inst_inst_first_level_0__13__q ) # 
// (Xd_0__inst_inst_first_level_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__13__q ),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_57 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_55  ) + ( Xd_0__inst_inst_inst_add_3_54  ))
// Xd_0__inst_inst_inst_add_3_58  = CARRY(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_55  ) + ( Xd_0__inst_inst_inst_add_3_54  ))
// Xd_0__inst_inst_inst_add_3_59  = SHARE((!Xd_0__inst_inst_first_level_4__13__q  & (Xd_0__inst_inst_first_level_3__13__q  & Xd_0__inst_inst_first_level_5__13__q )) # (Xd_0__inst_inst_first_level_4__13__q  & ((Xd_0__inst_inst_first_level_5__13__q ) # 
// (Xd_0__inst_inst_first_level_3__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__13__q ),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_5__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_54 ),
	.sharein(Xd_0__inst_inst_inst_add_3_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_57_sumout ),
	.cout(Xd_0__inst_inst_inst_add_3_58 ),
	.shareout(Xd_0__inst_inst_inst_add_3_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_2__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q  $ (Xd_0__inst_inst_first_level_0__13__q )) ) + ( Xd_0__inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_add_0_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_2__13__q ),
	.datac(!Xd_0__inst_inst_first_level_1__13__q ),
	.datad(!Xd_0__inst_inst_first_level_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_3_61 (
// Equation(s):
// Xd_0__inst_inst_inst_add_3_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_4__13__q  $ (!Xd_0__inst_inst_first_level_3__13__q  $ (Xd_0__inst_inst_first_level_5__13__q )) ) + ( Xd_0__inst_inst_inst_add_3_59  ) + ( Xd_0__inst_inst_inst_add_3_58  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_inst_first_level_4__13__q ),
	.datac(!Xd_0__inst_inst_first_level_3__13__q ),
	.datad(!Xd_0__inst_inst_first_level_5__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_3_58 ),
	.sharein(Xd_0__inst_inst_inst_add_3_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_3_61_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_35 (
// Equation(s):
// Xd_0__inst_mult_20_36  = SUM(( GND ) + ( Xd_0__inst_mult_20_42  ) + ( Xd_0__inst_mult_20_41  ))
// Xd_0__inst_mult_20_37  = CARRY(( GND ) + ( Xd_0__inst_mult_20_42  ) + ( Xd_0__inst_mult_20_41  ))
// Xd_0__inst_mult_20_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_41 ),
	.sharein(Xd_0__inst_mult_20_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_36 ),
	.cout(Xd_0__inst_mult_20_37 ),
	.shareout(Xd_0__inst_mult_20_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_35 (
// Equation(s):
// Xd_0__inst_mult_23_36  = SUM(( GND ) + ( Xd_0__inst_mult_23_42  ) + ( Xd_0__inst_mult_23_41  ))
// Xd_0__inst_mult_23_37  = CARRY(( GND ) + ( Xd_0__inst_mult_23_42  ) + ( Xd_0__inst_mult_23_41  ))
// Xd_0__inst_mult_23_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_41 ),
	.sharein(Xd_0__inst_mult_23_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_36 ),
	.cout(Xd_0__inst_mult_23_37 ),
	.shareout(Xd_0__inst_mult_23_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_16 (
// Equation(s):
// Xd_0__inst_mult_24_44  = CARRY(( GND ) + ( Xd_0__inst_i17_3  ) + ( Xd_0__inst_i17_2  ))
// Xd_0__inst_mult_24_45  = SHARE((din_b[147] & din_a[145]))

	.dataa(!din_b[147]),
	.datab(!din_a[145]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_2 ),
	.sharein(Xd_0__inst_i17_3 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_44 ),
	.shareout(Xd_0__inst_mult_24_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_1 (
// Equation(s):
// Xd_0__inst_inst_add_4_1_sumout  = SUM(( !Xd_0__inst_r_sum1_8__0__q  $ (!Xd_0__inst_r_sum1_7__0__q  $ (Xd_0__inst_r_sum1_6__0__q )) ) + ( Xd_0__inst_mult_26_38  ) + ( Xd_0__inst_mult_26_37  ))
// Xd_0__inst_inst_add_4_2  = CARRY(( !Xd_0__inst_r_sum1_8__0__q  $ (!Xd_0__inst_r_sum1_7__0__q  $ (Xd_0__inst_r_sum1_6__0__q )) ) + ( Xd_0__inst_mult_26_38  ) + ( Xd_0__inst_mult_26_37  ))
// Xd_0__inst_inst_add_4_3  = SHARE((!Xd_0__inst_r_sum1_8__0__q  & (Xd_0__inst_r_sum1_7__0__q  & Xd_0__inst_r_sum1_6__0__q )) # (Xd_0__inst_r_sum1_8__0__q  & ((Xd_0__inst_r_sum1_6__0__q ) # (Xd_0__inst_r_sum1_7__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__0__q ),
	.datac(!Xd_0__inst_r_sum1_7__0__q ),
	.datad(!Xd_0__inst_r_sum1_6__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_37 ),
	.sharein(Xd_0__inst_mult_26_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_1_sumout ),
	.cout(Xd_0__inst_inst_add_4_2 ),
	.shareout(Xd_0__inst_inst_add_4_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_1 (
// Equation(s):
// Xd_0__inst_inst_add_2_1_sumout  = SUM(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_mult_28_38  ) + ( Xd_0__inst_mult_28_37  ))
// Xd_0__inst_inst_add_2_2  = CARRY(( !Xd_0__inst_r_sum1_5__0__q  $ (!Xd_0__inst_r_sum1_4__0__q  $ (Xd_0__inst_r_sum1_3__0__q )) ) + ( Xd_0__inst_mult_28_38  ) + ( Xd_0__inst_mult_28_37  ))
// Xd_0__inst_inst_add_2_3  = SHARE((!Xd_0__inst_r_sum1_5__0__q  & (Xd_0__inst_r_sum1_4__0__q  & Xd_0__inst_r_sum1_3__0__q )) # (Xd_0__inst_r_sum1_5__0__q  & ((Xd_0__inst_r_sum1_3__0__q ) # (Xd_0__inst_r_sum1_4__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__0__q ),
	.datac(!Xd_0__inst_r_sum1_4__0__q ),
	.datad(!Xd_0__inst_r_sum1_3__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_37 ),
	.sharein(Xd_0__inst_mult_28_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_1_sumout ),
	.cout(Xd_0__inst_inst_add_2_2 ),
	.shareout(Xd_0__inst_inst_add_2_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_30_38  ) + ( Xd_0__inst_mult_30_37  ))
// Xd_0__inst_inst_add_0_2  = CARRY(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_30_38  ) + ( Xd_0__inst_mult_30_37  ))
// Xd_0__inst_inst_add_0_3  = SHARE((!Xd_0__inst_r_sum1_2__0__q  & (Xd_0__inst_r_sum1_1__0__q  & Xd_0__inst_r_sum1_0__0__q )) # (Xd_0__inst_r_sum1_2__0__q  & ((Xd_0__inst_r_sum1_0__0__q ) # (Xd_0__inst_r_sum1_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__0__q ),
	.datac(!Xd_0__inst_r_sum1_1__0__q ),
	.datad(!Xd_0__inst_r_sum1_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_37 ),
	.sharein(Xd_0__inst_mult_30_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20 (
// Equation(s):
// Xd_0__inst_mult_20_40  = SUM(( (!din_a[124] & (((din_a[123] & din_b[121])))) # (din_a[124] & (!din_b[120] $ (((!din_a[123]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_20_45  ) + ( Xd_0__inst_mult_20_44  ))
// Xd_0__inst_mult_20_41  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[121])))) # (din_a[124] & (!din_b[120] $ (((!din_a[123]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_20_45  ) + ( Xd_0__inst_mult_20_44  ))
// Xd_0__inst_mult_20_42  = SHARE((din_a[124] & (din_b[120] & (din_a[123] & din_b[121]))))

	.dataa(!din_a[124]),
	.datab(!din_b[120]),
	.datac(!din_a[123]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_44 ),
	.sharein(Xd_0__inst_mult_20_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_40 ),
	.cout(Xd_0__inst_mult_20_41 ),
	.shareout(Xd_0__inst_mult_20_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_1 (
// Equation(s):
// Xd_0__inst_inst_add_8_1_sumout  = SUM(( !Xd_0__inst_r_sum1_14__0__q  $ (!Xd_0__inst_r_sum1_13__0__q  $ (Xd_0__inst_r_sum1_12__0__q )) ) + ( Xd_0__inst_mult_22_38  ) + ( Xd_0__inst_mult_22_37  ))
// Xd_0__inst_inst_add_8_2  = CARRY(( !Xd_0__inst_r_sum1_14__0__q  $ (!Xd_0__inst_r_sum1_13__0__q  $ (Xd_0__inst_r_sum1_12__0__q )) ) + ( Xd_0__inst_mult_22_38  ) + ( Xd_0__inst_mult_22_37  ))
// Xd_0__inst_inst_add_8_3  = SHARE((!Xd_0__inst_r_sum1_14__0__q  & (Xd_0__inst_r_sum1_13__0__q  & Xd_0__inst_r_sum1_12__0__q )) # (Xd_0__inst_r_sum1_14__0__q  & ((Xd_0__inst_r_sum1_12__0__q ) # (Xd_0__inst_r_sum1_13__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__0__q ),
	.datac(!Xd_0__inst_r_sum1_13__0__q ),
	.datad(!Xd_0__inst_r_sum1_12__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_37 ),
	.sharein(Xd_0__inst_mult_22_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_1_sumout ),
	.cout(Xd_0__inst_inst_add_8_2 ),
	.shareout(Xd_0__inst_inst_add_8_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_1 (
// Equation(s):
// Xd_0__inst_inst_add_6_1_sumout  = SUM(( !Xd_0__inst_r_sum1_11__0__q  $ (!Xd_0__inst_r_sum1_10__0__q  $ (Xd_0__inst_r_sum1_9__0__q )) ) + ( Xd_0__inst_mult_19_38  ) + ( Xd_0__inst_mult_19_37  ))
// Xd_0__inst_inst_add_6_2  = CARRY(( !Xd_0__inst_r_sum1_11__0__q  $ (!Xd_0__inst_r_sum1_10__0__q  $ (Xd_0__inst_r_sum1_9__0__q )) ) + ( Xd_0__inst_mult_19_38  ) + ( Xd_0__inst_mult_19_37  ))
// Xd_0__inst_inst_add_6_3  = SHARE((!Xd_0__inst_r_sum1_11__0__q  & (Xd_0__inst_r_sum1_10__0__q  & Xd_0__inst_r_sum1_9__0__q )) # (Xd_0__inst_r_sum1_11__0__q  & ((Xd_0__inst_r_sum1_9__0__q ) # (Xd_0__inst_r_sum1_10__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__0__q ),
	.datac(!Xd_0__inst_r_sum1_10__0__q ),
	.datad(!Xd_0__inst_r_sum1_9__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_37 ),
	.sharein(Xd_0__inst_mult_19_38 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_1_sumout ),
	.cout(Xd_0__inst_inst_add_6_2 ),
	.shareout(Xd_0__inst_inst_add_6_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23 (
// Equation(s):
// Xd_0__inst_mult_23_40  = SUM(( (!din_a[142] & (((din_a[141] & din_b[139])))) # (din_a[142] & (!din_b[138] $ (((!din_a[141]) # (!din_b[139]))))) ) + ( Xd_0__inst_mult_23_45  ) + ( Xd_0__inst_mult_23_44  ))
// Xd_0__inst_mult_23_41  = CARRY(( (!din_a[142] & (((din_a[141] & din_b[139])))) # (din_a[142] & (!din_b[138] $ (((!din_a[141]) # (!din_b[139]))))) ) + ( Xd_0__inst_mult_23_45  ) + ( Xd_0__inst_mult_23_44  ))
// Xd_0__inst_mult_23_42  = SHARE((din_a[142] & (din_b[138] & (din_a[141] & din_b[139]))))

	.dataa(!din_a[142]),
	.datab(!din_b[138]),
	.datac(!din_a[141]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_44 ),
	.sharein(Xd_0__inst_mult_23_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_40 ),
	.cout(Xd_0__inst_mult_23_41 ),
	.shareout(Xd_0__inst_mult_23_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_1 (
// Equation(s):
// Xd_0__inst_i17_1_sumout  = SUM(( !din_a[71] $ (!din_b[71]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_2  = CARRY(( !din_a[71] $ (!din_b[71]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_3  = SHARE(GND)

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_1_sumout ),
	.cout(Xd_0__inst_i17_2 ),
	.shareout(Xd_0__inst_i17_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_5 (
// Equation(s):
// Xd_0__inst_inst_add_4_5_sumout  = SUM(( !Xd_0__inst_r_sum1_8__1__q  $ (!Xd_0__inst_r_sum1_7__1__q  $ (Xd_0__inst_r_sum1_6__1__q )) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_6  = CARRY(( !Xd_0__inst_r_sum1_8__1__q  $ (!Xd_0__inst_r_sum1_7__1__q  $ (Xd_0__inst_r_sum1_6__1__q )) ) + ( Xd_0__inst_inst_add_4_3  ) + ( Xd_0__inst_inst_add_4_2  ))
// Xd_0__inst_inst_add_4_7  = SHARE((!Xd_0__inst_r_sum1_8__1__q  & (Xd_0__inst_r_sum1_7__1__q  & Xd_0__inst_r_sum1_6__1__q )) # (Xd_0__inst_r_sum1_8__1__q  & ((Xd_0__inst_r_sum1_6__1__q ) # (Xd_0__inst_r_sum1_7__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__1__q ),
	.datac(!Xd_0__inst_r_sum1_7__1__q ),
	.datad(!Xd_0__inst_r_sum1_6__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_2 ),
	.sharein(Xd_0__inst_inst_add_4_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_5_sumout ),
	.cout(Xd_0__inst_inst_add_4_6 ),
	.shareout(Xd_0__inst_inst_add_4_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_5 (
// Equation(s):
// Xd_0__inst_inst_add_2_5_sumout  = SUM(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_6  = CARRY(( !Xd_0__inst_r_sum1_5__1__q  $ (!Xd_0__inst_r_sum1_4__1__q  $ (Xd_0__inst_r_sum1_3__1__q )) ) + ( Xd_0__inst_inst_add_2_3  ) + ( Xd_0__inst_inst_add_2_2  ))
// Xd_0__inst_inst_add_2_7  = SHARE((!Xd_0__inst_r_sum1_5__1__q  & (Xd_0__inst_r_sum1_4__1__q  & Xd_0__inst_r_sum1_3__1__q )) # (Xd_0__inst_r_sum1_5__1__q  & ((Xd_0__inst_r_sum1_3__1__q ) # (Xd_0__inst_r_sum1_4__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__1__q ),
	.datac(!Xd_0__inst_r_sum1_4__1__q ),
	.datad(!Xd_0__inst_r_sum1_3__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_2 ),
	.sharein(Xd_0__inst_inst_add_2_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_5_sumout ),
	.cout(Xd_0__inst_inst_add_2_6 ),
	.shareout(Xd_0__inst_inst_add_2_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_6  = CARRY(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_7  = SHARE((!Xd_0__inst_r_sum1_2__1__q  & (Xd_0__inst_r_sum1_1__1__q  & Xd_0__inst_r_sum1_0__1__q )) # (Xd_0__inst_r_sum1_2__1__q  & ((Xd_0__inst_r_sum1_0__1__q ) # (Xd_0__inst_r_sum1_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__1__q ),
	.datad(!Xd_0__inst_r_sum1_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_5 (
// Equation(s):
// Xd_0__inst_inst_add_8_5_sumout  = SUM(( !Xd_0__inst_r_sum1_14__1__q  $ (!Xd_0__inst_r_sum1_13__1__q  $ (Xd_0__inst_r_sum1_12__1__q )) ) + ( Xd_0__inst_inst_add_8_3  ) + ( Xd_0__inst_inst_add_8_2  ))
// Xd_0__inst_inst_add_8_6  = CARRY(( !Xd_0__inst_r_sum1_14__1__q  $ (!Xd_0__inst_r_sum1_13__1__q  $ (Xd_0__inst_r_sum1_12__1__q )) ) + ( Xd_0__inst_inst_add_8_3  ) + ( Xd_0__inst_inst_add_8_2  ))
// Xd_0__inst_inst_add_8_7  = SHARE((!Xd_0__inst_r_sum1_14__1__q  & (Xd_0__inst_r_sum1_13__1__q  & Xd_0__inst_r_sum1_12__1__q )) # (Xd_0__inst_r_sum1_14__1__q  & ((Xd_0__inst_r_sum1_12__1__q ) # (Xd_0__inst_r_sum1_13__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__1__q ),
	.datac(!Xd_0__inst_r_sum1_13__1__q ),
	.datad(!Xd_0__inst_r_sum1_12__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_2 ),
	.sharein(Xd_0__inst_inst_add_8_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_5_sumout ),
	.cout(Xd_0__inst_inst_add_8_6 ),
	.shareout(Xd_0__inst_inst_add_8_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_5 (
// Equation(s):
// Xd_0__inst_inst_add_6_5_sumout  = SUM(( !Xd_0__inst_r_sum1_11__1__q  $ (!Xd_0__inst_r_sum1_10__1__q  $ (Xd_0__inst_r_sum1_9__1__q )) ) + ( Xd_0__inst_inst_add_6_3  ) + ( Xd_0__inst_inst_add_6_2  ))
// Xd_0__inst_inst_add_6_6  = CARRY(( !Xd_0__inst_r_sum1_11__1__q  $ (!Xd_0__inst_r_sum1_10__1__q  $ (Xd_0__inst_r_sum1_9__1__q )) ) + ( Xd_0__inst_inst_add_6_3  ) + ( Xd_0__inst_inst_add_6_2  ))
// Xd_0__inst_inst_add_6_7  = SHARE((!Xd_0__inst_r_sum1_11__1__q  & (Xd_0__inst_r_sum1_10__1__q  & Xd_0__inst_r_sum1_9__1__q )) # (Xd_0__inst_r_sum1_11__1__q  & ((Xd_0__inst_r_sum1_9__1__q ) # (Xd_0__inst_r_sum1_10__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__1__q ),
	.datac(!Xd_0__inst_r_sum1_10__1__q ),
	.datad(!Xd_0__inst_r_sum1_9__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_2 ),
	.sharein(Xd_0__inst_inst_add_6_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_5_sumout ),
	.cout(Xd_0__inst_inst_add_6_6 ),
	.shareout(Xd_0__inst_inst_add_6_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_9 (
// Equation(s):
// Xd_0__inst_inst_add_4_9_sumout  = SUM(( !Xd_0__inst_r_sum1_8__2__q  $ (!Xd_0__inst_r_sum1_7__2__q  $ (Xd_0__inst_r_sum1_6__2__q )) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_10  = CARRY(( !Xd_0__inst_r_sum1_8__2__q  $ (!Xd_0__inst_r_sum1_7__2__q  $ (Xd_0__inst_r_sum1_6__2__q )) ) + ( Xd_0__inst_inst_add_4_7  ) + ( Xd_0__inst_inst_add_4_6  ))
// Xd_0__inst_inst_add_4_11  = SHARE((!Xd_0__inst_r_sum1_8__2__q  & (Xd_0__inst_r_sum1_7__2__q  & Xd_0__inst_r_sum1_6__2__q )) # (Xd_0__inst_r_sum1_8__2__q  & ((Xd_0__inst_r_sum1_6__2__q ) # (Xd_0__inst_r_sum1_7__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__2__q ),
	.datac(!Xd_0__inst_r_sum1_7__2__q ),
	.datad(!Xd_0__inst_r_sum1_6__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_6 ),
	.sharein(Xd_0__inst_inst_add_4_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_9_sumout ),
	.cout(Xd_0__inst_inst_add_4_10 ),
	.shareout(Xd_0__inst_inst_add_4_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_9 (
// Equation(s):
// Xd_0__inst_inst_add_2_9_sumout  = SUM(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_10  = CARRY(( !Xd_0__inst_r_sum1_5__2__q  $ (!Xd_0__inst_r_sum1_4__2__q  $ (Xd_0__inst_r_sum1_3__2__q )) ) + ( Xd_0__inst_inst_add_2_7  ) + ( Xd_0__inst_inst_add_2_6  ))
// Xd_0__inst_inst_add_2_11  = SHARE((!Xd_0__inst_r_sum1_5__2__q  & (Xd_0__inst_r_sum1_4__2__q  & Xd_0__inst_r_sum1_3__2__q )) # (Xd_0__inst_r_sum1_5__2__q  & ((Xd_0__inst_r_sum1_3__2__q ) # (Xd_0__inst_r_sum1_4__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__2__q ),
	.datac(!Xd_0__inst_r_sum1_4__2__q ),
	.datad(!Xd_0__inst_r_sum1_3__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_6 ),
	.sharein(Xd_0__inst_inst_add_2_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_9_sumout ),
	.cout(Xd_0__inst_inst_add_2_10 ),
	.shareout(Xd_0__inst_inst_add_2_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_10  = CARRY(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_11  = SHARE((!Xd_0__inst_r_sum1_2__2__q  & (Xd_0__inst_r_sum1_1__2__q  & Xd_0__inst_r_sum1_0__2__q )) # (Xd_0__inst_r_sum1_2__2__q  & ((Xd_0__inst_r_sum1_0__2__q ) # (Xd_0__inst_r_sum1_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__2__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_9 (
// Equation(s):
// Xd_0__inst_inst_add_8_9_sumout  = SUM(( !Xd_0__inst_r_sum1_14__2__q  $ (!Xd_0__inst_r_sum1_13__2__q  $ (Xd_0__inst_r_sum1_12__2__q )) ) + ( Xd_0__inst_inst_add_8_7  ) + ( Xd_0__inst_inst_add_8_6  ))
// Xd_0__inst_inst_add_8_10  = CARRY(( !Xd_0__inst_r_sum1_14__2__q  $ (!Xd_0__inst_r_sum1_13__2__q  $ (Xd_0__inst_r_sum1_12__2__q )) ) + ( Xd_0__inst_inst_add_8_7  ) + ( Xd_0__inst_inst_add_8_6  ))
// Xd_0__inst_inst_add_8_11  = SHARE((!Xd_0__inst_r_sum1_14__2__q  & (Xd_0__inst_r_sum1_13__2__q  & Xd_0__inst_r_sum1_12__2__q )) # (Xd_0__inst_r_sum1_14__2__q  & ((Xd_0__inst_r_sum1_12__2__q ) # (Xd_0__inst_r_sum1_13__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__2__q ),
	.datac(!Xd_0__inst_r_sum1_13__2__q ),
	.datad(!Xd_0__inst_r_sum1_12__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_6 ),
	.sharein(Xd_0__inst_inst_add_8_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_9_sumout ),
	.cout(Xd_0__inst_inst_add_8_10 ),
	.shareout(Xd_0__inst_inst_add_8_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_9 (
// Equation(s):
// Xd_0__inst_inst_add_6_9_sumout  = SUM(( !Xd_0__inst_r_sum1_11__2__q  $ (!Xd_0__inst_r_sum1_10__2__q  $ (Xd_0__inst_r_sum1_9__2__q )) ) + ( Xd_0__inst_inst_add_6_7  ) + ( Xd_0__inst_inst_add_6_6  ))
// Xd_0__inst_inst_add_6_10  = CARRY(( !Xd_0__inst_r_sum1_11__2__q  $ (!Xd_0__inst_r_sum1_10__2__q  $ (Xd_0__inst_r_sum1_9__2__q )) ) + ( Xd_0__inst_inst_add_6_7  ) + ( Xd_0__inst_inst_add_6_6  ))
// Xd_0__inst_inst_add_6_11  = SHARE((!Xd_0__inst_r_sum1_11__2__q  & (Xd_0__inst_r_sum1_10__2__q  & Xd_0__inst_r_sum1_9__2__q )) # (Xd_0__inst_r_sum1_11__2__q  & ((Xd_0__inst_r_sum1_9__2__q ) # (Xd_0__inst_r_sum1_10__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__2__q ),
	.datac(!Xd_0__inst_r_sum1_10__2__q ),
	.datad(!Xd_0__inst_r_sum1_9__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_6 ),
	.sharein(Xd_0__inst_inst_add_6_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_9_sumout ),
	.cout(Xd_0__inst_inst_add_6_10 ),
	.shareout(Xd_0__inst_inst_add_6_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_13 (
// Equation(s):
// Xd_0__inst_inst_add_4_13_sumout  = SUM(( !Xd_0__inst_r_sum1_8__3__q  $ (!Xd_0__inst_r_sum1_7__3__q  $ (Xd_0__inst_r_sum1_6__3__q )) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_14  = CARRY(( !Xd_0__inst_r_sum1_8__3__q  $ (!Xd_0__inst_r_sum1_7__3__q  $ (Xd_0__inst_r_sum1_6__3__q )) ) + ( Xd_0__inst_inst_add_4_11  ) + ( Xd_0__inst_inst_add_4_10  ))
// Xd_0__inst_inst_add_4_15  = SHARE((!Xd_0__inst_r_sum1_8__3__q  & (Xd_0__inst_r_sum1_7__3__q  & Xd_0__inst_r_sum1_6__3__q )) # (Xd_0__inst_r_sum1_8__3__q  & ((Xd_0__inst_r_sum1_6__3__q ) # (Xd_0__inst_r_sum1_7__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__3__q ),
	.datac(!Xd_0__inst_r_sum1_7__3__q ),
	.datad(!Xd_0__inst_r_sum1_6__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_10 ),
	.sharein(Xd_0__inst_inst_add_4_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_13_sumout ),
	.cout(Xd_0__inst_inst_add_4_14 ),
	.shareout(Xd_0__inst_inst_add_4_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_13 (
// Equation(s):
// Xd_0__inst_inst_add_2_13_sumout  = SUM(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_14  = CARRY(( !Xd_0__inst_r_sum1_5__3__q  $ (!Xd_0__inst_r_sum1_4__3__q  $ (Xd_0__inst_r_sum1_3__3__q )) ) + ( Xd_0__inst_inst_add_2_11  ) + ( Xd_0__inst_inst_add_2_10  ))
// Xd_0__inst_inst_add_2_15  = SHARE((!Xd_0__inst_r_sum1_5__3__q  & (Xd_0__inst_r_sum1_4__3__q  & Xd_0__inst_r_sum1_3__3__q )) # (Xd_0__inst_r_sum1_5__3__q  & ((Xd_0__inst_r_sum1_3__3__q ) # (Xd_0__inst_r_sum1_4__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__3__q ),
	.datac(!Xd_0__inst_r_sum1_4__3__q ),
	.datad(!Xd_0__inst_r_sum1_3__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_10 ),
	.sharein(Xd_0__inst_inst_add_2_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_13_sumout ),
	.cout(Xd_0__inst_inst_add_2_14 ),
	.shareout(Xd_0__inst_inst_add_2_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_14  = CARRY(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_15  = SHARE((!Xd_0__inst_r_sum1_2__3__q  & (Xd_0__inst_r_sum1_1__3__q  & Xd_0__inst_r_sum1_0__3__q )) # (Xd_0__inst_r_sum1_2__3__q  & ((Xd_0__inst_r_sum1_0__3__q ) # (Xd_0__inst_r_sum1_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__3__q ),
	.datad(!Xd_0__inst_r_sum1_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_13 (
// Equation(s):
// Xd_0__inst_inst_add_8_13_sumout  = SUM(( !Xd_0__inst_r_sum1_14__3__q  $ (!Xd_0__inst_r_sum1_13__3__q  $ (Xd_0__inst_r_sum1_12__3__q )) ) + ( Xd_0__inst_inst_add_8_11  ) + ( Xd_0__inst_inst_add_8_10  ))
// Xd_0__inst_inst_add_8_14  = CARRY(( !Xd_0__inst_r_sum1_14__3__q  $ (!Xd_0__inst_r_sum1_13__3__q  $ (Xd_0__inst_r_sum1_12__3__q )) ) + ( Xd_0__inst_inst_add_8_11  ) + ( Xd_0__inst_inst_add_8_10  ))
// Xd_0__inst_inst_add_8_15  = SHARE((!Xd_0__inst_r_sum1_14__3__q  & (Xd_0__inst_r_sum1_13__3__q  & Xd_0__inst_r_sum1_12__3__q )) # (Xd_0__inst_r_sum1_14__3__q  & ((Xd_0__inst_r_sum1_12__3__q ) # (Xd_0__inst_r_sum1_13__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__3__q ),
	.datac(!Xd_0__inst_r_sum1_13__3__q ),
	.datad(!Xd_0__inst_r_sum1_12__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_10 ),
	.sharein(Xd_0__inst_inst_add_8_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_13_sumout ),
	.cout(Xd_0__inst_inst_add_8_14 ),
	.shareout(Xd_0__inst_inst_add_8_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_13 (
// Equation(s):
// Xd_0__inst_inst_add_6_13_sumout  = SUM(( !Xd_0__inst_r_sum1_11__3__q  $ (!Xd_0__inst_r_sum1_10__3__q  $ (Xd_0__inst_r_sum1_9__3__q )) ) + ( Xd_0__inst_inst_add_6_11  ) + ( Xd_0__inst_inst_add_6_10  ))
// Xd_0__inst_inst_add_6_14  = CARRY(( !Xd_0__inst_r_sum1_11__3__q  $ (!Xd_0__inst_r_sum1_10__3__q  $ (Xd_0__inst_r_sum1_9__3__q )) ) + ( Xd_0__inst_inst_add_6_11  ) + ( Xd_0__inst_inst_add_6_10  ))
// Xd_0__inst_inst_add_6_15  = SHARE((!Xd_0__inst_r_sum1_11__3__q  & (Xd_0__inst_r_sum1_10__3__q  & Xd_0__inst_r_sum1_9__3__q )) # (Xd_0__inst_r_sum1_11__3__q  & ((Xd_0__inst_r_sum1_9__3__q ) # (Xd_0__inst_r_sum1_10__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__3__q ),
	.datac(!Xd_0__inst_r_sum1_10__3__q ),
	.datad(!Xd_0__inst_r_sum1_9__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_10 ),
	.sharein(Xd_0__inst_inst_add_6_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_13_sumout ),
	.cout(Xd_0__inst_inst_add_6_14 ),
	.shareout(Xd_0__inst_inst_add_6_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_17 (
// Equation(s):
// Xd_0__inst_inst_add_4_17_sumout  = SUM(( !Xd_0__inst_r_sum1_8__4__q  $ (!Xd_0__inst_r_sum1_7__4__q  $ (Xd_0__inst_r_sum1_6__4__q )) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_18  = CARRY(( !Xd_0__inst_r_sum1_8__4__q  $ (!Xd_0__inst_r_sum1_7__4__q  $ (Xd_0__inst_r_sum1_6__4__q )) ) + ( Xd_0__inst_inst_add_4_15  ) + ( Xd_0__inst_inst_add_4_14  ))
// Xd_0__inst_inst_add_4_19  = SHARE((!Xd_0__inst_r_sum1_8__4__q  & (Xd_0__inst_r_sum1_7__4__q  & Xd_0__inst_r_sum1_6__4__q )) # (Xd_0__inst_r_sum1_8__4__q  & ((Xd_0__inst_r_sum1_6__4__q ) # (Xd_0__inst_r_sum1_7__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__4__q ),
	.datac(!Xd_0__inst_r_sum1_7__4__q ),
	.datad(!Xd_0__inst_r_sum1_6__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_14 ),
	.sharein(Xd_0__inst_inst_add_4_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_17_sumout ),
	.cout(Xd_0__inst_inst_add_4_18 ),
	.shareout(Xd_0__inst_inst_add_4_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_17 (
// Equation(s):
// Xd_0__inst_inst_add_2_17_sumout  = SUM(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_18  = CARRY(( !Xd_0__inst_r_sum1_5__4__q  $ (!Xd_0__inst_r_sum1_4__4__q  $ (Xd_0__inst_r_sum1_3__4__q )) ) + ( Xd_0__inst_inst_add_2_15  ) + ( Xd_0__inst_inst_add_2_14  ))
// Xd_0__inst_inst_add_2_19  = SHARE((!Xd_0__inst_r_sum1_5__4__q  & (Xd_0__inst_r_sum1_4__4__q  & Xd_0__inst_r_sum1_3__4__q )) # (Xd_0__inst_r_sum1_5__4__q  & ((Xd_0__inst_r_sum1_3__4__q ) # (Xd_0__inst_r_sum1_4__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__4__q ),
	.datac(!Xd_0__inst_r_sum1_4__4__q ),
	.datad(!Xd_0__inst_r_sum1_3__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_14 ),
	.sharein(Xd_0__inst_inst_add_2_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_17_sumout ),
	.cout(Xd_0__inst_inst_add_2_18 ),
	.shareout(Xd_0__inst_inst_add_2_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_18  = CARRY(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_19  = SHARE((!Xd_0__inst_r_sum1_2__4__q  & (Xd_0__inst_r_sum1_1__4__q  & Xd_0__inst_r_sum1_0__4__q )) # (Xd_0__inst_r_sum1_2__4__q  & ((Xd_0__inst_r_sum1_0__4__q ) # (Xd_0__inst_r_sum1_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__4__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_17 (
// Equation(s):
// Xd_0__inst_inst_add_8_17_sumout  = SUM(( !Xd_0__inst_r_sum1_14__4__q  $ (!Xd_0__inst_r_sum1_13__4__q  $ (Xd_0__inst_r_sum1_12__4__q )) ) + ( Xd_0__inst_inst_add_8_15  ) + ( Xd_0__inst_inst_add_8_14  ))
// Xd_0__inst_inst_add_8_18  = CARRY(( !Xd_0__inst_r_sum1_14__4__q  $ (!Xd_0__inst_r_sum1_13__4__q  $ (Xd_0__inst_r_sum1_12__4__q )) ) + ( Xd_0__inst_inst_add_8_15  ) + ( Xd_0__inst_inst_add_8_14  ))
// Xd_0__inst_inst_add_8_19  = SHARE((!Xd_0__inst_r_sum1_14__4__q  & (Xd_0__inst_r_sum1_13__4__q  & Xd_0__inst_r_sum1_12__4__q )) # (Xd_0__inst_r_sum1_14__4__q  & ((Xd_0__inst_r_sum1_12__4__q ) # (Xd_0__inst_r_sum1_13__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__4__q ),
	.datac(!Xd_0__inst_r_sum1_13__4__q ),
	.datad(!Xd_0__inst_r_sum1_12__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_14 ),
	.sharein(Xd_0__inst_inst_add_8_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_17_sumout ),
	.cout(Xd_0__inst_inst_add_8_18 ),
	.shareout(Xd_0__inst_inst_add_8_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_17 (
// Equation(s):
// Xd_0__inst_inst_add_6_17_sumout  = SUM(( !Xd_0__inst_r_sum1_11__4__q  $ (!Xd_0__inst_r_sum1_10__4__q  $ (Xd_0__inst_r_sum1_9__4__q )) ) + ( Xd_0__inst_inst_add_6_15  ) + ( Xd_0__inst_inst_add_6_14  ))
// Xd_0__inst_inst_add_6_18  = CARRY(( !Xd_0__inst_r_sum1_11__4__q  $ (!Xd_0__inst_r_sum1_10__4__q  $ (Xd_0__inst_r_sum1_9__4__q )) ) + ( Xd_0__inst_inst_add_6_15  ) + ( Xd_0__inst_inst_add_6_14  ))
// Xd_0__inst_inst_add_6_19  = SHARE((!Xd_0__inst_r_sum1_11__4__q  & (Xd_0__inst_r_sum1_10__4__q  & Xd_0__inst_r_sum1_9__4__q )) # (Xd_0__inst_r_sum1_11__4__q  & ((Xd_0__inst_r_sum1_9__4__q ) # (Xd_0__inst_r_sum1_10__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__4__q ),
	.datac(!Xd_0__inst_r_sum1_10__4__q ),
	.datad(!Xd_0__inst_r_sum1_9__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_14 ),
	.sharein(Xd_0__inst_inst_add_6_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_17_sumout ),
	.cout(Xd_0__inst_inst_add_6_18 ),
	.shareout(Xd_0__inst_inst_add_6_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_21 (
// Equation(s):
// Xd_0__inst_inst_add_4_21_sumout  = SUM(( !Xd_0__inst_r_sum1_8__5__q  $ (!Xd_0__inst_r_sum1_7__5__q  $ (Xd_0__inst_r_sum1_6__5__q )) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_22  = CARRY(( !Xd_0__inst_r_sum1_8__5__q  $ (!Xd_0__inst_r_sum1_7__5__q  $ (Xd_0__inst_r_sum1_6__5__q )) ) + ( Xd_0__inst_inst_add_4_19  ) + ( Xd_0__inst_inst_add_4_18  ))
// Xd_0__inst_inst_add_4_23  = SHARE((!Xd_0__inst_r_sum1_8__5__q  & (Xd_0__inst_r_sum1_7__5__q  & Xd_0__inst_r_sum1_6__5__q )) # (Xd_0__inst_r_sum1_8__5__q  & ((Xd_0__inst_r_sum1_6__5__q ) # (Xd_0__inst_r_sum1_7__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__5__q ),
	.datac(!Xd_0__inst_r_sum1_7__5__q ),
	.datad(!Xd_0__inst_r_sum1_6__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_18 ),
	.sharein(Xd_0__inst_inst_add_4_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_21_sumout ),
	.cout(Xd_0__inst_inst_add_4_22 ),
	.shareout(Xd_0__inst_inst_add_4_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_21 (
// Equation(s):
// Xd_0__inst_inst_add_2_21_sumout  = SUM(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_22  = CARRY(( !Xd_0__inst_r_sum1_5__5__q  $ (!Xd_0__inst_r_sum1_4__5__q  $ (Xd_0__inst_r_sum1_3__5__q )) ) + ( Xd_0__inst_inst_add_2_19  ) + ( Xd_0__inst_inst_add_2_18  ))
// Xd_0__inst_inst_add_2_23  = SHARE((!Xd_0__inst_r_sum1_5__5__q  & (Xd_0__inst_r_sum1_4__5__q  & Xd_0__inst_r_sum1_3__5__q )) # (Xd_0__inst_r_sum1_5__5__q  & ((Xd_0__inst_r_sum1_3__5__q ) # (Xd_0__inst_r_sum1_4__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__5__q ),
	.datac(!Xd_0__inst_r_sum1_4__5__q ),
	.datad(!Xd_0__inst_r_sum1_3__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_18 ),
	.sharein(Xd_0__inst_inst_add_2_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_21_sumout ),
	.cout(Xd_0__inst_inst_add_2_22 ),
	.shareout(Xd_0__inst_inst_add_2_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_22  = CARRY(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_23  = SHARE((!Xd_0__inst_r_sum1_2__5__q  & (Xd_0__inst_r_sum1_1__5__q  & Xd_0__inst_r_sum1_0__5__q )) # (Xd_0__inst_r_sum1_2__5__q  & ((Xd_0__inst_r_sum1_0__5__q ) # (Xd_0__inst_r_sum1_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__5__q ),
	.datad(!Xd_0__inst_r_sum1_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_21 (
// Equation(s):
// Xd_0__inst_inst_add_8_21_sumout  = SUM(( !Xd_0__inst_r_sum1_14__5__q  $ (!Xd_0__inst_r_sum1_13__5__q  $ (Xd_0__inst_r_sum1_12__5__q )) ) + ( Xd_0__inst_inst_add_8_19  ) + ( Xd_0__inst_inst_add_8_18  ))
// Xd_0__inst_inst_add_8_22  = CARRY(( !Xd_0__inst_r_sum1_14__5__q  $ (!Xd_0__inst_r_sum1_13__5__q  $ (Xd_0__inst_r_sum1_12__5__q )) ) + ( Xd_0__inst_inst_add_8_19  ) + ( Xd_0__inst_inst_add_8_18  ))
// Xd_0__inst_inst_add_8_23  = SHARE((!Xd_0__inst_r_sum1_14__5__q  & (Xd_0__inst_r_sum1_13__5__q  & Xd_0__inst_r_sum1_12__5__q )) # (Xd_0__inst_r_sum1_14__5__q  & ((Xd_0__inst_r_sum1_12__5__q ) # (Xd_0__inst_r_sum1_13__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__5__q ),
	.datac(!Xd_0__inst_r_sum1_13__5__q ),
	.datad(!Xd_0__inst_r_sum1_12__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_18 ),
	.sharein(Xd_0__inst_inst_add_8_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_21_sumout ),
	.cout(Xd_0__inst_inst_add_8_22 ),
	.shareout(Xd_0__inst_inst_add_8_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_21 (
// Equation(s):
// Xd_0__inst_inst_add_6_21_sumout  = SUM(( !Xd_0__inst_r_sum1_11__5__q  $ (!Xd_0__inst_r_sum1_10__5__q  $ (Xd_0__inst_r_sum1_9__5__q )) ) + ( Xd_0__inst_inst_add_6_19  ) + ( Xd_0__inst_inst_add_6_18  ))
// Xd_0__inst_inst_add_6_22  = CARRY(( !Xd_0__inst_r_sum1_11__5__q  $ (!Xd_0__inst_r_sum1_10__5__q  $ (Xd_0__inst_r_sum1_9__5__q )) ) + ( Xd_0__inst_inst_add_6_19  ) + ( Xd_0__inst_inst_add_6_18  ))
// Xd_0__inst_inst_add_6_23  = SHARE((!Xd_0__inst_r_sum1_11__5__q  & (Xd_0__inst_r_sum1_10__5__q  & Xd_0__inst_r_sum1_9__5__q )) # (Xd_0__inst_r_sum1_11__5__q  & ((Xd_0__inst_r_sum1_9__5__q ) # (Xd_0__inst_r_sum1_10__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__5__q ),
	.datac(!Xd_0__inst_r_sum1_10__5__q ),
	.datad(!Xd_0__inst_r_sum1_9__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_18 ),
	.sharein(Xd_0__inst_inst_add_6_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_21_sumout ),
	.cout(Xd_0__inst_inst_add_6_22 ),
	.shareout(Xd_0__inst_inst_add_6_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_25 (
// Equation(s):
// Xd_0__inst_inst_add_4_25_sumout  = SUM(( !Xd_0__inst_r_sum1_8__6__q  $ (!Xd_0__inst_r_sum1_7__6__q  $ (Xd_0__inst_r_sum1_6__6__q )) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_26  = CARRY(( !Xd_0__inst_r_sum1_8__6__q  $ (!Xd_0__inst_r_sum1_7__6__q  $ (Xd_0__inst_r_sum1_6__6__q )) ) + ( Xd_0__inst_inst_add_4_23  ) + ( Xd_0__inst_inst_add_4_22  ))
// Xd_0__inst_inst_add_4_27  = SHARE((!Xd_0__inst_r_sum1_8__6__q  & (Xd_0__inst_r_sum1_7__6__q  & Xd_0__inst_r_sum1_6__6__q )) # (Xd_0__inst_r_sum1_8__6__q  & ((Xd_0__inst_r_sum1_6__6__q ) # (Xd_0__inst_r_sum1_7__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__6__q ),
	.datac(!Xd_0__inst_r_sum1_7__6__q ),
	.datad(!Xd_0__inst_r_sum1_6__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_22 ),
	.sharein(Xd_0__inst_inst_add_4_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_25_sumout ),
	.cout(Xd_0__inst_inst_add_4_26 ),
	.shareout(Xd_0__inst_inst_add_4_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_25 (
// Equation(s):
// Xd_0__inst_inst_add_2_25_sumout  = SUM(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_26  = CARRY(( !Xd_0__inst_r_sum1_5__6__q  $ (!Xd_0__inst_r_sum1_4__6__q  $ (Xd_0__inst_r_sum1_3__6__q )) ) + ( Xd_0__inst_inst_add_2_23  ) + ( Xd_0__inst_inst_add_2_22  ))
// Xd_0__inst_inst_add_2_27  = SHARE((!Xd_0__inst_r_sum1_5__6__q  & (Xd_0__inst_r_sum1_4__6__q  & Xd_0__inst_r_sum1_3__6__q )) # (Xd_0__inst_r_sum1_5__6__q  & ((Xd_0__inst_r_sum1_3__6__q ) # (Xd_0__inst_r_sum1_4__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__6__q ),
	.datac(!Xd_0__inst_r_sum1_4__6__q ),
	.datad(!Xd_0__inst_r_sum1_3__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_22 ),
	.sharein(Xd_0__inst_inst_add_2_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_25_sumout ),
	.cout(Xd_0__inst_inst_add_2_26 ),
	.shareout(Xd_0__inst_inst_add_2_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_26  = CARRY(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_27  = SHARE((!Xd_0__inst_r_sum1_2__6__q  & (Xd_0__inst_r_sum1_1__6__q  & Xd_0__inst_r_sum1_0__6__q )) # (Xd_0__inst_r_sum1_2__6__q  & ((Xd_0__inst_r_sum1_0__6__q ) # (Xd_0__inst_r_sum1_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__6__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_25 (
// Equation(s):
// Xd_0__inst_inst_add_8_25_sumout  = SUM(( !Xd_0__inst_r_sum1_14__6__q  $ (!Xd_0__inst_r_sum1_13__6__q  $ (Xd_0__inst_r_sum1_12__6__q )) ) + ( Xd_0__inst_inst_add_8_23  ) + ( Xd_0__inst_inst_add_8_22  ))
// Xd_0__inst_inst_add_8_26  = CARRY(( !Xd_0__inst_r_sum1_14__6__q  $ (!Xd_0__inst_r_sum1_13__6__q  $ (Xd_0__inst_r_sum1_12__6__q )) ) + ( Xd_0__inst_inst_add_8_23  ) + ( Xd_0__inst_inst_add_8_22  ))
// Xd_0__inst_inst_add_8_27  = SHARE((!Xd_0__inst_r_sum1_14__6__q  & (Xd_0__inst_r_sum1_13__6__q  & Xd_0__inst_r_sum1_12__6__q )) # (Xd_0__inst_r_sum1_14__6__q  & ((Xd_0__inst_r_sum1_12__6__q ) # (Xd_0__inst_r_sum1_13__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__6__q ),
	.datac(!Xd_0__inst_r_sum1_13__6__q ),
	.datad(!Xd_0__inst_r_sum1_12__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_22 ),
	.sharein(Xd_0__inst_inst_add_8_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_25_sumout ),
	.cout(Xd_0__inst_inst_add_8_26 ),
	.shareout(Xd_0__inst_inst_add_8_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_25 (
// Equation(s):
// Xd_0__inst_inst_add_6_25_sumout  = SUM(( !Xd_0__inst_r_sum1_11__6__q  $ (!Xd_0__inst_r_sum1_10__6__q  $ (Xd_0__inst_r_sum1_9__6__q )) ) + ( Xd_0__inst_inst_add_6_23  ) + ( Xd_0__inst_inst_add_6_22  ))
// Xd_0__inst_inst_add_6_26  = CARRY(( !Xd_0__inst_r_sum1_11__6__q  $ (!Xd_0__inst_r_sum1_10__6__q  $ (Xd_0__inst_r_sum1_9__6__q )) ) + ( Xd_0__inst_inst_add_6_23  ) + ( Xd_0__inst_inst_add_6_22  ))
// Xd_0__inst_inst_add_6_27  = SHARE((!Xd_0__inst_r_sum1_11__6__q  & (Xd_0__inst_r_sum1_10__6__q  & Xd_0__inst_r_sum1_9__6__q )) # (Xd_0__inst_r_sum1_11__6__q  & ((Xd_0__inst_r_sum1_9__6__q ) # (Xd_0__inst_r_sum1_10__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__6__q ),
	.datac(!Xd_0__inst_r_sum1_10__6__q ),
	.datad(!Xd_0__inst_r_sum1_9__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_22 ),
	.sharein(Xd_0__inst_inst_add_6_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_25_sumout ),
	.cout(Xd_0__inst_inst_add_6_26 ),
	.shareout(Xd_0__inst_inst_add_6_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_29 (
// Equation(s):
// Xd_0__inst_inst_add_4_29_sumout  = SUM(( !Xd_0__inst_r_sum1_8__7__q  $ (!Xd_0__inst_r_sum1_7__7__q  $ (Xd_0__inst_r_sum1_6__7__q )) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_30  = CARRY(( !Xd_0__inst_r_sum1_8__7__q  $ (!Xd_0__inst_r_sum1_7__7__q  $ (Xd_0__inst_r_sum1_6__7__q )) ) + ( Xd_0__inst_inst_add_4_27  ) + ( Xd_0__inst_inst_add_4_26  ))
// Xd_0__inst_inst_add_4_31  = SHARE((!Xd_0__inst_r_sum1_8__7__q  & (Xd_0__inst_r_sum1_7__7__q  & Xd_0__inst_r_sum1_6__7__q )) # (Xd_0__inst_r_sum1_8__7__q  & ((Xd_0__inst_r_sum1_6__7__q ) # (Xd_0__inst_r_sum1_7__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__7__q ),
	.datac(!Xd_0__inst_r_sum1_7__7__q ),
	.datad(!Xd_0__inst_r_sum1_6__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_26 ),
	.sharein(Xd_0__inst_inst_add_4_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_29_sumout ),
	.cout(Xd_0__inst_inst_add_4_30 ),
	.shareout(Xd_0__inst_inst_add_4_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_29 (
// Equation(s):
// Xd_0__inst_inst_add_2_29_sumout  = SUM(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_30  = CARRY(( !Xd_0__inst_r_sum1_5__7__q  $ (!Xd_0__inst_r_sum1_4__7__q  $ (Xd_0__inst_r_sum1_3__7__q )) ) + ( Xd_0__inst_inst_add_2_27  ) + ( Xd_0__inst_inst_add_2_26  ))
// Xd_0__inst_inst_add_2_31  = SHARE((!Xd_0__inst_r_sum1_5__7__q  & (Xd_0__inst_r_sum1_4__7__q  & Xd_0__inst_r_sum1_3__7__q )) # (Xd_0__inst_r_sum1_5__7__q  & ((Xd_0__inst_r_sum1_3__7__q ) # (Xd_0__inst_r_sum1_4__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__7__q ),
	.datac(!Xd_0__inst_r_sum1_4__7__q ),
	.datad(!Xd_0__inst_r_sum1_3__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_26 ),
	.sharein(Xd_0__inst_inst_add_2_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_29_sumout ),
	.cout(Xd_0__inst_inst_add_2_30 ),
	.shareout(Xd_0__inst_inst_add_2_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_30  = CARRY(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_31  = SHARE((!Xd_0__inst_r_sum1_2__7__q  & (Xd_0__inst_r_sum1_1__7__q  & Xd_0__inst_r_sum1_0__7__q )) # (Xd_0__inst_r_sum1_2__7__q  & ((Xd_0__inst_r_sum1_0__7__q ) # (Xd_0__inst_r_sum1_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__7__q ),
	.datad(!Xd_0__inst_r_sum1_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_29 (
// Equation(s):
// Xd_0__inst_inst_add_8_29_sumout  = SUM(( !Xd_0__inst_r_sum1_14__7__q  $ (!Xd_0__inst_r_sum1_13__7__q  $ (Xd_0__inst_r_sum1_12__7__q )) ) + ( Xd_0__inst_inst_add_8_27  ) + ( Xd_0__inst_inst_add_8_26  ))
// Xd_0__inst_inst_add_8_30  = CARRY(( !Xd_0__inst_r_sum1_14__7__q  $ (!Xd_0__inst_r_sum1_13__7__q  $ (Xd_0__inst_r_sum1_12__7__q )) ) + ( Xd_0__inst_inst_add_8_27  ) + ( Xd_0__inst_inst_add_8_26  ))
// Xd_0__inst_inst_add_8_31  = SHARE((!Xd_0__inst_r_sum1_14__7__q  & (Xd_0__inst_r_sum1_13__7__q  & Xd_0__inst_r_sum1_12__7__q )) # (Xd_0__inst_r_sum1_14__7__q  & ((Xd_0__inst_r_sum1_12__7__q ) # (Xd_0__inst_r_sum1_13__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__7__q ),
	.datac(!Xd_0__inst_r_sum1_13__7__q ),
	.datad(!Xd_0__inst_r_sum1_12__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_26 ),
	.sharein(Xd_0__inst_inst_add_8_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_29_sumout ),
	.cout(Xd_0__inst_inst_add_8_30 ),
	.shareout(Xd_0__inst_inst_add_8_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_29 (
// Equation(s):
// Xd_0__inst_inst_add_6_29_sumout  = SUM(( !Xd_0__inst_r_sum1_11__7__q  $ (!Xd_0__inst_r_sum1_10__7__q  $ (Xd_0__inst_r_sum1_9__7__q )) ) + ( Xd_0__inst_inst_add_6_27  ) + ( Xd_0__inst_inst_add_6_26  ))
// Xd_0__inst_inst_add_6_30  = CARRY(( !Xd_0__inst_r_sum1_11__7__q  $ (!Xd_0__inst_r_sum1_10__7__q  $ (Xd_0__inst_r_sum1_9__7__q )) ) + ( Xd_0__inst_inst_add_6_27  ) + ( Xd_0__inst_inst_add_6_26  ))
// Xd_0__inst_inst_add_6_31  = SHARE((!Xd_0__inst_r_sum1_11__7__q  & (Xd_0__inst_r_sum1_10__7__q  & Xd_0__inst_r_sum1_9__7__q )) # (Xd_0__inst_r_sum1_11__7__q  & ((Xd_0__inst_r_sum1_9__7__q ) # (Xd_0__inst_r_sum1_10__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__7__q ),
	.datac(!Xd_0__inst_r_sum1_10__7__q ),
	.datad(!Xd_0__inst_r_sum1_9__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_26 ),
	.sharein(Xd_0__inst_inst_add_6_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_29_sumout ),
	.cout(Xd_0__inst_inst_add_6_30 ),
	.shareout(Xd_0__inst_inst_add_6_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_33 (
// Equation(s):
// Xd_0__inst_inst_add_4_33_sumout  = SUM(( !Xd_0__inst_r_sum1_8__8__q  $ (!Xd_0__inst_r_sum1_7__8__q  $ (Xd_0__inst_r_sum1_6__8__q )) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_34  = CARRY(( !Xd_0__inst_r_sum1_8__8__q  $ (!Xd_0__inst_r_sum1_7__8__q  $ (Xd_0__inst_r_sum1_6__8__q )) ) + ( Xd_0__inst_inst_add_4_31  ) + ( Xd_0__inst_inst_add_4_30  ))
// Xd_0__inst_inst_add_4_35  = SHARE((!Xd_0__inst_r_sum1_8__8__q  & (Xd_0__inst_r_sum1_7__8__q  & Xd_0__inst_r_sum1_6__8__q )) # (Xd_0__inst_r_sum1_8__8__q  & ((Xd_0__inst_r_sum1_6__8__q ) # (Xd_0__inst_r_sum1_7__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__8__q ),
	.datac(!Xd_0__inst_r_sum1_7__8__q ),
	.datad(!Xd_0__inst_r_sum1_6__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_30 ),
	.sharein(Xd_0__inst_inst_add_4_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_33_sumout ),
	.cout(Xd_0__inst_inst_add_4_34 ),
	.shareout(Xd_0__inst_inst_add_4_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_33 (
// Equation(s):
// Xd_0__inst_inst_add_2_33_sumout  = SUM(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_34  = CARRY(( !Xd_0__inst_r_sum1_5__8__q  $ (!Xd_0__inst_r_sum1_4__8__q  $ (Xd_0__inst_r_sum1_3__8__q )) ) + ( Xd_0__inst_inst_add_2_31  ) + ( Xd_0__inst_inst_add_2_30  ))
// Xd_0__inst_inst_add_2_35  = SHARE((!Xd_0__inst_r_sum1_5__8__q  & (Xd_0__inst_r_sum1_4__8__q  & Xd_0__inst_r_sum1_3__8__q )) # (Xd_0__inst_r_sum1_5__8__q  & ((Xd_0__inst_r_sum1_3__8__q ) # (Xd_0__inst_r_sum1_4__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__8__q ),
	.datac(!Xd_0__inst_r_sum1_4__8__q ),
	.datad(!Xd_0__inst_r_sum1_3__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_30 ),
	.sharein(Xd_0__inst_inst_add_2_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_33_sumout ),
	.cout(Xd_0__inst_inst_add_2_34 ),
	.shareout(Xd_0__inst_inst_add_2_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_34  = CARRY(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_35  = SHARE((!Xd_0__inst_r_sum1_2__8__q  & (Xd_0__inst_r_sum1_1__8__q  & Xd_0__inst_r_sum1_0__8__q )) # (Xd_0__inst_r_sum1_2__8__q  & ((Xd_0__inst_r_sum1_0__8__q ) # (Xd_0__inst_r_sum1_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__8__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_33 (
// Equation(s):
// Xd_0__inst_inst_add_8_33_sumout  = SUM(( !Xd_0__inst_r_sum1_14__8__q  $ (!Xd_0__inst_r_sum1_13__8__q  $ (Xd_0__inst_r_sum1_12__8__q )) ) + ( Xd_0__inst_inst_add_8_31  ) + ( Xd_0__inst_inst_add_8_30  ))
// Xd_0__inst_inst_add_8_34  = CARRY(( !Xd_0__inst_r_sum1_14__8__q  $ (!Xd_0__inst_r_sum1_13__8__q  $ (Xd_0__inst_r_sum1_12__8__q )) ) + ( Xd_0__inst_inst_add_8_31  ) + ( Xd_0__inst_inst_add_8_30  ))
// Xd_0__inst_inst_add_8_35  = SHARE((!Xd_0__inst_r_sum1_14__8__q  & (Xd_0__inst_r_sum1_13__8__q  & Xd_0__inst_r_sum1_12__8__q )) # (Xd_0__inst_r_sum1_14__8__q  & ((Xd_0__inst_r_sum1_12__8__q ) # (Xd_0__inst_r_sum1_13__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__8__q ),
	.datac(!Xd_0__inst_r_sum1_13__8__q ),
	.datad(!Xd_0__inst_r_sum1_12__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_30 ),
	.sharein(Xd_0__inst_inst_add_8_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_33_sumout ),
	.cout(Xd_0__inst_inst_add_8_34 ),
	.shareout(Xd_0__inst_inst_add_8_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_33 (
// Equation(s):
// Xd_0__inst_inst_add_6_33_sumout  = SUM(( !Xd_0__inst_r_sum1_11__8__q  $ (!Xd_0__inst_r_sum1_10__8__q  $ (Xd_0__inst_r_sum1_9__8__q )) ) + ( Xd_0__inst_inst_add_6_31  ) + ( Xd_0__inst_inst_add_6_30  ))
// Xd_0__inst_inst_add_6_34  = CARRY(( !Xd_0__inst_r_sum1_11__8__q  $ (!Xd_0__inst_r_sum1_10__8__q  $ (Xd_0__inst_r_sum1_9__8__q )) ) + ( Xd_0__inst_inst_add_6_31  ) + ( Xd_0__inst_inst_add_6_30  ))
// Xd_0__inst_inst_add_6_35  = SHARE((!Xd_0__inst_r_sum1_11__8__q  & (Xd_0__inst_r_sum1_10__8__q  & Xd_0__inst_r_sum1_9__8__q )) # (Xd_0__inst_r_sum1_11__8__q  & ((Xd_0__inst_r_sum1_9__8__q ) # (Xd_0__inst_r_sum1_10__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__8__q ),
	.datac(!Xd_0__inst_r_sum1_10__8__q ),
	.datad(!Xd_0__inst_r_sum1_9__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_30 ),
	.sharein(Xd_0__inst_inst_add_6_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_33_sumout ),
	.cout(Xd_0__inst_inst_add_6_34 ),
	.shareout(Xd_0__inst_inst_add_6_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_37 (
// Equation(s):
// Xd_0__inst_inst_add_4_37_sumout  = SUM(( !Xd_0__inst_r_sum1_8__9__q  $ (!Xd_0__inst_r_sum1_7__9__q  $ (Xd_0__inst_r_sum1_6__9__q )) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_38  = CARRY(( !Xd_0__inst_r_sum1_8__9__q  $ (!Xd_0__inst_r_sum1_7__9__q  $ (Xd_0__inst_r_sum1_6__9__q )) ) + ( Xd_0__inst_inst_add_4_35  ) + ( Xd_0__inst_inst_add_4_34  ))
// Xd_0__inst_inst_add_4_39  = SHARE((!Xd_0__inst_r_sum1_8__9__q  & (Xd_0__inst_r_sum1_7__9__q  & Xd_0__inst_r_sum1_6__9__q )) # (Xd_0__inst_r_sum1_8__9__q  & ((Xd_0__inst_r_sum1_6__9__q ) # (Xd_0__inst_r_sum1_7__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__9__q ),
	.datac(!Xd_0__inst_r_sum1_7__9__q ),
	.datad(!Xd_0__inst_r_sum1_6__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_34 ),
	.sharein(Xd_0__inst_inst_add_4_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_37_sumout ),
	.cout(Xd_0__inst_inst_add_4_38 ),
	.shareout(Xd_0__inst_inst_add_4_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_37 (
// Equation(s):
// Xd_0__inst_inst_add_2_37_sumout  = SUM(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_38  = CARRY(( !Xd_0__inst_r_sum1_5__9__q  $ (!Xd_0__inst_r_sum1_4__9__q  $ (Xd_0__inst_r_sum1_3__9__q )) ) + ( Xd_0__inst_inst_add_2_35  ) + ( Xd_0__inst_inst_add_2_34  ))
// Xd_0__inst_inst_add_2_39  = SHARE((!Xd_0__inst_r_sum1_5__9__q  & (Xd_0__inst_r_sum1_4__9__q  & Xd_0__inst_r_sum1_3__9__q )) # (Xd_0__inst_r_sum1_5__9__q  & ((Xd_0__inst_r_sum1_3__9__q ) # (Xd_0__inst_r_sum1_4__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__9__q ),
	.datac(!Xd_0__inst_r_sum1_4__9__q ),
	.datad(!Xd_0__inst_r_sum1_3__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_34 ),
	.sharein(Xd_0__inst_inst_add_2_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_37_sumout ),
	.cout(Xd_0__inst_inst_add_2_38 ),
	.shareout(Xd_0__inst_inst_add_2_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_38  = CARRY(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_39  = SHARE((!Xd_0__inst_r_sum1_2__9__q  & (Xd_0__inst_r_sum1_1__9__q  & Xd_0__inst_r_sum1_0__9__q )) # (Xd_0__inst_r_sum1_2__9__q  & ((Xd_0__inst_r_sum1_0__9__q ) # (Xd_0__inst_r_sum1_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__9__q ),
	.datad(!Xd_0__inst_r_sum1_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_37 (
// Equation(s):
// Xd_0__inst_inst_add_8_37_sumout  = SUM(( !Xd_0__inst_r_sum1_14__9__q  $ (!Xd_0__inst_r_sum1_13__9__q  $ (Xd_0__inst_r_sum1_12__9__q )) ) + ( Xd_0__inst_inst_add_8_35  ) + ( Xd_0__inst_inst_add_8_34  ))
// Xd_0__inst_inst_add_8_38  = CARRY(( !Xd_0__inst_r_sum1_14__9__q  $ (!Xd_0__inst_r_sum1_13__9__q  $ (Xd_0__inst_r_sum1_12__9__q )) ) + ( Xd_0__inst_inst_add_8_35  ) + ( Xd_0__inst_inst_add_8_34  ))
// Xd_0__inst_inst_add_8_39  = SHARE((!Xd_0__inst_r_sum1_14__9__q  & (Xd_0__inst_r_sum1_13__9__q  & Xd_0__inst_r_sum1_12__9__q )) # (Xd_0__inst_r_sum1_14__9__q  & ((Xd_0__inst_r_sum1_12__9__q ) # (Xd_0__inst_r_sum1_13__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__9__q ),
	.datac(!Xd_0__inst_r_sum1_13__9__q ),
	.datad(!Xd_0__inst_r_sum1_12__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_34 ),
	.sharein(Xd_0__inst_inst_add_8_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_37_sumout ),
	.cout(Xd_0__inst_inst_add_8_38 ),
	.shareout(Xd_0__inst_inst_add_8_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_37 (
// Equation(s):
// Xd_0__inst_inst_add_6_37_sumout  = SUM(( !Xd_0__inst_r_sum1_11__9__q  $ (!Xd_0__inst_r_sum1_10__9__q  $ (Xd_0__inst_r_sum1_9__9__q )) ) + ( Xd_0__inst_inst_add_6_35  ) + ( Xd_0__inst_inst_add_6_34  ))
// Xd_0__inst_inst_add_6_38  = CARRY(( !Xd_0__inst_r_sum1_11__9__q  $ (!Xd_0__inst_r_sum1_10__9__q  $ (Xd_0__inst_r_sum1_9__9__q )) ) + ( Xd_0__inst_inst_add_6_35  ) + ( Xd_0__inst_inst_add_6_34  ))
// Xd_0__inst_inst_add_6_39  = SHARE((!Xd_0__inst_r_sum1_11__9__q  & (Xd_0__inst_r_sum1_10__9__q  & Xd_0__inst_r_sum1_9__9__q )) # (Xd_0__inst_r_sum1_11__9__q  & ((Xd_0__inst_r_sum1_9__9__q ) # (Xd_0__inst_r_sum1_10__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__9__q ),
	.datac(!Xd_0__inst_r_sum1_10__9__q ),
	.datad(!Xd_0__inst_r_sum1_9__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_34 ),
	.sharein(Xd_0__inst_inst_add_6_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_37_sumout ),
	.cout(Xd_0__inst_inst_add_6_38 ),
	.shareout(Xd_0__inst_inst_add_6_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_41 (
// Equation(s):
// Xd_0__inst_inst_add_4_41_sumout  = SUM(( !Xd_0__inst_r_sum1_8__10__q  $ (!Xd_0__inst_r_sum1_7__10__q  $ (Xd_0__inst_r_sum1_6__10__q )) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_42  = CARRY(( !Xd_0__inst_r_sum1_8__10__q  $ (!Xd_0__inst_r_sum1_7__10__q  $ (Xd_0__inst_r_sum1_6__10__q )) ) + ( Xd_0__inst_inst_add_4_39  ) + ( Xd_0__inst_inst_add_4_38  ))
// Xd_0__inst_inst_add_4_43  = SHARE((!Xd_0__inst_r_sum1_8__10__q  & (Xd_0__inst_r_sum1_7__10__q  & Xd_0__inst_r_sum1_6__10__q )) # (Xd_0__inst_r_sum1_8__10__q  & ((Xd_0__inst_r_sum1_6__10__q ) # (Xd_0__inst_r_sum1_7__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__10__q ),
	.datac(!Xd_0__inst_r_sum1_7__10__q ),
	.datad(!Xd_0__inst_r_sum1_6__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_38 ),
	.sharein(Xd_0__inst_inst_add_4_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_41_sumout ),
	.cout(Xd_0__inst_inst_add_4_42 ),
	.shareout(Xd_0__inst_inst_add_4_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_41 (
// Equation(s):
// Xd_0__inst_inst_add_2_41_sumout  = SUM(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_42  = CARRY(( !Xd_0__inst_r_sum1_5__10__q  $ (!Xd_0__inst_r_sum1_4__10__q  $ (Xd_0__inst_r_sum1_3__10__q )) ) + ( Xd_0__inst_inst_add_2_39  ) + ( Xd_0__inst_inst_add_2_38  ))
// Xd_0__inst_inst_add_2_43  = SHARE((!Xd_0__inst_r_sum1_5__10__q  & (Xd_0__inst_r_sum1_4__10__q  & Xd_0__inst_r_sum1_3__10__q )) # (Xd_0__inst_r_sum1_5__10__q  & ((Xd_0__inst_r_sum1_3__10__q ) # (Xd_0__inst_r_sum1_4__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__10__q ),
	.datac(!Xd_0__inst_r_sum1_4__10__q ),
	.datad(!Xd_0__inst_r_sum1_3__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_38 ),
	.sharein(Xd_0__inst_inst_add_2_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_41_sumout ),
	.cout(Xd_0__inst_inst_add_2_42 ),
	.shareout(Xd_0__inst_inst_add_2_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_42  = CARRY(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_43  = SHARE((!Xd_0__inst_r_sum1_2__10__q  & (Xd_0__inst_r_sum1_1__10__q  & Xd_0__inst_r_sum1_0__10__q )) # (Xd_0__inst_r_sum1_2__10__q  & ((Xd_0__inst_r_sum1_0__10__q ) # (Xd_0__inst_r_sum1_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__10__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_41 (
// Equation(s):
// Xd_0__inst_inst_add_8_41_sumout  = SUM(( !Xd_0__inst_r_sum1_14__10__q  $ (!Xd_0__inst_r_sum1_13__10__q  $ (Xd_0__inst_r_sum1_12__10__q )) ) + ( Xd_0__inst_inst_add_8_39  ) + ( Xd_0__inst_inst_add_8_38  ))
// Xd_0__inst_inst_add_8_42  = CARRY(( !Xd_0__inst_r_sum1_14__10__q  $ (!Xd_0__inst_r_sum1_13__10__q  $ (Xd_0__inst_r_sum1_12__10__q )) ) + ( Xd_0__inst_inst_add_8_39  ) + ( Xd_0__inst_inst_add_8_38  ))
// Xd_0__inst_inst_add_8_43  = SHARE((!Xd_0__inst_r_sum1_14__10__q  & (Xd_0__inst_r_sum1_13__10__q  & Xd_0__inst_r_sum1_12__10__q )) # (Xd_0__inst_r_sum1_14__10__q  & ((Xd_0__inst_r_sum1_12__10__q ) # (Xd_0__inst_r_sum1_13__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__10__q ),
	.datac(!Xd_0__inst_r_sum1_13__10__q ),
	.datad(!Xd_0__inst_r_sum1_12__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_38 ),
	.sharein(Xd_0__inst_inst_add_8_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_41_sumout ),
	.cout(Xd_0__inst_inst_add_8_42 ),
	.shareout(Xd_0__inst_inst_add_8_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_41 (
// Equation(s):
// Xd_0__inst_inst_add_6_41_sumout  = SUM(( !Xd_0__inst_r_sum1_11__10__q  $ (!Xd_0__inst_r_sum1_10__10__q  $ (Xd_0__inst_r_sum1_9__10__q )) ) + ( Xd_0__inst_inst_add_6_39  ) + ( Xd_0__inst_inst_add_6_38  ))
// Xd_0__inst_inst_add_6_42  = CARRY(( !Xd_0__inst_r_sum1_11__10__q  $ (!Xd_0__inst_r_sum1_10__10__q  $ (Xd_0__inst_r_sum1_9__10__q )) ) + ( Xd_0__inst_inst_add_6_39  ) + ( Xd_0__inst_inst_add_6_38  ))
// Xd_0__inst_inst_add_6_43  = SHARE((!Xd_0__inst_r_sum1_11__10__q  & (Xd_0__inst_r_sum1_10__10__q  & Xd_0__inst_r_sum1_9__10__q )) # (Xd_0__inst_r_sum1_11__10__q  & ((Xd_0__inst_r_sum1_9__10__q ) # (Xd_0__inst_r_sum1_10__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__10__q ),
	.datac(!Xd_0__inst_r_sum1_10__10__q ),
	.datad(!Xd_0__inst_r_sum1_9__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_38 ),
	.sharein(Xd_0__inst_inst_add_6_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_41_sumout ),
	.cout(Xd_0__inst_inst_add_6_42 ),
	.shareout(Xd_0__inst_inst_add_6_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_45 (
// Equation(s):
// Xd_0__inst_inst_add_4_45_sumout  = SUM(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_46  = CARRY(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_43  ) + ( Xd_0__inst_inst_add_4_42  ))
// Xd_0__inst_inst_add_4_47  = SHARE((!Xd_0__inst_r_sum1_8__11__q  & (Xd_0__inst_r_sum1_7__11__q  & Xd_0__inst_r_sum1_6__11__q )) # (Xd_0__inst_r_sum1_8__11__q  & ((Xd_0__inst_r_sum1_6__11__q ) # (Xd_0__inst_r_sum1_7__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__11__q ),
	.datad(!Xd_0__inst_r_sum1_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_42 ),
	.sharein(Xd_0__inst_inst_add_4_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_45_sumout ),
	.cout(Xd_0__inst_inst_add_4_46 ),
	.shareout(Xd_0__inst_inst_add_4_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_45 (
// Equation(s):
// Xd_0__inst_inst_add_2_45_sumout  = SUM(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_46  = CARRY(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_43  ) + ( Xd_0__inst_inst_add_2_42  ))
// Xd_0__inst_inst_add_2_47  = SHARE((!Xd_0__inst_r_sum1_5__11__q  & (Xd_0__inst_r_sum1_4__11__q  & Xd_0__inst_r_sum1_3__11__q )) # (Xd_0__inst_r_sum1_5__11__q  & ((Xd_0__inst_r_sum1_3__11__q ) # (Xd_0__inst_r_sum1_4__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__11__q ),
	.datad(!Xd_0__inst_r_sum1_3__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_42 ),
	.sharein(Xd_0__inst_inst_add_2_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_45_sumout ),
	.cout(Xd_0__inst_inst_add_2_46 ),
	.shareout(Xd_0__inst_inst_add_2_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_46  = CARRY(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_47  = SHARE((!Xd_0__inst_r_sum1_2__11__q  & (Xd_0__inst_r_sum1_1__11__q  & Xd_0__inst_r_sum1_0__11__q )) # (Xd_0__inst_r_sum1_2__11__q  & ((Xd_0__inst_r_sum1_0__11__q ) # (Xd_0__inst_r_sum1_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_45 (
// Equation(s):
// Xd_0__inst_inst_add_8_45_sumout  = SUM(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_43  ) + ( Xd_0__inst_inst_add_8_42  ))
// Xd_0__inst_inst_add_8_46  = CARRY(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_43  ) + ( Xd_0__inst_inst_add_8_42  ))
// Xd_0__inst_inst_add_8_47  = SHARE((!Xd_0__inst_r_sum1_14__11__q  & (Xd_0__inst_r_sum1_13__11__q  & Xd_0__inst_r_sum1_12__11__q )) # (Xd_0__inst_r_sum1_14__11__q  & ((Xd_0__inst_r_sum1_12__11__q ) # (Xd_0__inst_r_sum1_13__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__11__q ),
	.datad(!Xd_0__inst_r_sum1_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_42 ),
	.sharein(Xd_0__inst_inst_add_8_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_45_sumout ),
	.cout(Xd_0__inst_inst_add_8_46 ),
	.shareout(Xd_0__inst_inst_add_8_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_45 (
// Equation(s):
// Xd_0__inst_inst_add_6_45_sumout  = SUM(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_43  ) + ( Xd_0__inst_inst_add_6_42  ))
// Xd_0__inst_inst_add_6_46  = CARRY(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_43  ) + ( Xd_0__inst_inst_add_6_42  ))
// Xd_0__inst_inst_add_6_47  = SHARE((!Xd_0__inst_r_sum1_11__11__q  & (Xd_0__inst_r_sum1_10__11__q  & Xd_0__inst_r_sum1_9__11__q )) # (Xd_0__inst_r_sum1_11__11__q  & ((Xd_0__inst_r_sum1_9__11__q ) # (Xd_0__inst_r_sum1_10__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__11__q ),
	.datad(!Xd_0__inst_r_sum1_9__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_42 ),
	.sharein(Xd_0__inst_inst_add_6_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_45_sumout ),
	.cout(Xd_0__inst_inst_add_6_46 ),
	.shareout(Xd_0__inst_inst_add_6_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_49 (
// Equation(s):
// Xd_0__inst_inst_add_4_49_sumout  = SUM(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_50  = CARRY(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_47  ) + ( Xd_0__inst_inst_add_4_46  ))
// Xd_0__inst_inst_add_4_51  = SHARE((!Xd_0__inst_r_sum1_8__11__q  & (Xd_0__inst_r_sum1_7__11__q  & Xd_0__inst_r_sum1_6__11__q )) # (Xd_0__inst_r_sum1_8__11__q  & ((Xd_0__inst_r_sum1_6__11__q ) # (Xd_0__inst_r_sum1_7__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__11__q ),
	.datad(!Xd_0__inst_r_sum1_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_46 ),
	.sharein(Xd_0__inst_inst_add_4_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_49_sumout ),
	.cout(Xd_0__inst_inst_add_4_50 ),
	.shareout(Xd_0__inst_inst_add_4_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_49 (
// Equation(s):
// Xd_0__inst_inst_add_2_49_sumout  = SUM(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_50  = CARRY(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_47  ) + ( Xd_0__inst_inst_add_2_46  ))
// Xd_0__inst_inst_add_2_51  = SHARE((!Xd_0__inst_r_sum1_5__11__q  & (Xd_0__inst_r_sum1_4__11__q  & Xd_0__inst_r_sum1_3__11__q )) # (Xd_0__inst_r_sum1_5__11__q  & ((Xd_0__inst_r_sum1_3__11__q ) # (Xd_0__inst_r_sum1_4__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__11__q ),
	.datad(!Xd_0__inst_r_sum1_3__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_46 ),
	.sharein(Xd_0__inst_inst_add_2_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_49_sumout ),
	.cout(Xd_0__inst_inst_add_2_50 ),
	.shareout(Xd_0__inst_inst_add_2_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_50  = CARRY(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_51  = SHARE((!Xd_0__inst_r_sum1_2__11__q  & (Xd_0__inst_r_sum1_1__11__q  & Xd_0__inst_r_sum1_0__11__q )) # (Xd_0__inst_r_sum1_2__11__q  & ((Xd_0__inst_r_sum1_0__11__q ) # (Xd_0__inst_r_sum1_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_49 (
// Equation(s):
// Xd_0__inst_inst_add_8_49_sumout  = SUM(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_47  ) + ( Xd_0__inst_inst_add_8_46  ))
// Xd_0__inst_inst_add_8_50  = CARRY(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_47  ) + ( Xd_0__inst_inst_add_8_46  ))
// Xd_0__inst_inst_add_8_51  = SHARE((!Xd_0__inst_r_sum1_14__11__q  & (Xd_0__inst_r_sum1_13__11__q  & Xd_0__inst_r_sum1_12__11__q )) # (Xd_0__inst_r_sum1_14__11__q  & ((Xd_0__inst_r_sum1_12__11__q ) # (Xd_0__inst_r_sum1_13__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__11__q ),
	.datad(!Xd_0__inst_r_sum1_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_46 ),
	.sharein(Xd_0__inst_inst_add_8_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_49_sumout ),
	.cout(Xd_0__inst_inst_add_8_50 ),
	.shareout(Xd_0__inst_inst_add_8_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_49 (
// Equation(s):
// Xd_0__inst_inst_add_6_49_sumout  = SUM(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_47  ) + ( Xd_0__inst_inst_add_6_46  ))
// Xd_0__inst_inst_add_6_50  = CARRY(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_47  ) + ( Xd_0__inst_inst_add_6_46  ))
// Xd_0__inst_inst_add_6_51  = SHARE((!Xd_0__inst_r_sum1_11__11__q  & (Xd_0__inst_r_sum1_10__11__q  & Xd_0__inst_r_sum1_9__11__q )) # (Xd_0__inst_r_sum1_11__11__q  & ((Xd_0__inst_r_sum1_9__11__q ) # (Xd_0__inst_r_sum1_10__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__11__q ),
	.datad(!Xd_0__inst_r_sum1_9__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_46 ),
	.sharein(Xd_0__inst_inst_add_6_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_49_sumout ),
	.cout(Xd_0__inst_inst_add_6_50 ),
	.shareout(Xd_0__inst_inst_add_6_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_4_53 (
// Equation(s):
// Xd_0__inst_inst_add_4_53_sumout  = SUM(( !Xd_0__inst_r_sum1_8__11__q  $ (!Xd_0__inst_r_sum1_7__11__q  $ (Xd_0__inst_r_sum1_6__11__q )) ) + ( Xd_0__inst_inst_add_4_51  ) + ( Xd_0__inst_inst_add_4_50  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_8__11__q ),
	.datac(!Xd_0__inst_r_sum1_7__11__q ),
	.datad(!Xd_0__inst_r_sum1_6__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_4_50 ),
	.sharein(Xd_0__inst_inst_add_4_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_4_53_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_2_53 (
// Equation(s):
// Xd_0__inst_inst_add_2_53_sumout  = SUM(( !Xd_0__inst_r_sum1_5__11__q  $ (!Xd_0__inst_r_sum1_4__11__q  $ (Xd_0__inst_r_sum1_3__11__q )) ) + ( Xd_0__inst_inst_add_2_51  ) + ( Xd_0__inst_inst_add_2_50  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_5__11__q ),
	.datac(!Xd_0__inst_r_sum1_4__11__q ),
	.datad(!Xd_0__inst_r_sum1_3__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_2_50 ),
	.sharein(Xd_0__inst_inst_add_2_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_2_53_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_53_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_8_53 (
// Equation(s):
// Xd_0__inst_inst_add_8_53_sumout  = SUM(( !Xd_0__inst_r_sum1_14__11__q  $ (!Xd_0__inst_r_sum1_13__11__q  $ (Xd_0__inst_r_sum1_12__11__q )) ) + ( Xd_0__inst_inst_add_8_51  ) + ( Xd_0__inst_inst_add_8_50  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_14__11__q ),
	.datac(!Xd_0__inst_r_sum1_13__11__q ),
	.datad(!Xd_0__inst_r_sum1_12__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_8_50 ),
	.sharein(Xd_0__inst_inst_add_8_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_8_53_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_6_53 (
// Equation(s):
// Xd_0__inst_inst_add_6_53_sumout  = SUM(( !Xd_0__inst_r_sum1_11__11__q  $ (!Xd_0__inst_r_sum1_10__11__q  $ (Xd_0__inst_r_sum1_9__11__q )) ) + ( Xd_0__inst_inst_add_6_51  ) + ( Xd_0__inst_inst_add_6_50  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_11__11__q ),
	.datac(!Xd_0__inst_r_sum1_10__11__q ),
	.datad(!Xd_0__inst_r_sum1_9__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_6_50 ),
	.sharein(Xd_0__inst_inst_add_6_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_6_53_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_35 (
// Equation(s):
// Xd_0__inst_mult_26_36  = SUM(( GND ) + ( Xd_0__inst_mult_26_42  ) + ( Xd_0__inst_mult_26_41  ))
// Xd_0__inst_mult_26_37  = CARRY(( GND ) + ( Xd_0__inst_mult_26_42  ) + ( Xd_0__inst_mult_26_41  ))
// Xd_0__inst_mult_26_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_41 ),
	.sharein(Xd_0__inst_mult_26_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_36 ),
	.cout(Xd_0__inst_mult_26_37 ),
	.shareout(Xd_0__inst_mult_26_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_35 (
// Equation(s):
// Xd_0__inst_mult_28_36  = SUM(( GND ) + ( Xd_0__inst_mult_28_42  ) + ( Xd_0__inst_mult_28_41  ))
// Xd_0__inst_mult_28_37  = CARRY(( GND ) + ( Xd_0__inst_mult_28_42  ) + ( Xd_0__inst_mult_28_41  ))
// Xd_0__inst_mult_28_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_41 ),
	.sharein(Xd_0__inst_mult_28_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_36 ),
	.cout(Xd_0__inst_mult_28_37 ),
	.shareout(Xd_0__inst_mult_28_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_35 (
// Equation(s):
// Xd_0__inst_mult_30_36  = SUM(( GND ) + ( Xd_0__inst_mult_30_42  ) + ( Xd_0__inst_mult_30_41  ))
// Xd_0__inst_mult_30_37  = CARRY(( GND ) + ( Xd_0__inst_mult_30_42  ) + ( Xd_0__inst_mult_30_41  ))
// Xd_0__inst_mult_30_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_41 ),
	.sharein(Xd_0__inst_mult_30_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_36 ),
	.cout(Xd_0__inst_mult_30_37 ),
	.shareout(Xd_0__inst_mult_30_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_16 (
// Equation(s):
// Xd_0__inst_mult_20_44  = CARRY(( GND ) + ( Xd_0__inst_i17_7  ) + ( Xd_0__inst_i17_6  ))
// Xd_0__inst_mult_20_45  = SHARE((din_b[123] & din_a[121]))

	.dataa(!din_b[123]),
	.datab(!din_a[121]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_6 ),
	.sharein(Xd_0__inst_i17_7 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_44 ),
	.shareout(Xd_0__inst_mult_20_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_35 (
// Equation(s):
// Xd_0__inst_mult_22_36  = SUM(( GND ) + ( Xd_0__inst_mult_22_42  ) + ( Xd_0__inst_mult_22_41  ))
// Xd_0__inst_mult_22_37  = CARRY(( GND ) + ( Xd_0__inst_mult_22_42  ) + ( Xd_0__inst_mult_22_41  ))
// Xd_0__inst_mult_22_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_41 ),
	.sharein(Xd_0__inst_mult_22_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_36 ),
	.cout(Xd_0__inst_mult_22_37 ),
	.shareout(Xd_0__inst_mult_22_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_35 (
// Equation(s):
// Xd_0__inst_mult_19_36  = SUM(( GND ) + ( Xd_0__inst_mult_19_42  ) + ( Xd_0__inst_mult_19_41  ))
// Xd_0__inst_mult_19_37  = CARRY(( GND ) + ( Xd_0__inst_mult_19_42  ) + ( Xd_0__inst_mult_19_41  ))
// Xd_0__inst_mult_19_38  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_41 ),
	.sharein(Xd_0__inst_mult_19_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_36 ),
	.cout(Xd_0__inst_mult_19_37 ),
	.shareout(Xd_0__inst_mult_19_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_30__0__q  $ (!Xd_0__inst_product_31__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_30__0__q  $ (!Xd_0__inst_product_31__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_30__0__q  & ((!Xd_0__inst_sign [31] & ((Xd_0__inst_sign [30]))) # (Xd_0__inst_sign [31] & (!Xd_0__inst_product_31__0__q )))) # (Xd_0__inst_product_30__0__q  & ((!Xd_0__inst_sign [31] 
// & (Xd_0__inst_product_31__0__q )) # (Xd_0__inst_sign [31] & ((!Xd_0__inst_sign [30]))))))

	.dataa(!Xd_0__inst_product_30__0__q ),
	.datab(!Xd_0__inst_product_31__0__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_16 (
// Equation(s):
// Xd_0__inst_mult_23_44  = CARRY(( GND ) + ( Xd_0__inst_i17_11  ) + ( Xd_0__inst_i17_10  ))
// Xd_0__inst_mult_23_45  = SHARE((din_b[141] & din_a[139]))

	.dataa(!din_b[141]),
	.datab(!din_a[139]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_10 ),
	.sharein(Xd_0__inst_i17_11 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_44 ),
	.shareout(Xd_0__inst_mult_23_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_30__1__q  $ (!Xd_0__inst_product_31__1__q  $ (((Xd_0__inst_sign [31]) # (Xd_0__inst_sign [30])))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_30__1__q  $ (!Xd_0__inst_product_31__1__q  $ (((Xd_0__inst_sign [31]) # (Xd_0__inst_sign [30])))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [30] & (Xd_0__inst_product_30__1__q  & (!Xd_0__inst_product_31__1__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_sign [30] & ((!Xd_0__inst_product_31__1__q  & ((Xd_0__inst_sign [31]))) 
// # (Xd_0__inst_product_31__1__q  & (!Xd_0__inst_product_30__1__q )))))

	.dataa(!Xd_0__inst_product_30__1__q ),
	.datab(!Xd_0__inst_product_31__1__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_30__2__q  $ (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_30__2__q  $ (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__2__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__2__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__2__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__2__q ),
	.datab(!Xd_0__inst_product_31__2__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_30__3__q  $ (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_30__3__q  $ (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__3__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__3__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__3__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__3__q ),
	.datab(!Xd_0__inst_product_31__3__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_30__4__q  $ (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_30__4__q  $ (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__4__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__4__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__4__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__4__q ),
	.datab(!Xd_0__inst_product_31__4__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_30__5__q  $ (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_30__5__q  $ (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__5__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__5__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__5__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__5__q ),
	.datab(!Xd_0__inst_product_31__5__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_30__6__q  $ (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_30__6__q  $ (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__6__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__6__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__6__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__6__q ),
	.datab(!Xd_0__inst_product_31__6__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_30__7__q  $ (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_30__7__q  $ (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__7__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__7__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__7__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__7__q ),
	.datab(!Xd_0__inst_product_31__7__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_30__8__q  $ (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_30__8__q  $ (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__8__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__8__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__8__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__8__q ),
	.datab(!Xd_0__inst_product_31__8__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_30__9__q  $ (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_30__9__q  $ (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]))) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_30__9__q  & (Xd_0__inst_sign [30] & (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [31])))) # (Xd_0__inst_product_30__9__q  & (!Xd_0__inst_sign [30] & 
// (!Xd_0__inst_product_31__9__q  $ (!Xd_0__inst_sign [31])))))

	.dataa(!Xd_0__inst_product_30__9__q ),
	.datab(!Xd_0__inst_product_31__9__q ),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_15__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_15__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [30] & Xd_0__inst_sign [31]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [30]),
	.datad(!Xd_0__inst_sign [31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_15__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_34 (
// Equation(s):
// Xd_0__inst_mult_2_35  = SUM(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_2_36  = CARRY(( !Xd_0__inst_sign [30] $ (!Xd_0__inst_sign [31]) ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_15__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_2_37  = SHARE((Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_1_q ))

	.dataa(!Xd_0__inst_sign [30]),
	.datab(!Xd_0__inst_sign [31]),
	.datac(!Xd_0__inst_mult_2_0_q ),
	.datad(!Xd_0__inst_mult_2_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_15__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_15__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_35 ),
	.cout(Xd_0__inst_mult_2_36 ),
	.shareout(Xd_0__inst_mult_2_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_16__0__q  $ (!Xd_0__inst_product_17__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_16__0__q  $ (!Xd_0__inst_product_17__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_16__0__q  & ((!Xd_0__inst_sign [17] & ((Xd_0__inst_sign [16]))) # (Xd_0__inst_sign [17] & (!Xd_0__inst_product_17__0__q )))) # (Xd_0__inst_product_16__0__q  & ((!Xd_0__inst_sign [17] 
// & (Xd_0__inst_product_17__0__q )) # (Xd_0__inst_sign [17] & ((!Xd_0__inst_sign [16]))))))

	.dataa(!Xd_0__inst_product_16__0__q ),
	.datab(!Xd_0__inst_product_17__0__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_14__0__q  $ (!Xd_0__inst_product_15__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] & ((Xd_0__inst_sign [14]))) # (Xd_0__inst_sign [15] & (!Xd_0__inst_product_15__0__q )))) # (Xd_0__inst_product_14__0__q  & ((!Xd_0__inst_sign [15] 
// & (Xd_0__inst_product_15__0__q )) # (Xd_0__inst_sign [15] & ((!Xd_0__inst_sign [14]))))))

	.dataa(!Xd_0__inst_product_14__0__q ),
	.datab(!Xd_0__inst_product_15__0__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_12__0__q  $ (!Xd_0__inst_product_13__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] & ((Xd_0__inst_sign [12]))) # (Xd_0__inst_sign [13] & (!Xd_0__inst_product_13__0__q )))) # (Xd_0__inst_product_12__0__q  & ((!Xd_0__inst_sign [13] 
// & (Xd_0__inst_product_13__0__q )) # (Xd_0__inst_sign [13] & ((!Xd_0__inst_sign [12]))))))

	.dataa(!Xd_0__inst_product_12__0__q ),
	.datab(!Xd_0__inst_product_13__0__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26 (
// Equation(s):
// Xd_0__inst_mult_26_40  = SUM(( (!din_a[160] & (((din_a[159] & din_b[157])))) # (din_a[160] & (!din_b[156] $ (((!din_a[159]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_26_49  ) + ( Xd_0__inst_mult_26_48  ))
// Xd_0__inst_mult_26_41  = CARRY(( (!din_a[160] & (((din_a[159] & din_b[157])))) # (din_a[160] & (!din_b[156] $ (((!din_a[159]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_26_49  ) + ( Xd_0__inst_mult_26_48  ))
// Xd_0__inst_mult_26_42  = SHARE((din_a[160] & (din_b[156] & (din_a[159] & din_b[157]))))

	.dataa(!din_a[160]),
	.datab(!din_b[156]),
	.datac(!din_a[159]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_48 ),
	.sharein(Xd_0__inst_mult_26_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_40 ),
	.cout(Xd_0__inst_mult_26_41 ),
	.shareout(Xd_0__inst_mult_26_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_10__0__q  $ (!Xd_0__inst_product_11__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] & ((Xd_0__inst_sign [10]))) # (Xd_0__inst_sign [11] & (!Xd_0__inst_product_11__0__q )))) # (Xd_0__inst_product_10__0__q  & ((!Xd_0__inst_sign [11] 
// & (Xd_0__inst_product_11__0__q )) # (Xd_0__inst_sign [11] & ((!Xd_0__inst_sign [10]))))))

	.dataa(!Xd_0__inst_product_10__0__q ),
	.datab(!Xd_0__inst_product_11__0__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_4__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_8__0__q  $ (!Xd_0__inst_product_9__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & ((Xd_0__inst_sign [8]))) # (Xd_0__inst_sign [9] & (!Xd_0__inst_product_9__0__q )))) # (Xd_0__inst_product_8__0__q  & ((!Xd_0__inst_sign [9] & 
// (Xd_0__inst_product_9__0__q )) # (Xd_0__inst_sign [9] & ((!Xd_0__inst_sign [8]))))))

	.dataa(!Xd_0__inst_product_8__0__q ),
	.datab(!Xd_0__inst_product_9__0__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_3__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & ((Xd_0__inst_sign [6]))) # (Xd_0__inst_sign [7] & (!Xd_0__inst_product_7__0__q )))) # (Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & 
// (Xd_0__inst_product_7__0__q )) # (Xd_0__inst_sign [7] & ((!Xd_0__inst_sign [6]))))))

	.dataa(!Xd_0__inst_product_6__0__q ),
	.datab(!Xd_0__inst_product_7__0__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28 (
// Equation(s):
// Xd_0__inst_mult_28_40  = SUM(( (!din_a[172] & (((din_a[171] & din_b[169])))) # (din_a[172] & (!din_b[168] $ (((!din_a[171]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_28_49  ) + ( Xd_0__inst_mult_28_48  ))
// Xd_0__inst_mult_28_41  = CARRY(( (!din_a[172] & (((din_a[171] & din_b[169])))) # (din_a[172] & (!din_b[168] $ (((!din_a[171]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_28_49  ) + ( Xd_0__inst_mult_28_48  ))
// Xd_0__inst_mult_28_42  = SHARE((din_a[172] & (din_b[168] & (din_a[171] & din_b[169]))))

	.dataa(!din_a[172]),
	.datab(!din_b[168]),
	.datac(!din_a[171]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_48 ),
	.sharein(Xd_0__inst_mult_28_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_40 ),
	.cout(Xd_0__inst_mult_28_41 ),
	.shareout(Xd_0__inst_mult_28_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_2__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & ((Xd_0__inst_sign [4]))) # (Xd_0__inst_sign [5] & (!Xd_0__inst_product_5__0__q )))) # (Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & 
// (Xd_0__inst_product_5__0__q )) # (Xd_0__inst_sign [5] & ((!Xd_0__inst_sign [4]))))))

	.dataa(!Xd_0__inst_product_4__0__q ),
	.datab(!Xd_0__inst_product_5__0__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_1__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & ((Xd_0__inst_sign [2]))) # (Xd_0__inst_sign [3] & (!Xd_0__inst_product_3__0__q )))) # (Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & 
// (Xd_0__inst_product_3__0__q )) # (Xd_0__inst_sign [3] & ((!Xd_0__inst_sign [2]))))))

	.dataa(!Xd_0__inst_product_2__0__q ),
	.datab(!Xd_0__inst_product_3__0__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_0__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & ((Xd_0__inst_sign [0]))) # (Xd_0__inst_sign [1] & (!Xd_0__inst_product_1__0__q )))) # (Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & 
// (Xd_0__inst_product_1__0__q )) # (Xd_0__inst_sign [1] & ((!Xd_0__inst_sign [0]))))))

	.dataa(!Xd_0__inst_product_0__0__q ),
	.datab(!Xd_0__inst_product_1__0__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30 (
// Equation(s):
// Xd_0__inst_mult_30_40  = SUM(( (!din_a[184] & (((din_a[183] & din_b[181])))) # (din_a[184] & (!din_b[180] $ (((!din_a[183]) # (!din_b[181]))))) ) + ( Xd_0__inst_mult_30_49  ) + ( Xd_0__inst_mult_30_48  ))
// Xd_0__inst_mult_30_41  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[181])))) # (din_a[184] & (!din_b[180] $ (((!din_a[183]) # (!din_b[181]))))) ) + ( Xd_0__inst_mult_30_49  ) + ( Xd_0__inst_mult_30_48  ))
// Xd_0__inst_mult_30_42  = SHARE((din_a[184] & (din_b[180] & (din_a[183] & din_b[181]))))

	.dataa(!din_a[184]),
	.datab(!din_b[180]),
	.datac(!din_a[183]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_48 ),
	.sharein(Xd_0__inst_mult_30_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_40 ),
	.cout(Xd_0__inst_mult_30_41 ),
	.shareout(Xd_0__inst_mult_30_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_5 (
// Equation(s):
// Xd_0__inst_i17_5_sumout  = SUM(( !din_a[107] $ (!din_b[107]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_6  = CARRY(( !din_a[107] $ (!din_b[107]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_7  = SHARE(GND)

	.dataa(!din_a[107]),
	.datab(!din_b[107]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_5_sumout ),
	.cout(Xd_0__inst_i17_6 ),
	.shareout(Xd_0__inst_i17_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_28__0__q  $ (!Xd_0__inst_product_29__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_28__0__q  $ (!Xd_0__inst_product_29__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_28__0__q  & ((!Xd_0__inst_sign [29] & ((Xd_0__inst_sign [28]))) # (Xd_0__inst_sign [29] & (!Xd_0__inst_product_29__0__q )))) # (Xd_0__inst_product_28__0__q  & ((!Xd_0__inst_sign [29] 
// & (Xd_0__inst_product_29__0__q )) # (Xd_0__inst_sign [29] & ((!Xd_0__inst_sign [28]))))))

	.dataa(!Xd_0__inst_product_28__0__q ),
	.datab(!Xd_0__inst_product_29__0__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_26__0__q  $ (!Xd_0__inst_product_27__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_26__0__q  $ (!Xd_0__inst_product_27__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_26__0__q  & ((!Xd_0__inst_sign [27] & ((Xd_0__inst_sign [26]))) # (Xd_0__inst_sign [27] & (!Xd_0__inst_product_27__0__q )))) # (Xd_0__inst_product_26__0__q  & ((!Xd_0__inst_sign [27] 
// & (Xd_0__inst_product_27__0__q )) # (Xd_0__inst_sign [27] & ((!Xd_0__inst_sign [26]))))))

	.dataa(!Xd_0__inst_product_26__0__q ),
	.datab(!Xd_0__inst_product_27__0__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_24__0__q  $ (!Xd_0__inst_product_25__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_24__0__q  $ (!Xd_0__inst_product_25__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_24__0__q  & ((!Xd_0__inst_sign [25] & ((Xd_0__inst_sign [24]))) # (Xd_0__inst_sign [25] & (!Xd_0__inst_product_25__0__q )))) # (Xd_0__inst_product_24__0__q  & ((!Xd_0__inst_sign [25] 
// & (Xd_0__inst_product_25__0__q )) # (Xd_0__inst_sign [25] & ((!Xd_0__inst_sign [24]))))))

	.dataa(!Xd_0__inst_product_24__0__q ),
	.datab(!Xd_0__inst_product_25__0__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22 (
// Equation(s):
// Xd_0__inst_mult_22_40  = SUM(( (!din_a[136] & (((din_a[135] & din_b[133])))) # (din_a[136] & (!din_b[132] $ (((!din_a[135]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_22_49  ) + ( Xd_0__inst_mult_22_48  ))
// Xd_0__inst_mult_22_41  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[133])))) # (din_a[136] & (!din_b[132] $ (((!din_a[135]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_22_49  ) + ( Xd_0__inst_mult_22_48  ))
// Xd_0__inst_mult_22_42  = SHARE((din_a[136] & (din_b[132] & (din_a[135] & din_b[133]))))

	.dataa(!din_a[136]),
	.datab(!din_b[132]),
	.datac(!din_a[135]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_48 ),
	.sharein(Xd_0__inst_mult_22_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_40 ),
	.cout(Xd_0__inst_mult_22_41 ),
	.shareout(Xd_0__inst_mult_22_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_22__0__q  $ (!Xd_0__inst_product_23__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_22__0__q  $ (!Xd_0__inst_product_23__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_22__0__q  & ((!Xd_0__inst_sign [23] & ((Xd_0__inst_sign [22]))) # (Xd_0__inst_sign [23] & (!Xd_0__inst_product_23__0__q )))) # (Xd_0__inst_product_22__0__q  & ((!Xd_0__inst_sign [23] 
// & (Xd_0__inst_product_23__0__q )) # (Xd_0__inst_sign [23] & ((!Xd_0__inst_sign [22]))))))

	.dataa(!Xd_0__inst_product_22__0__q ),
	.datab(!Xd_0__inst_product_23__0__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_20__0__q  $ (!Xd_0__inst_product_21__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_20__0__q  $ (!Xd_0__inst_product_21__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_20__0__q  & ((!Xd_0__inst_sign [21] & ((Xd_0__inst_sign [20]))) # (Xd_0__inst_sign [21] & (!Xd_0__inst_product_21__0__q )))) # (Xd_0__inst_product_20__0__q  & ((!Xd_0__inst_sign [21] 
// & (Xd_0__inst_product_21__0__q )) # (Xd_0__inst_sign [21] & ((!Xd_0__inst_sign [20]))))))

	.dataa(!Xd_0__inst_product_20__0__q ),
	.datab(!Xd_0__inst_product_21__0__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_18__0__q  $ (!Xd_0__inst_product_19__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_18__0__q  $ (!Xd_0__inst_product_19__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_18__0__q  & ((!Xd_0__inst_sign [19] & ((Xd_0__inst_sign [18]))) # (Xd_0__inst_sign [19] & (!Xd_0__inst_product_19__0__q )))) # (Xd_0__inst_product_18__0__q  & ((!Xd_0__inst_sign [19] 
// & (Xd_0__inst_product_19__0__q )) # (Xd_0__inst_sign [19] & ((!Xd_0__inst_sign [18]))))))

	.dataa(!Xd_0__inst_product_18__0__q ),
	.datab(!Xd_0__inst_product_19__0__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19 (
// Equation(s):
// Xd_0__inst_mult_19_40  = SUM(( (!din_a[118] & (((din_a[117] & din_b[115])))) # (din_a[118] & (!din_b[114] $ (((!din_a[117]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_19_45  ) + ( Xd_0__inst_mult_19_44  ))
// Xd_0__inst_mult_19_41  = CARRY(( (!din_a[118] & (((din_a[117] & din_b[115])))) # (din_a[118] & (!din_b[114] $ (((!din_a[117]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_19_45  ) + ( Xd_0__inst_mult_19_44  ))
// Xd_0__inst_mult_19_42  = SHARE((din_a[118] & (din_b[114] & (din_a[117] & din_b[115]))))

	.dataa(!din_a[118]),
	.datab(!din_b[114]),
	.datac(!din_a[117]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_44 ),
	.sharein(Xd_0__inst_mult_19_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_40 ),
	.cout(Xd_0__inst_mult_19_41 ),
	.shareout(Xd_0__inst_mult_19_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_9 (
// Equation(s):
// Xd_0__inst_i17_9_sumout  = SUM(( !din_a[161] $ (!din_b[161]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_10  = CARRY(( !din_a[161] $ (!din_b[161]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_11  = SHARE(GND)

	.dataa(!din_a[161]),
	.datab(!din_b[161]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_9_sumout ),
	.cout(Xd_0__inst_i17_10 ),
	.shareout(Xd_0__inst_i17_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_16__1__q  $ (!Xd_0__inst_product_17__1__q  $ (((Xd_0__inst_sign [17]) # (Xd_0__inst_sign [16])))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_16__1__q  $ (!Xd_0__inst_product_17__1__q  $ (((Xd_0__inst_sign [17]) # (Xd_0__inst_sign [16])))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [16] & (Xd_0__inst_product_16__1__q  & (!Xd_0__inst_product_17__1__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_sign [16] & ((!Xd_0__inst_product_17__1__q  & ((Xd_0__inst_sign [17]))) # 
// (Xd_0__inst_product_17__1__q  & (!Xd_0__inst_product_16__1__q )))))

	.dataa(!Xd_0__inst_product_16__1__q ),
	.datab(!Xd_0__inst_product_17__1__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_14__1__q  $ (!Xd_0__inst_product_15__1__q  $ (((Xd_0__inst_sign [15]) # (Xd_0__inst_sign [14])))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [14] & (Xd_0__inst_product_14__1__q  & (!Xd_0__inst_product_15__1__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_sign [14] & ((!Xd_0__inst_product_15__1__q  & ((Xd_0__inst_sign [15]))) # 
// (Xd_0__inst_product_15__1__q  & (!Xd_0__inst_product_14__1__q )))))

	.dataa(!Xd_0__inst_product_14__1__q ),
	.datab(!Xd_0__inst_product_15__1__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_12__1__q  $ (!Xd_0__inst_product_13__1__q  $ (((Xd_0__inst_sign [13]) # (Xd_0__inst_sign [12])))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [12] & (Xd_0__inst_product_12__1__q  & (!Xd_0__inst_product_13__1__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_sign [12] & ((!Xd_0__inst_product_13__1__q  & ((Xd_0__inst_sign [13]))) # 
// (Xd_0__inst_product_13__1__q  & (!Xd_0__inst_product_12__1__q )))))

	.dataa(!Xd_0__inst_product_12__1__q ),
	.datab(!Xd_0__inst_product_13__1__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_10__1__q  $ (!Xd_0__inst_product_11__1__q  $ (((Xd_0__inst_sign [11]) # (Xd_0__inst_sign [10])))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [10] & (Xd_0__inst_product_10__1__q  & (!Xd_0__inst_product_11__1__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_sign [10] & ((!Xd_0__inst_product_11__1__q  & ((Xd_0__inst_sign [11]))) # 
// (Xd_0__inst_product_11__1__q  & (!Xd_0__inst_product_10__1__q )))))

	.dataa(!Xd_0__inst_product_10__1__q ),
	.datab(!Xd_0__inst_product_11__1__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_8__1__q  $ (!Xd_0__inst_product_9__1__q  $ (((Xd_0__inst_sign [9]) # (Xd_0__inst_sign [8])))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [8] & (Xd_0__inst_product_8__1__q  & (!Xd_0__inst_product_9__1__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_sign [8] & ((!Xd_0__inst_product_9__1__q  & ((Xd_0__inst_sign [9]))) # 
// (Xd_0__inst_product_9__1__q  & (!Xd_0__inst_product_8__1__q )))))

	.dataa(!Xd_0__inst_product_8__1__q ),
	.datab(!Xd_0__inst_product_9__1__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [6] & (Xd_0__inst_product_6__1__q  & (!Xd_0__inst_product_7__1__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_sign [6] & ((!Xd_0__inst_product_7__1__q  & ((Xd_0__inst_sign [7]))) # 
// (Xd_0__inst_product_7__1__q  & (!Xd_0__inst_product_6__1__q )))))

	.dataa(!Xd_0__inst_product_6__1__q ),
	.datab(!Xd_0__inst_product_7__1__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [4] & (Xd_0__inst_product_4__1__q  & (!Xd_0__inst_product_5__1__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_sign [4] & ((!Xd_0__inst_product_5__1__q  & ((Xd_0__inst_sign [5]))) # 
// (Xd_0__inst_product_5__1__q  & (!Xd_0__inst_product_4__1__q )))))

	.dataa(!Xd_0__inst_product_4__1__q ),
	.datab(!Xd_0__inst_product_5__1__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [2] & (Xd_0__inst_product_2__1__q  & (!Xd_0__inst_product_3__1__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_sign [2] & ((!Xd_0__inst_product_3__1__q  & ((Xd_0__inst_sign [3]))) # 
// (Xd_0__inst_product_3__1__q  & (!Xd_0__inst_product_2__1__q )))))

	.dataa(!Xd_0__inst_product_2__1__q ),
	.datab(!Xd_0__inst_product_3__1__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [0] & (Xd_0__inst_product_0__1__q  & (!Xd_0__inst_product_1__1__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_sign [0] & ((!Xd_0__inst_product_1__1__q  & ((Xd_0__inst_sign [1]))) # 
// (Xd_0__inst_product_1__1__q  & (!Xd_0__inst_product_0__1__q )))))

	.dataa(!Xd_0__inst_product_0__1__q ),
	.datab(!Xd_0__inst_product_1__1__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_28__1__q  $ (!Xd_0__inst_product_29__1__q  $ (((Xd_0__inst_sign [29]) # (Xd_0__inst_sign [28])))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_28__1__q  $ (!Xd_0__inst_product_29__1__q  $ (((Xd_0__inst_sign [29]) # (Xd_0__inst_sign [28])))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [28] & (Xd_0__inst_product_28__1__q  & (!Xd_0__inst_product_29__1__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_sign [28] & ((!Xd_0__inst_product_29__1__q  & ((Xd_0__inst_sign [29]))) 
// # (Xd_0__inst_product_29__1__q  & (!Xd_0__inst_product_28__1__q )))))

	.dataa(!Xd_0__inst_product_28__1__q ),
	.datab(!Xd_0__inst_product_29__1__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_26__1__q  $ (!Xd_0__inst_product_27__1__q  $ (((Xd_0__inst_sign [27]) # (Xd_0__inst_sign [26])))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_26__1__q  $ (!Xd_0__inst_product_27__1__q  $ (((Xd_0__inst_sign [27]) # (Xd_0__inst_sign [26])))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [26] & (Xd_0__inst_product_26__1__q  & (!Xd_0__inst_product_27__1__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_sign [26] & ((!Xd_0__inst_product_27__1__q  & ((Xd_0__inst_sign [27]))) 
// # (Xd_0__inst_product_27__1__q  & (!Xd_0__inst_product_26__1__q )))))

	.dataa(!Xd_0__inst_product_26__1__q ),
	.datab(!Xd_0__inst_product_27__1__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_24__1__q  $ (!Xd_0__inst_product_25__1__q  $ (((Xd_0__inst_sign [25]) # (Xd_0__inst_sign [24])))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_24__1__q  $ (!Xd_0__inst_product_25__1__q  $ (((Xd_0__inst_sign [25]) # (Xd_0__inst_sign [24])))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [24] & (Xd_0__inst_product_24__1__q  & (!Xd_0__inst_product_25__1__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_sign [24] & ((!Xd_0__inst_product_25__1__q  & ((Xd_0__inst_sign [25]))) 
// # (Xd_0__inst_product_25__1__q  & (!Xd_0__inst_product_24__1__q )))))

	.dataa(!Xd_0__inst_product_24__1__q ),
	.datab(!Xd_0__inst_product_25__1__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_22__1__q  $ (!Xd_0__inst_product_23__1__q  $ (((Xd_0__inst_sign [23]) # (Xd_0__inst_sign [22])))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_22__1__q  $ (!Xd_0__inst_product_23__1__q  $ (((Xd_0__inst_sign [23]) # (Xd_0__inst_sign [22])))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [22] & (Xd_0__inst_product_22__1__q  & (!Xd_0__inst_product_23__1__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_sign [22] & ((!Xd_0__inst_product_23__1__q  & ((Xd_0__inst_sign [23]))) 
// # (Xd_0__inst_product_23__1__q  & (!Xd_0__inst_product_22__1__q )))))

	.dataa(!Xd_0__inst_product_22__1__q ),
	.datab(!Xd_0__inst_product_23__1__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_20__1__q  $ (!Xd_0__inst_product_21__1__q  $ (((Xd_0__inst_sign [21]) # (Xd_0__inst_sign [20])))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_20__1__q  $ (!Xd_0__inst_product_21__1__q  $ (((Xd_0__inst_sign [21]) # (Xd_0__inst_sign [20])))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [20] & (Xd_0__inst_product_20__1__q  & (!Xd_0__inst_product_21__1__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_sign [20] & ((!Xd_0__inst_product_21__1__q  & ((Xd_0__inst_sign [21]))) 
// # (Xd_0__inst_product_21__1__q  & (!Xd_0__inst_product_20__1__q )))))

	.dataa(!Xd_0__inst_product_20__1__q ),
	.datab(!Xd_0__inst_product_21__1__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_18__1__q  $ (!Xd_0__inst_product_19__1__q  $ (((Xd_0__inst_sign [19]) # (Xd_0__inst_sign [18])))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_18__1__q  $ (!Xd_0__inst_product_19__1__q  $ (((Xd_0__inst_sign [19]) # (Xd_0__inst_sign [18])))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc0_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [18] & (Xd_0__inst_product_18__1__q  & (!Xd_0__inst_product_19__1__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_sign [18] & ((!Xd_0__inst_product_19__1__q  & ((Xd_0__inst_sign [19]))) # 
// (Xd_0__inst_product_19__1__q  & (!Xd_0__inst_product_18__1__q )))))

	.dataa(!Xd_0__inst_product_18__1__q ),
	.datab(!Xd_0__inst_product_19__1__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_16__2__q  $ (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_16__2__q  $ (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__2__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__2__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__2__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__2__q ),
	.datab(!Xd_0__inst_product_17__2__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_14__2__q  $ (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__2__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__2__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__2__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__2__q ),
	.datab(!Xd_0__inst_product_15__2__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_12__2__q  $ (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__2__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__2__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__2__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__2__q ),
	.datab(!Xd_0__inst_product_13__2__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_10__2__q  $ (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__2__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__2__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__2__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__2__q ),
	.datab(!Xd_0__inst_product_11__2__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_8__2__q  $ (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__2__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__2__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__2__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__2__q ),
	.datab(!Xd_0__inst_product_9__2__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__2__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__2__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__2__q ),
	.datab(!Xd_0__inst_product_7__2__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__2__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__2__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__2__q ),
	.datab(!Xd_0__inst_product_5__2__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__2__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__2__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__2__q ),
	.datab(!Xd_0__inst_product_3__2__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__2__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__2__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__2__q ),
	.datab(!Xd_0__inst_product_1__2__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_28__2__q  $ (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_28__2__q  $ (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__2__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__2__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__2__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__2__q ),
	.datab(!Xd_0__inst_product_29__2__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_26__2__q  $ (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_26__2__q  $ (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__2__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__2__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__2__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__2__q ),
	.datab(!Xd_0__inst_product_27__2__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_24__2__q  $ (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_24__2__q  $ (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__2__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__2__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__2__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__2__q ),
	.datab(!Xd_0__inst_product_25__2__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_22__2__q  $ (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_22__2__q  $ (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__2__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__2__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__2__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__2__q ),
	.datab(!Xd_0__inst_product_23__2__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_20__2__q  $ (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_20__2__q  $ (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__2__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__2__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__2__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__2__q ),
	.datab(!Xd_0__inst_product_21__2__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_18__2__q  $ (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_COUT  
// ))
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_18__2__q  $ (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__2__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__2__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__2__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__2__q ),
	.datab(!Xd_0__inst_product_19__2__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_16__3__q  $ (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_16__3__q  $ (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__3__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__3__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__3__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__3__q ),
	.datab(!Xd_0__inst_product_17__3__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_14__3__q  $ (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__3__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__3__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__3__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__3__q ),
	.datab(!Xd_0__inst_product_15__3__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_12__3__q  $ (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__3__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__3__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__3__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__3__q ),
	.datab(!Xd_0__inst_product_13__3__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_10__3__q  $ (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__3__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__3__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__3__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__3__q ),
	.datab(!Xd_0__inst_product_11__3__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_8__3__q  $ (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__3__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__3__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__3__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__3__q ),
	.datab(!Xd_0__inst_product_9__3__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__3__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__3__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__3__q ),
	.datab(!Xd_0__inst_product_7__3__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__3__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__3__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__3__q ),
	.datab(!Xd_0__inst_product_5__3__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__3__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__3__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__3__q ),
	.datab(!Xd_0__inst_product_3__3__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__3__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__3__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__3__q ),
	.datab(!Xd_0__inst_product_1__3__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_28__3__q  $ (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_28__3__q  $ (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__3__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__3__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__3__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__3__q ),
	.datab(!Xd_0__inst_product_29__3__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_26__3__q  $ (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_26__3__q  $ (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__3__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__3__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__3__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__3__q ),
	.datab(!Xd_0__inst_product_27__3__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_24__3__q  $ (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_24__3__q  $ (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__3__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__3__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__3__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__3__q ),
	.datab(!Xd_0__inst_product_25__3__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_22__3__q  $ (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_22__3__q  $ (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__3__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__3__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__3__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__3__q ),
	.datab(!Xd_0__inst_product_23__3__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_20__3__q  $ (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_20__3__q  $ (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__3__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__3__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__3__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__3__q ),
	.datab(!Xd_0__inst_product_21__3__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_18__3__q  $ (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_18__3__q  $ (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__3__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__3__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__3__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__3__q ),
	.datab(!Xd_0__inst_product_19__3__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_16__4__q  $ (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_16__4__q  $ (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__4__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__4__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__4__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__4__q ),
	.datab(!Xd_0__inst_product_17__4__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_14__4__q  $ (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__4__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__4__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__4__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__4__q ),
	.datab(!Xd_0__inst_product_15__4__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_12__4__q  $ (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__4__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__4__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__4__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__4__q ),
	.datab(!Xd_0__inst_product_13__4__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_10__4__q  $ (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__4__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__4__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__4__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__4__q ),
	.datab(!Xd_0__inst_product_11__4__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_8__4__q  $ (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__4__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__4__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__4__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__4__q ),
	.datab(!Xd_0__inst_product_9__4__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__4__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__4__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__4__q ),
	.datab(!Xd_0__inst_product_7__4__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__4__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__4__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__4__q ),
	.datab(!Xd_0__inst_product_5__4__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__4__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__4__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__4__q ),
	.datab(!Xd_0__inst_product_3__4__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__4__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__4__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__4__q ),
	.datab(!Xd_0__inst_product_1__4__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_28__4__q  $ (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_28__4__q  $ (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__4__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__4__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__4__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__4__q ),
	.datab(!Xd_0__inst_product_29__4__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_26__4__q  $ (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_26__4__q  $ (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__4__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__4__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__4__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__4__q ),
	.datab(!Xd_0__inst_product_27__4__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_24__4__q  $ (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_24__4__q  $ (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__4__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__4__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__4__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__4__q ),
	.datab(!Xd_0__inst_product_25__4__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_22__4__q  $ (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_22__4__q  $ (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__4__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__4__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__4__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__4__q ),
	.datab(!Xd_0__inst_product_23__4__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_20__4__q  $ (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_20__4__q  $ (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__4__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__4__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__4__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__4__q ),
	.datab(!Xd_0__inst_product_21__4__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_18__4__q  $ (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_18__4__q  $ (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__4__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__4__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__4__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__4__q ),
	.datab(!Xd_0__inst_product_19__4__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_16__5__q  $ (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_16__5__q  $ (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__5__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__5__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__5__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__5__q ),
	.datab(!Xd_0__inst_product_17__5__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_14__5__q  $ (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__5__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__5__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__5__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__5__q ),
	.datab(!Xd_0__inst_product_15__5__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_12__5__q  $ (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__5__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__5__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__5__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__5__q ),
	.datab(!Xd_0__inst_product_13__5__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_10__5__q  $ (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__5__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__5__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__5__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__5__q ),
	.datab(!Xd_0__inst_product_11__5__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_8__5__q  $ (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__5__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__5__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__5__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__5__q ),
	.datab(!Xd_0__inst_product_9__5__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__5__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__5__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__5__q ),
	.datab(!Xd_0__inst_product_7__5__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__5__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__5__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__5__q ),
	.datab(!Xd_0__inst_product_5__5__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__5__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__5__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__5__q ),
	.datab(!Xd_0__inst_product_3__5__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__5__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__5__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__5__q ),
	.datab(!Xd_0__inst_product_1__5__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_28__5__q  $ (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_28__5__q  $ (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__5__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__5__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__5__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__5__q ),
	.datab(!Xd_0__inst_product_29__5__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_26__5__q  $ (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_26__5__q  $ (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__5__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__5__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__5__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__5__q ),
	.datab(!Xd_0__inst_product_27__5__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_24__5__q  $ (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_24__5__q  $ (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__5__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__5__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__5__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__5__q ),
	.datab(!Xd_0__inst_product_25__5__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_22__5__q  $ (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_22__5__q  $ (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__5__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__5__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__5__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__5__q ),
	.datab(!Xd_0__inst_product_23__5__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_20__5__q  $ (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_20__5__q  $ (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__5__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__5__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__5__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__5__q ),
	.datab(!Xd_0__inst_product_21__5__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_18__5__q  $ (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_18__5__q  $ (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__5__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__5__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__5__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__5__q ),
	.datab(!Xd_0__inst_product_19__5__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_16__6__q  $ (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_16__6__q  $ (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__6__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__6__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__6__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__6__q ),
	.datab(!Xd_0__inst_product_17__6__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_14__6__q  $ (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__6__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__6__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__6__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__6__q ),
	.datab(!Xd_0__inst_product_15__6__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_12__6__q  $ (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__6__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__6__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__6__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__6__q ),
	.datab(!Xd_0__inst_product_13__6__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_10__6__q  $ (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__6__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__6__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__6__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__6__q ),
	.datab(!Xd_0__inst_product_11__6__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_8__6__q  $ (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__6__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__6__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__6__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__6__q ),
	.datab(!Xd_0__inst_product_9__6__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__6__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__6__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__6__q ),
	.datab(!Xd_0__inst_product_7__6__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__6__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__6__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__6__q ),
	.datab(!Xd_0__inst_product_5__6__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__6__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__6__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__6__q ),
	.datab(!Xd_0__inst_product_3__6__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__6__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__6__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__6__q ),
	.datab(!Xd_0__inst_product_1__6__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_28__6__q  $ (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_28__6__q  $ (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__6__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__6__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__6__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__6__q ),
	.datab(!Xd_0__inst_product_29__6__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_26__6__q  $ (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_26__6__q  $ (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__6__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__6__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__6__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__6__q ),
	.datab(!Xd_0__inst_product_27__6__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_24__6__q  $ (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_24__6__q  $ (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__6__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__6__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__6__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__6__q ),
	.datab(!Xd_0__inst_product_25__6__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_22__6__q  $ (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_22__6__q  $ (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__6__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__6__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__6__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__6__q ),
	.datab(!Xd_0__inst_product_23__6__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_20__6__q  $ (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_20__6__q  $ (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__6__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__6__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__6__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__6__q ),
	.datab(!Xd_0__inst_product_21__6__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_18__6__q  $ (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_18__6__q  $ (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__6__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__6__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__6__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__6__q ),
	.datab(!Xd_0__inst_product_19__6__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_16__7__q  $ (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_16__7__q  $ (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__7__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__7__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__7__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__7__q ),
	.datab(!Xd_0__inst_product_17__7__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_14__7__q  $ (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__7__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__7__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__7__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__7__q ),
	.datab(!Xd_0__inst_product_15__7__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_12__7__q  $ (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__7__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__7__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__7__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__7__q ),
	.datab(!Xd_0__inst_product_13__7__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_10__7__q  $ (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__7__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__7__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__7__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__7__q ),
	.datab(!Xd_0__inst_product_11__7__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_8__7__q  $ (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__7__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__7__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__7__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__7__q ),
	.datab(!Xd_0__inst_product_9__7__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__7__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__7__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__7__q ),
	.datab(!Xd_0__inst_product_7__7__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__7__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__7__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__7__q ),
	.datab(!Xd_0__inst_product_5__7__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__7__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__7__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__7__q ),
	.datab(!Xd_0__inst_product_3__7__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__7__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__7__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__7__q ),
	.datab(!Xd_0__inst_product_1__7__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_28__7__q  $ (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_28__7__q  $ (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__7__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__7__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__7__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__7__q ),
	.datab(!Xd_0__inst_product_29__7__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_26__7__q  $ (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_26__7__q  $ (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__7__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__7__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__7__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__7__q ),
	.datab(!Xd_0__inst_product_27__7__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_24__7__q  $ (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_24__7__q  $ (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__7__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__7__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__7__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__7__q ),
	.datab(!Xd_0__inst_product_25__7__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_22__7__q  $ (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_22__7__q  $ (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__7__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__7__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__7__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__7__q ),
	.datab(!Xd_0__inst_product_23__7__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_20__7__q  $ (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_20__7__q  $ (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__7__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__7__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__7__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__7__q ),
	.datab(!Xd_0__inst_product_21__7__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_18__7__q  $ (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_18__7__q  $ (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__7__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__7__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__7__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__7__q ),
	.datab(!Xd_0__inst_product_19__7__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_16__8__q  $ (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_16__8__q  $ (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__8__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__8__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__8__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__8__q ),
	.datab(!Xd_0__inst_product_17__8__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_14__8__q  $ (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__8__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__8__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__8__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__8__q ),
	.datab(!Xd_0__inst_product_15__8__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_12__8__q  $ (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__8__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__8__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__8__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__8__q ),
	.datab(!Xd_0__inst_product_13__8__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_10__8__q  $ (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__8__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__8__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__8__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__8__q ),
	.datab(!Xd_0__inst_product_11__8__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_8__8__q  $ (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__8__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__8__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__8__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__8__q ),
	.datab(!Xd_0__inst_product_9__8__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__8__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__8__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__8__q ),
	.datab(!Xd_0__inst_product_7__8__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__8__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__8__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__8__q ),
	.datab(!Xd_0__inst_product_5__8__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__8__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__8__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__8__q ),
	.datab(!Xd_0__inst_product_3__8__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__8__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__8__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__8__q ),
	.datab(!Xd_0__inst_product_1__8__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_28__8__q  $ (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_28__8__q  $ (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__8__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__8__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__8__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__8__q ),
	.datab(!Xd_0__inst_product_29__8__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_26__8__q  $ (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_26__8__q  $ (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__8__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__8__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__8__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__8__q ),
	.datab(!Xd_0__inst_product_27__8__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_24__8__q  $ (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_24__8__q  $ (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__8__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__8__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__8__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__8__q ),
	.datab(!Xd_0__inst_product_25__8__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_22__8__q  $ (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_22__8__q  $ (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__8__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__8__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__8__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__8__q ),
	.datab(!Xd_0__inst_product_23__8__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_20__8__q  $ (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_20__8__q  $ (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__8__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__8__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__8__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__8__q ),
	.datab(!Xd_0__inst_product_21__8__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_18__8__q  $ (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_18__8__q  $ (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__8__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__8__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__8__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__8__q ),
	.datab(!Xd_0__inst_product_19__8__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_16__9__q  $ (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_16__9__q  $ (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]))) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_16__9__q  & (Xd_0__inst_sign [16] & (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [17])))) # (Xd_0__inst_product_16__9__q  & (!Xd_0__inst_sign [16] & 
// (!Xd_0__inst_product_17__9__q  $ (!Xd_0__inst_sign [17])))))

	.dataa(!Xd_0__inst_product_16__9__q ),
	.datab(!Xd_0__inst_product_17__9__q ),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_14__9__q  $ (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]))) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_14__9__q  & (Xd_0__inst_sign [14] & (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))) # (Xd_0__inst_product_14__9__q  & (!Xd_0__inst_sign [14] & 
// (!Xd_0__inst_product_15__9__q  $ (!Xd_0__inst_sign [15])))))

	.dataa(!Xd_0__inst_product_14__9__q ),
	.datab(!Xd_0__inst_product_15__9__q ),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_12__9__q  $ (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]))) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_12__9__q  & (Xd_0__inst_sign [12] & (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))) # (Xd_0__inst_product_12__9__q  & (!Xd_0__inst_sign [12] & 
// (!Xd_0__inst_product_13__9__q  $ (!Xd_0__inst_sign [13])))))

	.dataa(!Xd_0__inst_product_12__9__q ),
	.datab(!Xd_0__inst_product_13__9__q ),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_10__9__q  $ (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]))) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_10__9__q  & (Xd_0__inst_sign [10] & (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))) # (Xd_0__inst_product_10__9__q  & (!Xd_0__inst_sign [10] & 
// (!Xd_0__inst_product_11__9__q  $ (!Xd_0__inst_sign [11])))))

	.dataa(!Xd_0__inst_product_10__9__q ),
	.datab(!Xd_0__inst_product_11__9__q ),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_8__9__q  $ (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]))) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_8__9__q  & (Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q  $ (!Xd_0__inst_sign [9])))) # (Xd_0__inst_product_8__9__q  & (!Xd_0__inst_sign [8] & (!Xd_0__inst_product_9__9__q 
//  $ (!Xd_0__inst_sign [9])))))

	.dataa(!Xd_0__inst_product_8__9__q ),
	.datab(!Xd_0__inst_product_9__9__q ),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__9__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__9__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__9__q ),
	.datab(!Xd_0__inst_product_7__9__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__9__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__9__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__9__q ),
	.datab(!Xd_0__inst_product_5__9__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__9__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__9__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__9__q ),
	.datab(!Xd_0__inst_product_3__9__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__9__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__9__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__9__q ),
	.datab(!Xd_0__inst_product_1__9__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_28__9__q  $ (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_28__9__q  $ (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]))) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_28__9__q  & (Xd_0__inst_sign [28] & (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [29])))) # (Xd_0__inst_product_28__9__q  & (!Xd_0__inst_sign [28] & 
// (!Xd_0__inst_product_29__9__q  $ (!Xd_0__inst_sign [29])))))

	.dataa(!Xd_0__inst_product_28__9__q ),
	.datab(!Xd_0__inst_product_29__9__q ),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_26__9__q  $ (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_26__9__q  $ (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]))) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_26__9__q  & (Xd_0__inst_sign [26] & (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [27])))) # (Xd_0__inst_product_26__9__q  & (!Xd_0__inst_sign [26] & 
// (!Xd_0__inst_product_27__9__q  $ (!Xd_0__inst_sign [27])))))

	.dataa(!Xd_0__inst_product_26__9__q ),
	.datab(!Xd_0__inst_product_27__9__q ),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_24__9__q  $ (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_24__9__q  $ (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]))) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_24__9__q  & (Xd_0__inst_sign [24] & (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [25])))) # (Xd_0__inst_product_24__9__q  & (!Xd_0__inst_sign [24] & 
// (!Xd_0__inst_product_25__9__q  $ (!Xd_0__inst_sign [25])))))

	.dataa(!Xd_0__inst_product_24__9__q ),
	.datab(!Xd_0__inst_product_25__9__q ),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_22__9__q  $ (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_22__9__q  $ (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]))) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_22__9__q  & (Xd_0__inst_sign [22] & (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [23])))) # (Xd_0__inst_product_22__9__q  & (!Xd_0__inst_sign [22] & 
// (!Xd_0__inst_product_23__9__q  $ (!Xd_0__inst_sign [23])))))

	.dataa(!Xd_0__inst_product_22__9__q ),
	.datab(!Xd_0__inst_product_23__9__q ),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_20__9__q  $ (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_20__9__q  $ (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]))) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_20__9__q  & (Xd_0__inst_sign [20] & (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [21])))) # (Xd_0__inst_product_20__9__q  & (!Xd_0__inst_sign [20] & 
// (!Xd_0__inst_product_21__9__q  $ (!Xd_0__inst_sign [21])))))

	.dataa(!Xd_0__inst_product_20__9__q ),
	.datab(!Xd_0__inst_product_21__9__q ),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_18__9__q  $ (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_18__9__q  $ (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]))) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_18__9__q  & (Xd_0__inst_sign [18] & (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [19])))) # (Xd_0__inst_product_18__9__q  & (!Xd_0__inst_sign [18] & 
// (!Xd_0__inst_product_19__9__q  $ (!Xd_0__inst_sign [19])))))

	.dataa(!Xd_0__inst_product_18__9__q ),
	.datab(!Xd_0__inst_product_19__9__q ),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_8__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_8__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [16] & Xd_0__inst_sign [17]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [16]),
	.datad(!Xd_0__inst_sign [17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_8__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_7__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_7__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [14] & Xd_0__inst_sign [15]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [14]),
	.datad(!Xd_0__inst_sign [15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_6__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_6__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [12] & Xd_0__inst_sign [13]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [12]),
	.datad(!Xd_0__inst_sign [13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_5__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_5__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [10] & Xd_0__inst_sign [11]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [10]),
	.datad(!Xd_0__inst_sign [11]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_4__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_4__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [8] & Xd_0__inst_sign [9]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [8]),
	.datad(!Xd_0__inst_sign [9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [6] & Xd_0__inst_sign [7]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [4] & Xd_0__inst_sign [5]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [2] & Xd_0__inst_sign [3]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [0] & Xd_0__inst_sign [1]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_14__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_14__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [28] & Xd_0__inst_sign [29]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [28]),
	.datad(!Xd_0__inst_sign [29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_14__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_13__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_13__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [26] & Xd_0__inst_sign [27]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [26]),
	.datad(!Xd_0__inst_sign [27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_13__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_12__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_12__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [24] & Xd_0__inst_sign [25]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [24]),
	.datad(!Xd_0__inst_sign [25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_12__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_11__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_11__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [22] & Xd_0__inst_sign [23]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [22]),
	.datad(!Xd_0__inst_sign [23]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_11__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_10__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_10__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [20] & Xd_0__inst_sign [21]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [20]),
	.datad(!Xd_0__inst_sign [21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_10__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_9__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_9__adder1_inst_dout [10] = SUM(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [18] & Xd_0__inst_sign [19]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [18]),
	.datad(!Xd_0__inst_sign [19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_9__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_34 (
// Equation(s):
// Xd_0__inst_mult_0_35  = SUM(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_0_36  = CARRY(( !Xd_0__inst_sign [16] $ (!Xd_0__inst_sign [17]) ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_8__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_0_37  = SHARE((Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_1_q ))

	.dataa(!Xd_0__inst_sign [16]),
	.datab(!Xd_0__inst_sign [17]),
	.datac(!Xd_0__inst_mult_0_0_q ),
	.datad(!Xd_0__inst_mult_0_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_8__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_8__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_35 ),
	.cout(Xd_0__inst_mult_0_36 ),
	.shareout(Xd_0__inst_mult_0_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_25_35 (
// Equation(s):
// Xd_0__inst_mult_25_36  = SUM(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_25_37  = CARRY(( !Xd_0__inst_sign [14] $ (!Xd_0__inst_sign [15]) ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_7__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_25_38  = SHARE((Xd_0__inst_mult_25_0_q  & Xd_0__inst_mult_25_1_q ))

	.dataa(!Xd_0__inst_sign [14]),
	.datab(!Xd_0__inst_sign [15]),
	.datac(!Xd_0__inst_mult_25_0_q ),
	.datad(!Xd_0__inst_mult_25_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_7__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_7__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_36 ),
	.cout(Xd_0__inst_mult_25_37 ),
	.shareout(Xd_0__inst_mult_25_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_24_17 (
// Equation(s):
// Xd_0__inst_mult_24_47  = SUM(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_24_48  = CARRY(( !Xd_0__inst_sign [12] $ (!Xd_0__inst_sign [13]) ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_6__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_24_49  = SHARE((Xd_0__inst_mult_24_0_q  & Xd_0__inst_mult_24_1_q ))

	.dataa(!Xd_0__inst_sign [12]),
	.datab(!Xd_0__inst_sign [13]),
	.datac(!Xd_0__inst_mult_24_0_q ),
	.datad(!Xd_0__inst_mult_24_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_6__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_6__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_47 ),
	.cout(Xd_0__inst_mult_24_48 ),
	.shareout(Xd_0__inst_mult_24_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_27_35 (
// Equation(s):
// Xd_0__inst_mult_27_36  = SUM(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_27_37  = CARRY(( !Xd_0__inst_sign [10] $ (!Xd_0__inst_sign [11]) ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_5__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_27_38  = SHARE((Xd_0__inst_mult_27_0_q  & Xd_0__inst_mult_27_1_q ))

	.dataa(!Xd_0__inst_sign [10]),
	.datab(!Xd_0__inst_sign [11]),
	.datac(!Xd_0__inst_mult_27_0_q ),
	.datad(!Xd_0__inst_mult_27_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_5__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_5__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_36 ),
	.cout(Xd_0__inst_mult_27_37 ),
	.shareout(Xd_0__inst_mult_27_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_26_16 (
// Equation(s):
// Xd_0__inst_mult_26_43  = SUM(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_26_44  = CARRY(( !Xd_0__inst_sign [8] $ (!Xd_0__inst_sign [9]) ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_4__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_26_45  = SHARE((Xd_0__inst_mult_26_0_q  & Xd_0__inst_mult_26_1_q ))

	.dataa(!Xd_0__inst_sign [8]),
	.datab(!Xd_0__inst_sign [9]),
	.datac(!Xd_0__inst_mult_26_0_q ),
	.datad(!Xd_0__inst_mult_26_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_4__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_4__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_43 ),
	.cout(Xd_0__inst_mult_26_44 ),
	.shareout(Xd_0__inst_mult_26_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_29_35 (
// Equation(s):
// Xd_0__inst_mult_29_36  = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_29_37  = CARRY(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_29_38  = SHARE((Xd_0__inst_mult_29_0_q  & Xd_0__inst_mult_29_1_q ))

	.dataa(!Xd_0__inst_sign [6]),
	.datab(!Xd_0__inst_sign [7]),
	.datac(!Xd_0__inst_mult_29_0_q ),
	.datad(!Xd_0__inst_mult_29_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_36 ),
	.cout(Xd_0__inst_mult_29_37 ),
	.shareout(Xd_0__inst_mult_29_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_28_16 (
// Equation(s):
// Xd_0__inst_mult_28_43  = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_28_44  = CARRY(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_28_45  = SHARE((Xd_0__inst_mult_28_0_q  & Xd_0__inst_mult_28_1_q ))

	.dataa(!Xd_0__inst_sign [4]),
	.datab(!Xd_0__inst_sign [5]),
	.datac(!Xd_0__inst_mult_28_0_q ),
	.datad(!Xd_0__inst_mult_28_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_43 ),
	.cout(Xd_0__inst_mult_28_44 ),
	.shareout(Xd_0__inst_mult_28_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_31_35 (
// Equation(s):
// Xd_0__inst_mult_31_36  = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_31_37  = CARRY(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_31_38  = SHARE((Xd_0__inst_mult_31_0_q  & Xd_0__inst_mult_31_1_q ))

	.dataa(!Xd_0__inst_sign [2]),
	.datab(!Xd_0__inst_sign [3]),
	.datac(!Xd_0__inst_mult_31_0_q ),
	.datad(!Xd_0__inst_mult_31_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_36 ),
	.cout(Xd_0__inst_mult_31_37 ),
	.shareout(Xd_0__inst_mult_31_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_20_17 (
// Equation(s):
// Xd_0__inst_mult_20_47  = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_20_48  = CARRY(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_20_49  = SHARE((Xd_0__inst_mult_20_0_q  & Xd_0__inst_mult_20_1_q ))

	.dataa(!Xd_0__inst_sign [0]),
	.datab(!Xd_0__inst_sign [1]),
	.datac(!Xd_0__inst_mult_20_0_q ),
	.datad(!Xd_0__inst_mult_20_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_47 ),
	.cout(Xd_0__inst_mult_20_48 ),
	.shareout(Xd_0__inst_mult_20_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_34 (
// Equation(s):
// Xd_0__inst_mult_3_35  = SUM(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_3_36  = CARRY(( !Xd_0__inst_sign [28] $ (!Xd_0__inst_sign [29]) ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_14__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_3_37  = SHARE((Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_1_q ))

	.dataa(!Xd_0__inst_sign [28]),
	.datab(!Xd_0__inst_sign [29]),
	.datac(!Xd_0__inst_mult_3_0_q ),
	.datad(!Xd_0__inst_mult_3_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_14__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_14__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_35 ),
	.cout(Xd_0__inst_mult_3_36 ),
	.shareout(Xd_0__inst_mult_3_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_34 (
// Equation(s):
// Xd_0__inst_mult_1_35  = SUM(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_1_36  = CARRY(( !Xd_0__inst_sign [26] $ (!Xd_0__inst_sign [27]) ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_13__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_1_37  = SHARE((Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_1_q ))

	.dataa(!Xd_0__inst_sign [26]),
	.datab(!Xd_0__inst_sign [27]),
	.datac(!Xd_0__inst_mult_1_0_q ),
	.datad(!Xd_0__inst_mult_1_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_13__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_13__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_35 ),
	.cout(Xd_0__inst_mult_1_36 ),
	.shareout(Xd_0__inst_mult_1_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_35 (
// Equation(s):
// Xd_0__inst_mult_11_36  = SUM(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_11_37  = CARRY(( !Xd_0__inst_sign [24] $ (!Xd_0__inst_sign [25]) ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_12__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_11_38  = SHARE((Xd_0__inst_mult_11_0_q  & Xd_0__inst_mult_11_1_q ))

	.dataa(!Xd_0__inst_sign [24]),
	.datab(!Xd_0__inst_sign [25]),
	.datac(!Xd_0__inst_mult_11_0_q ),
	.datad(!Xd_0__inst_mult_11_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_12__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_12__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_36 ),
	.cout(Xd_0__inst_mult_11_37 ),
	.shareout(Xd_0__inst_mult_11_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_30_16 (
// Equation(s):
// Xd_0__inst_mult_30_43  = SUM(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_30_44  = CARRY(( !Xd_0__inst_sign [22] $ (!Xd_0__inst_sign [23]) ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_11__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_30_45  = SHARE((Xd_0__inst_mult_30_0_q  & Xd_0__inst_mult_30_1_q ))

	.dataa(!Xd_0__inst_sign [22]),
	.datab(!Xd_0__inst_sign [23]),
	.datac(!Xd_0__inst_mult_30_0_q ),
	.datad(!Xd_0__inst_mult_30_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_11__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_11__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_43 ),
	.cout(Xd_0__inst_mult_30_44 ),
	.shareout(Xd_0__inst_mult_30_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_23_17 (
// Equation(s):
// Xd_0__inst_mult_23_47  = SUM(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_23_48  = CARRY(( !Xd_0__inst_sign [20] $ (!Xd_0__inst_sign [21]) ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_10__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_23_49  = SHARE((Xd_0__inst_mult_23_0_q  & Xd_0__inst_mult_23_1_q ))

	.dataa(!Xd_0__inst_sign [20]),
	.datab(!Xd_0__inst_sign [21]),
	.datac(!Xd_0__inst_mult_23_0_q ),
	.datad(!Xd_0__inst_mult_23_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_10__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_10__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_47 ),
	.cout(Xd_0__inst_mult_23_48 ),
	.shareout(Xd_0__inst_mult_23_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00006666),
	.shared_arith("on")
) Xd_0__inst_mult_22_16 (
// Equation(s):
// Xd_0__inst_mult_22_43  = SUM(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_22_44  = CARRY(( !Xd_0__inst_sign [18] $ (!Xd_0__inst_sign [19]) ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_9__adder1_inst_wc_n_COUT  ))
// Xd_0__inst_mult_22_45  = SHARE((Xd_0__inst_mult_22_0_q  & Xd_0__inst_mult_22_1_q ))

	.dataa(!Xd_0__inst_sign [18]),
	.datab(!Xd_0__inst_sign [19]),
	.datac(!Xd_0__inst_mult_22_0_q ),
	.datad(!Xd_0__inst_mult_22_1_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_9__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_9__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_43 ),
	.cout(Xd_0__inst_mult_22_44 ),
	.shareout(Xd_0__inst_mult_22_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_17 (
// Equation(s):
// Xd_0__inst_mult_26_48  = CARRY(( GND ) + ( Xd_0__inst_mult_29_42  ) + ( Xd_0__inst_mult_29_41  ))
// Xd_0__inst_mult_26_49  = SHARE((din_b[159] & din_a[157]))

	.dataa(!din_b[159]),
	.datab(!din_a[157]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_41 ),
	.sharein(Xd_0__inst_mult_29_42 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_48 ),
	.shareout(Xd_0__inst_mult_26_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_17 (
// Equation(s):
// Xd_0__inst_mult_28_48  = CARRY(( GND ) + ( Xd_0__inst_mult_31_69  ) + ( Xd_0__inst_mult_31_68  ))
// Xd_0__inst_mult_28_49  = SHARE((din_b[171] & din_a[169]))

	.dataa(!din_b[171]),
	.datab(!din_a[169]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_68 ),
	.sharein(Xd_0__inst_mult_31_69 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_48 ),
	.shareout(Xd_0__inst_mult_28_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_17 (
// Equation(s):
// Xd_0__inst_mult_30_48  = CARRY(( GND ) + ( Xd_0__inst_mult_11_42  ) + ( Xd_0__inst_mult_11_41  ))
// Xd_0__inst_mult_30_49  = SHARE((din_b[183] & din_a[181]))

	.dataa(!din_b[183]),
	.datab(!din_a[181]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_41 ),
	.sharein(Xd_0__inst_mult_11_42 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_48 ),
	.shareout(Xd_0__inst_mult_30_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_17 (
// Equation(s):
// Xd_0__inst_mult_22_48  = CARRY(( GND ) + ( Xd_0__inst_mult_25_42  ) + ( Xd_0__inst_mult_25_41  ))
// Xd_0__inst_mult_22_49  = SHARE((din_b[135] & din_a[133]))

	.dataa(!din_b[135]),
	.datab(!din_a[133]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_41 ),
	.sharein(Xd_0__inst_mult_25_42 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_48 ),
	.shareout(Xd_0__inst_mult_22_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_16 (
// Equation(s):
// Xd_0__inst_mult_19_44  = CARRY(( GND ) + ( Xd_0__inst_mult_27_42  ) + ( Xd_0__inst_mult_27_41  ))
// Xd_0__inst_mult_19_45  = SHARE((din_b[117] & din_a[115]))

	.dataa(!din_b[117]),
	.datab(!din_a[115]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_41 ),
	.sharein(Xd_0__inst_mult_27_42 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_44 ),
	.shareout(Xd_0__inst_mult_19_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_30_18 (
// Equation(s):
// Xd_0__inst_mult_30_51  = SUM(( Xd_0__inst_mult_30_5_q  ) + ( Xd_0__inst_mult_30_93  ) + ( Xd_0__inst_mult_30_92  ))
// Xd_0__inst_mult_30_52  = CARRY(( Xd_0__inst_mult_30_5_q  ) + ( Xd_0__inst_mult_30_93  ) + ( Xd_0__inst_mult_30_92  ))
// Xd_0__inst_mult_30_53  = SHARE((Xd_0__inst_mult_30_4_q  & Xd_0__inst_mult_30_2_q ))

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_2_q ),
	.datac(!Xd_0__inst_mult_30_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_92 ),
	.sharein(Xd_0__inst_mult_30_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_51 ),
	.cout(Xd_0__inst_mult_30_52 ),
	.shareout(Xd_0__inst_mult_30_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_31 (
// Equation(s):
// Xd_0__inst_mult_31_40  = SUM(( Xd_0__inst_mult_31_5_q  ) + ( Xd_0__inst_mult_31_85  ) + ( Xd_0__inst_mult_31_84  ))
// Xd_0__inst_mult_31_41  = CARRY(( Xd_0__inst_mult_31_5_q  ) + ( Xd_0__inst_mult_31_85  ) + ( Xd_0__inst_mult_31_84  ))
// Xd_0__inst_mult_31_42  = SHARE((Xd_0__inst_mult_31_4_q  & Xd_0__inst_mult_31_2_q ))

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_2_q ),
	.datac(!Xd_0__inst_mult_31_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_84 ),
	.sharein(Xd_0__inst_mult_31_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_40 ),
	.cout(Xd_0__inst_mult_31_41 ),
	.shareout(Xd_0__inst_mult_31_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_30_19 (
// Equation(s):
// Xd_0__inst_mult_30_55  = SUM(( !Xd_0__inst_mult_30_6_q  $ (!Xd_0__inst_mult_30_7_q ) ) + ( Xd_0__inst_mult_30_53  ) + ( Xd_0__inst_mult_30_52  ))
// Xd_0__inst_mult_30_56  = CARRY(( !Xd_0__inst_mult_30_6_q  $ (!Xd_0__inst_mult_30_7_q ) ) + ( Xd_0__inst_mult_30_53  ) + ( Xd_0__inst_mult_30_52  ))
// Xd_0__inst_mult_30_57  = SHARE((Xd_0__inst_mult_30_6_q  & Xd_0__inst_mult_30_7_q ))

	.dataa(!Xd_0__inst_mult_30_6_q ),
	.datab(!Xd_0__inst_mult_30_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_52 ),
	.sharein(Xd_0__inst_mult_30_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_55 ),
	.cout(Xd_0__inst_mult_30_56 ),
	.shareout(Xd_0__inst_mult_30_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_31_16 (
// Equation(s):
// Xd_0__inst_mult_31_43  = SUM(( !Xd_0__inst_mult_31_6_q  $ (!Xd_0__inst_mult_31_7_q ) ) + ( Xd_0__inst_mult_31_42  ) + ( Xd_0__inst_mult_31_41  ))
// Xd_0__inst_mult_31_44  = CARRY(( !Xd_0__inst_mult_31_6_q  $ (!Xd_0__inst_mult_31_7_q ) ) + ( Xd_0__inst_mult_31_42  ) + ( Xd_0__inst_mult_31_41  ))
// Xd_0__inst_mult_31_45  = SHARE((Xd_0__inst_mult_31_6_q  & Xd_0__inst_mult_31_7_q ))

	.dataa(!Xd_0__inst_mult_31_6_q ),
	.datab(!Xd_0__inst_mult_31_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_41 ),
	.sharein(Xd_0__inst_mult_31_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_43 ),
	.cout(Xd_0__inst_mult_31_44 ),
	.shareout(Xd_0__inst_mult_31_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_30_20 (
// Equation(s):
// Xd_0__inst_mult_30_59  = SUM(( !Xd_0__inst_mult_30_8_q  $ (!Xd_0__inst_mult_30_9_q  $ (((Xd_0__inst_mult_30_4_q  & Xd_0__inst_mult_30_10_q )))) ) + ( Xd_0__inst_mult_30_57  ) + ( Xd_0__inst_mult_30_56  ))
// Xd_0__inst_mult_30_60  = CARRY(( !Xd_0__inst_mult_30_8_q  $ (!Xd_0__inst_mult_30_9_q  $ (((Xd_0__inst_mult_30_4_q  & Xd_0__inst_mult_30_10_q )))) ) + ( Xd_0__inst_mult_30_57  ) + ( Xd_0__inst_mult_30_56  ))
// Xd_0__inst_mult_30_61  = SHARE((!Xd_0__inst_mult_30_8_q  & (Xd_0__inst_mult_30_9_q  & (Xd_0__inst_mult_30_4_q  & Xd_0__inst_mult_30_10_q ))) # (Xd_0__inst_mult_30_8_q  & (((Xd_0__inst_mult_30_4_q  & Xd_0__inst_mult_30_10_q )) # (Xd_0__inst_mult_30_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_30_8_q ),
	.datab(!Xd_0__inst_mult_30_9_q ),
	.datac(!Xd_0__inst_mult_30_4_q ),
	.datad(!Xd_0__inst_mult_30_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_56 ),
	.sharein(Xd_0__inst_mult_30_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_59 ),
	.cout(Xd_0__inst_mult_30_60 ),
	.shareout(Xd_0__inst_mult_30_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_31_17 (
// Equation(s):
// Xd_0__inst_mult_31_47  = SUM(( !Xd_0__inst_mult_31_8_q  $ (!Xd_0__inst_mult_31_9_q  $ (((Xd_0__inst_mult_31_4_q  & Xd_0__inst_mult_31_10_q )))) ) + ( Xd_0__inst_mult_31_45  ) + ( Xd_0__inst_mult_31_44  ))
// Xd_0__inst_mult_31_48  = CARRY(( !Xd_0__inst_mult_31_8_q  $ (!Xd_0__inst_mult_31_9_q  $ (((Xd_0__inst_mult_31_4_q  & Xd_0__inst_mult_31_10_q )))) ) + ( Xd_0__inst_mult_31_45  ) + ( Xd_0__inst_mult_31_44  ))
// Xd_0__inst_mult_31_49  = SHARE((!Xd_0__inst_mult_31_8_q  & (Xd_0__inst_mult_31_9_q  & (Xd_0__inst_mult_31_4_q  & Xd_0__inst_mult_31_10_q ))) # (Xd_0__inst_mult_31_8_q  & (((Xd_0__inst_mult_31_4_q  & Xd_0__inst_mult_31_10_q )) # (Xd_0__inst_mult_31_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_31_8_q ),
	.datab(!Xd_0__inst_mult_31_9_q ),
	.datac(!Xd_0__inst_mult_31_4_q ),
	.datad(!Xd_0__inst_mult_31_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_44 ),
	.sharein(Xd_0__inst_mult_31_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_47 ),
	.cout(Xd_0__inst_mult_31_48 ),
	.shareout(Xd_0__inst_mult_31_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_30_21 (
// Equation(s):
// Xd_0__inst_mult_30_63  = SUM(( !Xd_0__inst_mult_30_12_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_11_q ))) ) + ( Xd_0__inst_mult_30_61  ) + ( Xd_0__inst_mult_30_60  ))
// Xd_0__inst_mult_30_64  = CARRY(( !Xd_0__inst_mult_30_12_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_11_q ))) ) + ( Xd_0__inst_mult_30_61  ) + ( Xd_0__inst_mult_30_60  ))
// Xd_0__inst_mult_30_65  = SHARE((Xd_0__inst_mult_30_4_q  & (Xd_0__inst_mult_30_11_q  & Xd_0__inst_mult_30_12_q )))

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_11_q ),
	.datac(!Xd_0__inst_mult_30_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_60 ),
	.sharein(Xd_0__inst_mult_30_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_63 ),
	.cout(Xd_0__inst_mult_30_64 ),
	.shareout(Xd_0__inst_mult_30_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_31_18 (
// Equation(s):
// Xd_0__inst_mult_31_51  = SUM(( !Xd_0__inst_mult_31_12_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_11_q ))) ) + ( Xd_0__inst_mult_31_49  ) + ( Xd_0__inst_mult_31_48  ))
// Xd_0__inst_mult_31_52  = CARRY(( !Xd_0__inst_mult_31_12_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_11_q ))) ) + ( Xd_0__inst_mult_31_49  ) + ( Xd_0__inst_mult_31_48  ))
// Xd_0__inst_mult_31_53  = SHARE((Xd_0__inst_mult_31_4_q  & (Xd_0__inst_mult_31_11_q  & Xd_0__inst_mult_31_12_q )))

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_11_q ),
	.datac(!Xd_0__inst_mult_31_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_48 ),
	.sharein(Xd_0__inst_mult_31_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_51 ),
	.cout(Xd_0__inst_mult_31_52 ),
	.shareout(Xd_0__inst_mult_31_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_30_22 (
// Equation(s):
// Xd_0__inst_mult_30_67  = SUM(( !Xd_0__inst_mult_30_13_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_0_q ))) ) + ( Xd_0__inst_mult_30_65  ) + ( Xd_0__inst_mult_30_64  ))
// Xd_0__inst_mult_30_68  = CARRY(( !Xd_0__inst_mult_30_13_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_0_q ))) ) + ( Xd_0__inst_mult_30_65  ) + ( Xd_0__inst_mult_30_64  ))
// Xd_0__inst_mult_30_69  = SHARE((Xd_0__inst_mult_30_4_q  & (Xd_0__inst_mult_30_0_q  & Xd_0__inst_mult_30_13_q )))

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_0_q ),
	.datac(!Xd_0__inst_mult_30_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_64 ),
	.sharein(Xd_0__inst_mult_30_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_67 ),
	.cout(Xd_0__inst_mult_30_68 ),
	.shareout(Xd_0__inst_mult_30_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_31_19 (
// Equation(s):
// Xd_0__inst_mult_31_55  = SUM(( !Xd_0__inst_mult_31_13_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_0_q ))) ) + ( Xd_0__inst_mult_31_53  ) + ( Xd_0__inst_mult_31_52  ))
// Xd_0__inst_mult_31_56  = CARRY(( !Xd_0__inst_mult_31_13_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_0_q ))) ) + ( Xd_0__inst_mult_31_53  ) + ( Xd_0__inst_mult_31_52  ))
// Xd_0__inst_mult_31_57  = SHARE((Xd_0__inst_mult_31_4_q  & (Xd_0__inst_mult_31_0_q  & Xd_0__inst_mult_31_13_q )))

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_0_q ),
	.datac(!Xd_0__inst_mult_31_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_52 ),
	.sharein(Xd_0__inst_mult_31_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_55 ),
	.cout(Xd_0__inst_mult_31_56 ),
	.shareout(Xd_0__inst_mult_31_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_30_23 (
// Equation(s):
// Xd_0__inst_mult_30_71  = SUM(( !Xd_0__inst_mult_30_15_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_14_q ))) ) + ( Xd_0__inst_mult_30_69  ) + ( Xd_0__inst_mult_30_68  ))
// Xd_0__inst_mult_30_72  = CARRY(( !Xd_0__inst_mult_30_15_q  $ (((!Xd_0__inst_mult_30_4_q ) # (!Xd_0__inst_mult_30_14_q ))) ) + ( Xd_0__inst_mult_30_69  ) + ( Xd_0__inst_mult_30_68  ))
// Xd_0__inst_mult_30_73  = SHARE((Xd_0__inst_mult_30_4_q  & (Xd_0__inst_mult_30_14_q  & Xd_0__inst_mult_30_15_q )))

	.dataa(!Xd_0__inst_mult_30_4_q ),
	.datab(!Xd_0__inst_mult_30_14_q ),
	.datac(!Xd_0__inst_mult_30_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_68 ),
	.sharein(Xd_0__inst_mult_30_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_71 ),
	.cout(Xd_0__inst_mult_30_72 ),
	.shareout(Xd_0__inst_mult_30_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_31_20 (
// Equation(s):
// Xd_0__inst_mult_31_59  = SUM(( !Xd_0__inst_mult_31_15_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_14_q ))) ) + ( Xd_0__inst_mult_31_57  ) + ( Xd_0__inst_mult_31_56  ))
// Xd_0__inst_mult_31_60  = CARRY(( !Xd_0__inst_mult_31_15_q  $ (((!Xd_0__inst_mult_31_4_q ) # (!Xd_0__inst_mult_31_14_q ))) ) + ( Xd_0__inst_mult_31_57  ) + ( Xd_0__inst_mult_31_56  ))
// Xd_0__inst_mult_31_61  = SHARE((Xd_0__inst_mult_31_4_q  & (Xd_0__inst_mult_31_14_q  & Xd_0__inst_mult_31_15_q )))

	.dataa(!Xd_0__inst_mult_31_4_q ),
	.datab(!Xd_0__inst_mult_31_14_q ),
	.datac(!Xd_0__inst_mult_31_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_56 ),
	.sharein(Xd_0__inst_mult_31_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_59 ),
	.cout(Xd_0__inst_mult_31_60 ),
	.shareout(Xd_0__inst_mult_31_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_24 (
// Equation(s):
// Xd_0__inst_mult_30_75  = SUM(( GND ) + ( Xd_0__inst_mult_30_73  ) + ( Xd_0__inst_mult_30_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_72 ),
	.sharein(Xd_0__inst_mult_30_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_21 (
// Equation(s):
// Xd_0__inst_mult_31_63  = SUM(( GND ) + ( Xd_0__inst_mult_31_61  ) + ( Xd_0__inst_mult_31_60  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_60 ),
	.sharein(Xd_0__inst_mult_31_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29 (
// Equation(s):
// Xd_0__inst_mult_29_40  = SUM(( GND ) + ( Xd_0__inst_mult_29_73  ) + ( Xd_0__inst_mult_29_72  ))
// Xd_0__inst_mult_29_41  = CARRY(( GND ) + ( Xd_0__inst_mult_29_73  ) + ( Xd_0__inst_mult_29_72  ))
// Xd_0__inst_mult_29_42  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_72 ),
	.sharein(Xd_0__inst_mult_29_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_40 ),
	.cout(Xd_0__inst_mult_29_41 ),
	.shareout(Xd_0__inst_mult_29_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_22 (
// Equation(s):
// Xd_0__inst_mult_31_67  = SUM(( GND ) + ( Xd_0__inst_mult_31_89  ) + ( Xd_0__inst_mult_31_88  ))
// Xd_0__inst_mult_31_68  = CARRY(( GND ) + ( Xd_0__inst_mult_31_89  ) + ( Xd_0__inst_mult_31_88  ))
// Xd_0__inst_mult_31_69  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_88 ),
	.sharein(Xd_0__inst_mult_31_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_67 ),
	.cout(Xd_0__inst_mult_31_68 ),
	.shareout(Xd_0__inst_mult_31_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11 (
// Equation(s):
// Xd_0__inst_mult_11_40  = SUM(( GND ) + ( Xd_0__inst_mult_11_77  ) + ( Xd_0__inst_mult_11_76  ))
// Xd_0__inst_mult_11_41  = CARRY(( GND ) + ( Xd_0__inst_mult_11_77  ) + ( Xd_0__inst_mult_11_76  ))
// Xd_0__inst_mult_11_42  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_76 ),
	.sharein(Xd_0__inst_mult_11_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_40 ),
	.cout(Xd_0__inst_mult_11_41 ),
	.shareout(Xd_0__inst_mult_11_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25 (
// Equation(s):
// Xd_0__inst_mult_25_40  = SUM(( GND ) + ( Xd_0__inst_mult_25_77  ) + ( Xd_0__inst_mult_25_76  ))
// Xd_0__inst_mult_25_41  = CARRY(( GND ) + ( Xd_0__inst_mult_25_77  ) + ( Xd_0__inst_mult_25_76  ))
// Xd_0__inst_mult_25_42  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_76 ),
	.sharein(Xd_0__inst_mult_25_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_40 ),
	.cout(Xd_0__inst_mult_25_41 ),
	.shareout(Xd_0__inst_mult_25_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27 (
// Equation(s):
// Xd_0__inst_mult_27_40  = SUM(( GND ) + ( Xd_0__inst_mult_27_77  ) + ( Xd_0__inst_mult_27_76  ))
// Xd_0__inst_mult_27_41  = CARRY(( GND ) + ( Xd_0__inst_mult_27_77  ) + ( Xd_0__inst_mult_27_76  ))
// Xd_0__inst_mult_27_42  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_76 ),
	.sharein(Xd_0__inst_mult_27_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_40 ),
	.cout(Xd_0__inst_mult_27_41 ),
	.shareout(Xd_0__inst_mult_27_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_25 (
// Equation(s):
// Xd_0__inst_mult_30_79  = SUM(( (din_a[180] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_30_80  = CARRY(( (din_a[180] & din_b[180]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_30_81  = SHARE((din_b[180] & din_a[181]))

	.dataa(!din_a[180]),
	.datab(!din_b[180]),
	.datac(!din_a[181]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_30_79 ),
	.cout(Xd_0__inst_mult_30_80 ),
	.shareout(Xd_0__inst_mult_30_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_23 (
// Equation(s):
// Xd_0__inst_mult_31_71  = SUM(( (din_a[186] & din_b[186]) ) + ( Xd_0__inst_mult_30_97  ) + ( Xd_0__inst_mult_30_96  ))
// Xd_0__inst_mult_31_72  = CARRY(( (din_a[186] & din_b[186]) ) + ( Xd_0__inst_mult_30_97  ) + ( Xd_0__inst_mult_30_96  ))
// Xd_0__inst_mult_31_73  = SHARE((din_b[186] & din_a[187]))

	.dataa(!din_a[186]),
	.datab(!din_b[186]),
	.datac(!din_a[187]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_96 ),
	.sharein(Xd_0__inst_mult_30_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_71 ),
	.cout(Xd_0__inst_mult_31_72 ),
	.shareout(Xd_0__inst_mult_31_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_13 (
// Equation(s):
// Xd_0__inst_i17_13_sumout  = SUM(( !din_a[185] $ (!din_b[185]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_14  = CARRY(( !din_a[185] $ (!din_b[185]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_15  = SHARE(GND)

	.dataa(!din_a[185]),
	.datab(!din_b[185]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_13_sumout ),
	.cout(Xd_0__inst_i17_14 ),
	.shareout(Xd_0__inst_i17_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_17 (
// Equation(s):
// Xd_0__inst_i17_17_sumout  = SUM(( !din_a[191] $ (!din_b[191]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_18  = CARRY(( !din_a[191] $ (!din_b[191]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_19  = SHARE(GND)

	.dataa(!din_a[191]),
	.datab(!din_b[191]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_17_sumout ),
	.cout(Xd_0__inst_i17_18 ),
	.shareout(Xd_0__inst_i17_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_30_26 (
// Equation(s):
// Xd_0__inst_mult_30_83  = SUM(( (din_a[180] & din_b[181]) ) + ( Xd_0__inst_mult_30_81  ) + ( Xd_0__inst_mult_30_80  ))
// Xd_0__inst_mult_30_84  = CARRY(( (din_a[180] & din_b[181]) ) + ( Xd_0__inst_mult_30_81  ) + ( Xd_0__inst_mult_30_80  ))
// Xd_0__inst_mult_30_85  = SHARE((din_b[180] & din_a[182]))

	.dataa(!din_a[180]),
	.datab(!din_b[180]),
	.datac(!din_b[181]),
	.datad(!din_a[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_80 ),
	.sharein(Xd_0__inst_mult_30_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_83 ),
	.cout(Xd_0__inst_mult_30_84 ),
	.shareout(Xd_0__inst_mult_30_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_31_24 (
// Equation(s):
// Xd_0__inst_mult_31_75  = SUM(( (din_a[186] & din_b[187]) ) + ( Xd_0__inst_mult_31_73  ) + ( Xd_0__inst_mult_31_72  ))
// Xd_0__inst_mult_31_76  = CARRY(( (din_a[186] & din_b[187]) ) + ( Xd_0__inst_mult_31_73  ) + ( Xd_0__inst_mult_31_72  ))
// Xd_0__inst_mult_31_77  = SHARE((din_b[186] & din_a[188]))

	.dataa(!din_a[186]),
	.datab(!din_b[186]),
	.datac(!din_b[187]),
	.datad(!din_a[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_72 ),
	.sharein(Xd_0__inst_mult_31_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_75 ),
	.cout(Xd_0__inst_mult_31_76 ),
	.shareout(Xd_0__inst_mult_31_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_27 (
// Equation(s):
// Xd_0__inst_mult_30_87  = SUM(( (!din_a[181] & (((din_a[180] & din_b[182])))) # (din_a[181] & (!din_b[181] $ (((!din_a[180]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_30_85  ) + ( Xd_0__inst_mult_30_84  ))
// Xd_0__inst_mult_30_88  = CARRY(( (!din_a[181] & (((din_a[180] & din_b[182])))) # (din_a[181] & (!din_b[181] $ (((!din_a[180]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_30_85  ) + ( Xd_0__inst_mult_30_84  ))
// Xd_0__inst_mult_30_89  = SHARE((din_a[181] & (din_b[181] & (din_a[180] & din_b[182]))))

	.dataa(!din_a[181]),
	.datab(!din_b[181]),
	.datac(!din_a[180]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_84 ),
	.sharein(Xd_0__inst_mult_30_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_87 ),
	.cout(Xd_0__inst_mult_30_88 ),
	.shareout(Xd_0__inst_mult_30_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_25 (
// Equation(s):
// Xd_0__inst_mult_31_79  = SUM(( (!din_a[187] & (((din_a[186] & din_b[188])))) # (din_a[187] & (!din_b[187] $ (((!din_a[186]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_31_77  ) + ( Xd_0__inst_mult_31_76  ))
// Xd_0__inst_mult_31_80  = CARRY(( (!din_a[187] & (((din_a[186] & din_b[188])))) # (din_a[187] & (!din_b[187] $ (((!din_a[186]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_31_77  ) + ( Xd_0__inst_mult_31_76  ))
// Xd_0__inst_mult_31_81  = SHARE((din_a[187] & (din_b[187] & (din_a[186] & din_b[188]))))

	.dataa(!din_a[187]),
	.datab(!din_b[187]),
	.datac(!din_a[186]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_76 ),
	.sharein(Xd_0__inst_mult_31_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_79 ),
	.cout(Xd_0__inst_mult_31_80 ),
	.shareout(Xd_0__inst_mult_31_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_16_34 (
// Equation(s):
// Xd_0__inst_mult_16_35  = SUM(( Xd_0__inst_mult_16_5_q  ) + ( Xd_0__inst_mult_16_72  ) + ( Xd_0__inst_mult_16_71  ))
// Xd_0__inst_mult_16_36  = CARRY(( Xd_0__inst_mult_16_5_q  ) + ( Xd_0__inst_mult_16_72  ) + ( Xd_0__inst_mult_16_71  ))
// Xd_0__inst_mult_16_37  = SHARE((Xd_0__inst_mult_16_4_q  & Xd_0__inst_mult_16_2_q ))

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_2_q ),
	.datac(!Xd_0__inst_mult_16_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_71 ),
	.sharein(Xd_0__inst_mult_16_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_35 ),
	.cout(Xd_0__inst_mult_16_36 ),
	.shareout(Xd_0__inst_mult_16_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_17_35 (
// Equation(s):
// Xd_0__inst_mult_17_36  = SUM(( Xd_0__inst_mult_17_5_q  ) + ( Xd_0__inst_mult_17_81  ) + ( Xd_0__inst_mult_17_80  ))
// Xd_0__inst_mult_17_37  = CARRY(( Xd_0__inst_mult_17_5_q  ) + ( Xd_0__inst_mult_17_81  ) + ( Xd_0__inst_mult_17_80  ))
// Xd_0__inst_mult_17_38  = SHARE((Xd_0__inst_mult_17_4_q  & Xd_0__inst_mult_17_2_q ))

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_2_q ),
	.datac(!Xd_0__inst_mult_17_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_80 ),
	.sharein(Xd_0__inst_mult_17_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_36 ),
	.cout(Xd_0__inst_mult_17_37 ),
	.shareout(Xd_0__inst_mult_17_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_14_34 (
// Equation(s):
// Xd_0__inst_mult_14_35  = SUM(( Xd_0__inst_mult_14_5_q  ) + ( Xd_0__inst_mult_14_72  ) + ( Xd_0__inst_mult_14_71  ))
// Xd_0__inst_mult_14_36  = CARRY(( Xd_0__inst_mult_14_5_q  ) + ( Xd_0__inst_mult_14_72  ) + ( Xd_0__inst_mult_14_71  ))
// Xd_0__inst_mult_14_37  = SHARE((Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_2_q ))

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_2_q ),
	.datac(!Xd_0__inst_mult_14_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_71 ),
	.sharein(Xd_0__inst_mult_14_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_35 ),
	.cout(Xd_0__inst_mult_14_36 ),
	.shareout(Xd_0__inst_mult_14_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_15_35 (
// Equation(s):
// Xd_0__inst_mult_15_36  = SUM(( Xd_0__inst_mult_15_5_q  ) + ( Xd_0__inst_mult_15_81  ) + ( Xd_0__inst_mult_15_80  ))
// Xd_0__inst_mult_15_37  = CARRY(( Xd_0__inst_mult_15_5_q  ) + ( Xd_0__inst_mult_15_81  ) + ( Xd_0__inst_mult_15_80  ))
// Xd_0__inst_mult_15_38  = SHARE((Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_2_q ))

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_2_q ),
	.datac(!Xd_0__inst_mult_15_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_80 ),
	.sharein(Xd_0__inst_mult_15_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_36 ),
	.cout(Xd_0__inst_mult_15_37 ),
	.shareout(Xd_0__inst_mult_15_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_12_34 (
// Equation(s):
// Xd_0__inst_mult_12_35  = SUM(( Xd_0__inst_mult_12_5_q  ) + ( Xd_0__inst_mult_12_72  ) + ( Xd_0__inst_mult_12_71  ))
// Xd_0__inst_mult_12_36  = CARRY(( Xd_0__inst_mult_12_5_q  ) + ( Xd_0__inst_mult_12_72  ) + ( Xd_0__inst_mult_12_71  ))
// Xd_0__inst_mult_12_37  = SHARE((Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_2_q ))

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_2_q ),
	.datac(!Xd_0__inst_mult_12_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_71 ),
	.sharein(Xd_0__inst_mult_12_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_35 ),
	.cout(Xd_0__inst_mult_12_36 ),
	.shareout(Xd_0__inst_mult_12_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_13_35 (
// Equation(s):
// Xd_0__inst_mult_13_36  = SUM(( Xd_0__inst_mult_13_5_q  ) + ( Xd_0__inst_mult_13_81  ) + ( Xd_0__inst_mult_13_80  ))
// Xd_0__inst_mult_13_37  = CARRY(( Xd_0__inst_mult_13_5_q  ) + ( Xd_0__inst_mult_13_81  ) + ( Xd_0__inst_mult_13_80  ))
// Xd_0__inst_mult_13_38  = SHARE((Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_2_q ))

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_2_q ),
	.datac(!Xd_0__inst_mult_13_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_80 ),
	.sharein(Xd_0__inst_mult_13_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_36 ),
	.cout(Xd_0__inst_mult_13_37 ),
	.shareout(Xd_0__inst_mult_13_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_10_34 (
// Equation(s):
// Xd_0__inst_mult_10_35  = SUM(( Xd_0__inst_mult_10_5_q  ) + ( Xd_0__inst_mult_10_72  ) + ( Xd_0__inst_mult_10_71  ))
// Xd_0__inst_mult_10_36  = CARRY(( Xd_0__inst_mult_10_5_q  ) + ( Xd_0__inst_mult_10_72  ) + ( Xd_0__inst_mult_10_71  ))
// Xd_0__inst_mult_10_37  = SHARE((Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_2_q ))

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_2_q ),
	.datac(!Xd_0__inst_mult_10_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_71 ),
	.sharein(Xd_0__inst_mult_10_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_35 ),
	.cout(Xd_0__inst_mult_10_36 ),
	.shareout(Xd_0__inst_mult_10_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_11_16 (
// Equation(s):
// Xd_0__inst_mult_11_43  = SUM(( Xd_0__inst_mult_11_5_q  ) + ( Xd_0__inst_mult_11_89  ) + ( Xd_0__inst_mult_11_88  ))
// Xd_0__inst_mult_11_44  = CARRY(( Xd_0__inst_mult_11_5_q  ) + ( Xd_0__inst_mult_11_89  ) + ( Xd_0__inst_mult_11_88  ))
// Xd_0__inst_mult_11_45  = SHARE((Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_2_q ))

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_2_q ),
	.datac(!Xd_0__inst_mult_11_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_88 ),
	.sharein(Xd_0__inst_mult_11_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_43 ),
	.cout(Xd_0__inst_mult_11_44 ),
	.shareout(Xd_0__inst_mult_11_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_8_34 (
// Equation(s):
// Xd_0__inst_mult_8_35  = SUM(( Xd_0__inst_mult_8_5_q  ) + ( Xd_0__inst_mult_8_72  ) + ( Xd_0__inst_mult_8_71  ))
// Xd_0__inst_mult_8_36  = CARRY(( Xd_0__inst_mult_8_5_q  ) + ( Xd_0__inst_mult_8_72  ) + ( Xd_0__inst_mult_8_71  ))
// Xd_0__inst_mult_8_37  = SHARE((Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_2_q ))

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_2_q ),
	.datac(!Xd_0__inst_mult_8_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_71 ),
	.sharein(Xd_0__inst_mult_8_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_35 ),
	.cout(Xd_0__inst_mult_8_36 ),
	.shareout(Xd_0__inst_mult_8_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_9_35 (
// Equation(s):
// Xd_0__inst_mult_9_36  = SUM(( Xd_0__inst_mult_9_5_q  ) + ( Xd_0__inst_mult_9_81  ) + ( Xd_0__inst_mult_9_80  ))
// Xd_0__inst_mult_9_37  = CARRY(( Xd_0__inst_mult_9_5_q  ) + ( Xd_0__inst_mult_9_81  ) + ( Xd_0__inst_mult_9_80  ))
// Xd_0__inst_mult_9_38  = SHARE((Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_2_q ))

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_2_q ),
	.datac(!Xd_0__inst_mult_9_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_80 ),
	.sharein(Xd_0__inst_mult_9_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_36 ),
	.cout(Xd_0__inst_mult_9_37 ),
	.shareout(Xd_0__inst_mult_9_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_6_33 (
// Equation(s):
// Xd_0__inst_mult_6_34  = SUM(( Xd_0__inst_mult_6_5_q  ) + ( Xd_0__inst_mult_6_71  ) + ( Xd_0__inst_mult_6_70  ))
// Xd_0__inst_mult_6_35  = CARRY(( Xd_0__inst_mult_6_5_q  ) + ( Xd_0__inst_mult_6_71  ) + ( Xd_0__inst_mult_6_70  ))
// Xd_0__inst_mult_6_36  = SHARE((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_2_q ))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_2_q ),
	.datac(!Xd_0__inst_mult_6_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_70 ),
	.sharein(Xd_0__inst_mult_6_71 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_34 ),
	.cout(Xd_0__inst_mult_6_35 ),
	.shareout(Xd_0__inst_mult_6_36 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_7_34 (
// Equation(s):
// Xd_0__inst_mult_7_35  = SUM(( Xd_0__inst_mult_7_5_q  ) + ( Xd_0__inst_mult_7_80  ) + ( Xd_0__inst_mult_7_79  ))
// Xd_0__inst_mult_7_36  = CARRY(( Xd_0__inst_mult_7_5_q  ) + ( Xd_0__inst_mult_7_80  ) + ( Xd_0__inst_mult_7_79  ))
// Xd_0__inst_mult_7_37  = SHARE((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_2_q ))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_2_q ),
	.datac(!Xd_0__inst_mult_7_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_79 ),
	.sharein(Xd_0__inst_mult_7_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_35 ),
	.cout(Xd_0__inst_mult_7_36 ),
	.shareout(Xd_0__inst_mult_7_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_4_33 (
// Equation(s):
// Xd_0__inst_mult_4_34  = SUM(( Xd_0__inst_mult_4_5_q  ) + ( Xd_0__inst_mult_4_71  ) + ( Xd_0__inst_mult_4_70  ))
// Xd_0__inst_mult_4_35  = CARRY(( Xd_0__inst_mult_4_5_q  ) + ( Xd_0__inst_mult_4_71  ) + ( Xd_0__inst_mult_4_70  ))
// Xd_0__inst_mult_4_36  = SHARE((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_2_q ))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_2_q ),
	.datac(!Xd_0__inst_mult_4_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_70 ),
	.sharein(Xd_0__inst_mult_4_71 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_34 ),
	.cout(Xd_0__inst_mult_4_35 ),
	.shareout(Xd_0__inst_mult_4_36 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_5_34 (
// Equation(s):
// Xd_0__inst_mult_5_35  = SUM(( Xd_0__inst_mult_5_5_q  ) + ( Xd_0__inst_mult_5_80  ) + ( Xd_0__inst_mult_5_79  ))
// Xd_0__inst_mult_5_36  = CARRY(( Xd_0__inst_mult_5_5_q  ) + ( Xd_0__inst_mult_5_80  ) + ( Xd_0__inst_mult_5_79  ))
// Xd_0__inst_mult_5_37  = SHARE((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_2_q ))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_2_q ),
	.datac(!Xd_0__inst_mult_5_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_79 ),
	.sharein(Xd_0__inst_mult_5_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_35 ),
	.cout(Xd_0__inst_mult_5_36 ),
	.shareout(Xd_0__inst_mult_5_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_2 (
// Equation(s):
// Xd_0__inst_mult_2_39  = SUM(( Xd_0__inst_mult_2_5_q  ) + ( Xd_0__inst_mult_2_80  ) + ( Xd_0__inst_mult_2_79  ))
// Xd_0__inst_mult_2_40  = CARRY(( Xd_0__inst_mult_2_5_q  ) + ( Xd_0__inst_mult_2_80  ) + ( Xd_0__inst_mult_2_79  ))
// Xd_0__inst_mult_2_41  = SHARE((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_2_q ))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_2_q ),
	.datac(!Xd_0__inst_mult_2_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_79 ),
	.sharein(Xd_0__inst_mult_2_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_39 ),
	.cout(Xd_0__inst_mult_2_40 ),
	.shareout(Xd_0__inst_mult_2_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_3 (
// Equation(s):
// Xd_0__inst_mult_3_39  = SUM(( Xd_0__inst_mult_3_5_q  ) + ( Xd_0__inst_mult_3_80  ) + ( Xd_0__inst_mult_3_79  ))
// Xd_0__inst_mult_3_40  = CARRY(( Xd_0__inst_mult_3_5_q  ) + ( Xd_0__inst_mult_3_80  ) + ( Xd_0__inst_mult_3_79  ))
// Xd_0__inst_mult_3_41  = SHARE((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_2_q ))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_2_q ),
	.datac(!Xd_0__inst_mult_3_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_79 ),
	.sharein(Xd_0__inst_mult_3_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_39 ),
	.cout(Xd_0__inst_mult_3_40 ),
	.shareout(Xd_0__inst_mult_3_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_0 (
// Equation(s):
// Xd_0__inst_mult_0_39  = SUM(( Xd_0__inst_mult_0_5_q  ) + ( Xd_0__inst_mult_0_80  ) + ( Xd_0__inst_mult_0_79  ))
// Xd_0__inst_mult_0_40  = CARRY(( Xd_0__inst_mult_0_5_q  ) + ( Xd_0__inst_mult_0_80  ) + ( Xd_0__inst_mult_0_79  ))
// Xd_0__inst_mult_0_41  = SHARE((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_2_q ))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_2_q ),
	.datac(!Xd_0__inst_mult_0_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_79 ),
	.sharein(Xd_0__inst_mult_0_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_39 ),
	.cout(Xd_0__inst_mult_0_40 ),
	.shareout(Xd_0__inst_mult_0_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_1 (
// Equation(s):
// Xd_0__inst_mult_1_39  = SUM(( Xd_0__inst_mult_1_5_q  ) + ( Xd_0__inst_mult_1_80  ) + ( Xd_0__inst_mult_1_79  ))
// Xd_0__inst_mult_1_40  = CARRY(( Xd_0__inst_mult_1_5_q  ) + ( Xd_0__inst_mult_1_80  ) + ( Xd_0__inst_mult_1_79  ))
// Xd_0__inst_mult_1_41  = SHARE((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_2_q ))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_2_q ),
	.datac(!Xd_0__inst_mult_1_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_79 ),
	.sharein(Xd_0__inst_mult_1_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_39 ),
	.cout(Xd_0__inst_mult_1_40 ),
	.shareout(Xd_0__inst_mult_1_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_28_18 (
// Equation(s):
// Xd_0__inst_mult_28_51  = SUM(( Xd_0__inst_mult_28_5_q  ) + ( Xd_0__inst_mult_28_93  ) + ( Xd_0__inst_mult_28_92  ))
// Xd_0__inst_mult_28_52  = CARRY(( Xd_0__inst_mult_28_5_q  ) + ( Xd_0__inst_mult_28_93  ) + ( Xd_0__inst_mult_28_92  ))
// Xd_0__inst_mult_28_53  = SHARE((Xd_0__inst_mult_28_4_q  & Xd_0__inst_mult_28_2_q ))

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_2_q ),
	.datac(!Xd_0__inst_mult_28_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_92 ),
	.sharein(Xd_0__inst_mult_28_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_51 ),
	.cout(Xd_0__inst_mult_28_52 ),
	.shareout(Xd_0__inst_mult_28_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_29_16 (
// Equation(s):
// Xd_0__inst_mult_29_43  = SUM(( Xd_0__inst_mult_29_5_q  ) + ( Xd_0__inst_mult_29_89  ) + ( Xd_0__inst_mult_29_88  ))
// Xd_0__inst_mult_29_44  = CARRY(( Xd_0__inst_mult_29_5_q  ) + ( Xd_0__inst_mult_29_89  ) + ( Xd_0__inst_mult_29_88  ))
// Xd_0__inst_mult_29_45  = SHARE((Xd_0__inst_mult_29_4_q  & Xd_0__inst_mult_29_2_q ))

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_2_q ),
	.datac(!Xd_0__inst_mult_29_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_88 ),
	.sharein(Xd_0__inst_mult_29_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_43 ),
	.cout(Xd_0__inst_mult_29_44 ),
	.shareout(Xd_0__inst_mult_29_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_26_18 (
// Equation(s):
// Xd_0__inst_mult_26_51  = SUM(( Xd_0__inst_mult_26_5_q  ) + ( Xd_0__inst_mult_26_93  ) + ( Xd_0__inst_mult_26_92  ))
// Xd_0__inst_mult_26_52  = CARRY(( Xd_0__inst_mult_26_5_q  ) + ( Xd_0__inst_mult_26_93  ) + ( Xd_0__inst_mult_26_92  ))
// Xd_0__inst_mult_26_53  = SHARE((Xd_0__inst_mult_26_4_q  & Xd_0__inst_mult_26_2_q ))

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_2_q ),
	.datac(!Xd_0__inst_mult_26_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_92 ),
	.sharein(Xd_0__inst_mult_26_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_51 ),
	.cout(Xd_0__inst_mult_26_52 ),
	.shareout(Xd_0__inst_mult_26_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_27_16 (
// Equation(s):
// Xd_0__inst_mult_27_43  = SUM(( Xd_0__inst_mult_27_5_q  ) + ( Xd_0__inst_mult_27_89  ) + ( Xd_0__inst_mult_27_88  ))
// Xd_0__inst_mult_27_44  = CARRY(( Xd_0__inst_mult_27_5_q  ) + ( Xd_0__inst_mult_27_89  ) + ( Xd_0__inst_mult_27_88  ))
// Xd_0__inst_mult_27_45  = SHARE((Xd_0__inst_mult_27_4_q  & Xd_0__inst_mult_27_2_q ))

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_2_q ),
	.datac(!Xd_0__inst_mult_27_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_88 ),
	.sharein(Xd_0__inst_mult_27_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_43 ),
	.cout(Xd_0__inst_mult_27_44 ),
	.shareout(Xd_0__inst_mult_27_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_24_18 (
// Equation(s):
// Xd_0__inst_mult_24_51  = SUM(( Xd_0__inst_mult_24_5_q  ) + ( Xd_0__inst_mult_24_93  ) + ( Xd_0__inst_mult_24_92  ))
// Xd_0__inst_mult_24_52  = CARRY(( Xd_0__inst_mult_24_5_q  ) + ( Xd_0__inst_mult_24_93  ) + ( Xd_0__inst_mult_24_92  ))
// Xd_0__inst_mult_24_53  = SHARE((Xd_0__inst_mult_24_4_q  & Xd_0__inst_mult_24_2_q ))

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_2_q ),
	.datac(!Xd_0__inst_mult_24_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_92 ),
	.sharein(Xd_0__inst_mult_24_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_51 ),
	.cout(Xd_0__inst_mult_24_52 ),
	.shareout(Xd_0__inst_mult_24_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_25_16 (
// Equation(s):
// Xd_0__inst_mult_25_43  = SUM(( Xd_0__inst_mult_25_5_q  ) + ( Xd_0__inst_mult_25_89  ) + ( Xd_0__inst_mult_25_88  ))
// Xd_0__inst_mult_25_44  = CARRY(( Xd_0__inst_mult_25_5_q  ) + ( Xd_0__inst_mult_25_89  ) + ( Xd_0__inst_mult_25_88  ))
// Xd_0__inst_mult_25_45  = SHARE((Xd_0__inst_mult_25_4_q  & Xd_0__inst_mult_25_2_q ))

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_2_q ),
	.datac(!Xd_0__inst_mult_25_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_88 ),
	.sharein(Xd_0__inst_mult_25_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_43 ),
	.cout(Xd_0__inst_mult_25_44 ),
	.shareout(Xd_0__inst_mult_25_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_22_18 (
// Equation(s):
// Xd_0__inst_mult_22_51  = SUM(( Xd_0__inst_mult_22_5_q  ) + ( Xd_0__inst_mult_22_93  ) + ( Xd_0__inst_mult_22_92  ))
// Xd_0__inst_mult_22_52  = CARRY(( Xd_0__inst_mult_22_5_q  ) + ( Xd_0__inst_mult_22_93  ) + ( Xd_0__inst_mult_22_92  ))
// Xd_0__inst_mult_22_53  = SHARE((Xd_0__inst_mult_22_4_q  & Xd_0__inst_mult_22_2_q ))

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_2_q ),
	.datac(!Xd_0__inst_mult_22_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_92 ),
	.sharein(Xd_0__inst_mult_22_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_51 ),
	.cout(Xd_0__inst_mult_22_52 ),
	.shareout(Xd_0__inst_mult_22_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_23_18 (
// Equation(s):
// Xd_0__inst_mult_23_51  = SUM(( Xd_0__inst_mult_23_5_q  ) + ( Xd_0__inst_mult_23_93  ) + ( Xd_0__inst_mult_23_92  ))
// Xd_0__inst_mult_23_52  = CARRY(( Xd_0__inst_mult_23_5_q  ) + ( Xd_0__inst_mult_23_93  ) + ( Xd_0__inst_mult_23_92  ))
// Xd_0__inst_mult_23_53  = SHARE((Xd_0__inst_mult_23_4_q  & Xd_0__inst_mult_23_2_q ))

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_2_q ),
	.datac(!Xd_0__inst_mult_23_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_92 ),
	.sharein(Xd_0__inst_mult_23_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_51 ),
	.cout(Xd_0__inst_mult_23_52 ),
	.shareout(Xd_0__inst_mult_23_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_20_18 (
// Equation(s):
// Xd_0__inst_mult_20_51  = SUM(( Xd_0__inst_mult_20_5_q  ) + ( Xd_0__inst_mult_20_93  ) + ( Xd_0__inst_mult_20_92  ))
// Xd_0__inst_mult_20_52  = CARRY(( Xd_0__inst_mult_20_5_q  ) + ( Xd_0__inst_mult_20_93  ) + ( Xd_0__inst_mult_20_92  ))
// Xd_0__inst_mult_20_53  = SHARE((Xd_0__inst_mult_20_4_q  & Xd_0__inst_mult_20_2_q ))

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_2_q ),
	.datac(!Xd_0__inst_mult_20_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_92 ),
	.sharein(Xd_0__inst_mult_20_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_51 ),
	.cout(Xd_0__inst_mult_20_52 ),
	.shareout(Xd_0__inst_mult_20_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_21_35 (
// Equation(s):
// Xd_0__inst_mult_21_36  = SUM(( Xd_0__inst_mult_21_5_q  ) + ( Xd_0__inst_mult_21_81  ) + ( Xd_0__inst_mult_21_80  ))
// Xd_0__inst_mult_21_37  = CARRY(( Xd_0__inst_mult_21_5_q  ) + ( Xd_0__inst_mult_21_81  ) + ( Xd_0__inst_mult_21_80  ))
// Xd_0__inst_mult_21_38  = SHARE((Xd_0__inst_mult_21_4_q  & Xd_0__inst_mult_21_2_q ))

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_2_q ),
	.datac(!Xd_0__inst_mult_21_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_80 ),
	.sharein(Xd_0__inst_mult_21_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_36 ),
	.cout(Xd_0__inst_mult_21_37 ),
	.shareout(Xd_0__inst_mult_21_38 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_18_34 (
// Equation(s):
// Xd_0__inst_mult_18_35  = SUM(( Xd_0__inst_mult_18_5_q  ) + ( Xd_0__inst_mult_18_72  ) + ( Xd_0__inst_mult_18_71  ))
// Xd_0__inst_mult_18_36  = CARRY(( Xd_0__inst_mult_18_5_q  ) + ( Xd_0__inst_mult_18_72  ) + ( Xd_0__inst_mult_18_71  ))
// Xd_0__inst_mult_18_37  = SHARE((Xd_0__inst_mult_18_4_q  & Xd_0__inst_mult_18_2_q ))

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_2_q ),
	.datac(!Xd_0__inst_mult_18_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_71 ),
	.sharein(Xd_0__inst_mult_18_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_35 ),
	.cout(Xd_0__inst_mult_18_36 ),
	.shareout(Xd_0__inst_mult_18_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000F0F),
	.shared_arith("on")
) Xd_0__inst_mult_19_17 (
// Equation(s):
// Xd_0__inst_mult_19_47  = SUM(( Xd_0__inst_mult_19_5_q  ) + ( Xd_0__inst_mult_19_93  ) + ( Xd_0__inst_mult_19_92  ))
// Xd_0__inst_mult_19_48  = CARRY(( Xd_0__inst_mult_19_5_q  ) + ( Xd_0__inst_mult_19_93  ) + ( Xd_0__inst_mult_19_92  ))
// Xd_0__inst_mult_19_49  = SHARE((Xd_0__inst_mult_19_4_q  & Xd_0__inst_mult_19_2_q ))

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_2_q ),
	.datac(!Xd_0__inst_mult_19_5_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_92 ),
	.sharein(Xd_0__inst_mult_19_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_47 ),
	.cout(Xd_0__inst_mult_19_48 ),
	.shareout(Xd_0__inst_mult_19_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_28 (
// Equation(s):
// Xd_0__inst_mult_30_92  = CARRY(( (Xd_0__inst_mult_30_0_q  & Xd_0__inst_mult_30_1_q ) ) + ( Xd_0__inst_mult_30_45  ) + ( Xd_0__inst_mult_30_44  ))
// Xd_0__inst_mult_30_93  = SHARE((Xd_0__inst_mult_30_2_q  & Xd_0__inst_mult_30_3_q ))

	.dataa(!Xd_0__inst_mult_30_0_q ),
	.datab(!Xd_0__inst_mult_30_1_q ),
	.datac(!Xd_0__inst_mult_30_2_q ),
	.datad(!Xd_0__inst_mult_30_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_44 ),
	.sharein(Xd_0__inst_mult_30_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_30_92 ),
	.shareout(Xd_0__inst_mult_30_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_26 (
// Equation(s):
// Xd_0__inst_mult_31_84  = CARRY(( (Xd_0__inst_mult_31_0_q  & Xd_0__inst_mult_31_1_q ) ) + ( Xd_0__inst_mult_31_38  ) + ( Xd_0__inst_mult_31_37  ))
// Xd_0__inst_mult_31_85  = SHARE((Xd_0__inst_mult_31_2_q  & Xd_0__inst_mult_31_3_q ))

	.dataa(!Xd_0__inst_mult_31_0_q ),
	.datab(!Xd_0__inst_mult_31_1_q ),
	.datac(!Xd_0__inst_mult_31_2_q ),
	.datad(!Xd_0__inst_mult_31_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_37 ),
	.sharein(Xd_0__inst_mult_31_38 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_84 ),
	.shareout(Xd_0__inst_mult_31_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_16 (
// Equation(s):
// Xd_0__inst_mult_16_39  = SUM(( !Xd_0__inst_mult_16_6_q  $ (!Xd_0__inst_mult_16_7_q ) ) + ( Xd_0__inst_mult_16_37  ) + ( Xd_0__inst_mult_16_36  ))
// Xd_0__inst_mult_16_40  = CARRY(( !Xd_0__inst_mult_16_6_q  $ (!Xd_0__inst_mult_16_7_q ) ) + ( Xd_0__inst_mult_16_37  ) + ( Xd_0__inst_mult_16_36  ))
// Xd_0__inst_mult_16_41  = SHARE((Xd_0__inst_mult_16_6_q  & Xd_0__inst_mult_16_7_q ))

	.dataa(!Xd_0__inst_mult_16_6_q ),
	.datab(!Xd_0__inst_mult_16_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_36 ),
	.sharein(Xd_0__inst_mult_16_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_39 ),
	.cout(Xd_0__inst_mult_16_40 ),
	.shareout(Xd_0__inst_mult_16_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_17 (
// Equation(s):
// Xd_0__inst_mult_17_40  = SUM(( !Xd_0__inst_mult_17_6_q  $ (!Xd_0__inst_mult_17_7_q ) ) + ( Xd_0__inst_mult_17_38  ) + ( Xd_0__inst_mult_17_37  ))
// Xd_0__inst_mult_17_41  = CARRY(( !Xd_0__inst_mult_17_6_q  $ (!Xd_0__inst_mult_17_7_q ) ) + ( Xd_0__inst_mult_17_38  ) + ( Xd_0__inst_mult_17_37  ))
// Xd_0__inst_mult_17_42  = SHARE((Xd_0__inst_mult_17_6_q  & Xd_0__inst_mult_17_7_q ))

	.dataa(!Xd_0__inst_mult_17_6_q ),
	.datab(!Xd_0__inst_mult_17_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_37 ),
	.sharein(Xd_0__inst_mult_17_38 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_40 ),
	.cout(Xd_0__inst_mult_17_41 ),
	.shareout(Xd_0__inst_mult_17_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_14 (
// Equation(s):
// Xd_0__inst_mult_14_39  = SUM(( !Xd_0__inst_mult_14_6_q  $ (!Xd_0__inst_mult_14_7_q ) ) + ( Xd_0__inst_mult_14_37  ) + ( Xd_0__inst_mult_14_36  ))
// Xd_0__inst_mult_14_40  = CARRY(( !Xd_0__inst_mult_14_6_q  $ (!Xd_0__inst_mult_14_7_q ) ) + ( Xd_0__inst_mult_14_37  ) + ( Xd_0__inst_mult_14_36  ))
// Xd_0__inst_mult_14_41  = SHARE((Xd_0__inst_mult_14_6_q  & Xd_0__inst_mult_14_7_q ))

	.dataa(!Xd_0__inst_mult_14_6_q ),
	.datab(!Xd_0__inst_mult_14_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_36 ),
	.sharein(Xd_0__inst_mult_14_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_39 ),
	.cout(Xd_0__inst_mult_14_40 ),
	.shareout(Xd_0__inst_mult_14_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_15 (
// Equation(s):
// Xd_0__inst_mult_15_40  = SUM(( !Xd_0__inst_mult_15_6_q  $ (!Xd_0__inst_mult_15_7_q ) ) + ( Xd_0__inst_mult_15_38  ) + ( Xd_0__inst_mult_15_37  ))
// Xd_0__inst_mult_15_41  = CARRY(( !Xd_0__inst_mult_15_6_q  $ (!Xd_0__inst_mult_15_7_q ) ) + ( Xd_0__inst_mult_15_38  ) + ( Xd_0__inst_mult_15_37  ))
// Xd_0__inst_mult_15_42  = SHARE((Xd_0__inst_mult_15_6_q  & Xd_0__inst_mult_15_7_q ))

	.dataa(!Xd_0__inst_mult_15_6_q ),
	.datab(!Xd_0__inst_mult_15_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_37 ),
	.sharein(Xd_0__inst_mult_15_38 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_40 ),
	.cout(Xd_0__inst_mult_15_41 ),
	.shareout(Xd_0__inst_mult_15_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_12 (
// Equation(s):
// Xd_0__inst_mult_12_39  = SUM(( !Xd_0__inst_mult_12_6_q  $ (!Xd_0__inst_mult_12_7_q ) ) + ( Xd_0__inst_mult_12_37  ) + ( Xd_0__inst_mult_12_36  ))
// Xd_0__inst_mult_12_40  = CARRY(( !Xd_0__inst_mult_12_6_q  $ (!Xd_0__inst_mult_12_7_q ) ) + ( Xd_0__inst_mult_12_37  ) + ( Xd_0__inst_mult_12_36  ))
// Xd_0__inst_mult_12_41  = SHARE((Xd_0__inst_mult_12_6_q  & Xd_0__inst_mult_12_7_q ))

	.dataa(!Xd_0__inst_mult_12_6_q ),
	.datab(!Xd_0__inst_mult_12_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_36 ),
	.sharein(Xd_0__inst_mult_12_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_39 ),
	.cout(Xd_0__inst_mult_12_40 ),
	.shareout(Xd_0__inst_mult_12_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_13 (
// Equation(s):
// Xd_0__inst_mult_13_40  = SUM(( !Xd_0__inst_mult_13_6_q  $ (!Xd_0__inst_mult_13_7_q ) ) + ( Xd_0__inst_mult_13_38  ) + ( Xd_0__inst_mult_13_37  ))
// Xd_0__inst_mult_13_41  = CARRY(( !Xd_0__inst_mult_13_6_q  $ (!Xd_0__inst_mult_13_7_q ) ) + ( Xd_0__inst_mult_13_38  ) + ( Xd_0__inst_mult_13_37  ))
// Xd_0__inst_mult_13_42  = SHARE((Xd_0__inst_mult_13_6_q  & Xd_0__inst_mult_13_7_q ))

	.dataa(!Xd_0__inst_mult_13_6_q ),
	.datab(!Xd_0__inst_mult_13_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_37 ),
	.sharein(Xd_0__inst_mult_13_38 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_40 ),
	.cout(Xd_0__inst_mult_13_41 ),
	.shareout(Xd_0__inst_mult_13_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_10 (
// Equation(s):
// Xd_0__inst_mult_10_39  = SUM(( !Xd_0__inst_mult_10_6_q  $ (!Xd_0__inst_mult_10_7_q ) ) + ( Xd_0__inst_mult_10_37  ) + ( Xd_0__inst_mult_10_36  ))
// Xd_0__inst_mult_10_40  = CARRY(( !Xd_0__inst_mult_10_6_q  $ (!Xd_0__inst_mult_10_7_q ) ) + ( Xd_0__inst_mult_10_37  ) + ( Xd_0__inst_mult_10_36  ))
// Xd_0__inst_mult_10_41  = SHARE((Xd_0__inst_mult_10_6_q  & Xd_0__inst_mult_10_7_q ))

	.dataa(!Xd_0__inst_mult_10_6_q ),
	.datab(!Xd_0__inst_mult_10_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_36 ),
	.sharein(Xd_0__inst_mult_10_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_39 ),
	.cout(Xd_0__inst_mult_10_40 ),
	.shareout(Xd_0__inst_mult_10_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_11_17 (
// Equation(s):
// Xd_0__inst_mult_11_47  = SUM(( !Xd_0__inst_mult_11_6_q  $ (!Xd_0__inst_mult_11_7_q ) ) + ( Xd_0__inst_mult_11_45  ) + ( Xd_0__inst_mult_11_44  ))
// Xd_0__inst_mult_11_48  = CARRY(( !Xd_0__inst_mult_11_6_q  $ (!Xd_0__inst_mult_11_7_q ) ) + ( Xd_0__inst_mult_11_45  ) + ( Xd_0__inst_mult_11_44  ))
// Xd_0__inst_mult_11_49  = SHARE((Xd_0__inst_mult_11_6_q  & Xd_0__inst_mult_11_7_q ))

	.dataa(!Xd_0__inst_mult_11_6_q ),
	.datab(!Xd_0__inst_mult_11_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_44 ),
	.sharein(Xd_0__inst_mult_11_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_47 ),
	.cout(Xd_0__inst_mult_11_48 ),
	.shareout(Xd_0__inst_mult_11_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_8 (
// Equation(s):
// Xd_0__inst_mult_8_39  = SUM(( !Xd_0__inst_mult_8_6_q  $ (!Xd_0__inst_mult_8_7_q ) ) + ( Xd_0__inst_mult_8_37  ) + ( Xd_0__inst_mult_8_36  ))
// Xd_0__inst_mult_8_40  = CARRY(( !Xd_0__inst_mult_8_6_q  $ (!Xd_0__inst_mult_8_7_q ) ) + ( Xd_0__inst_mult_8_37  ) + ( Xd_0__inst_mult_8_36  ))
// Xd_0__inst_mult_8_41  = SHARE((Xd_0__inst_mult_8_6_q  & Xd_0__inst_mult_8_7_q ))

	.dataa(!Xd_0__inst_mult_8_6_q ),
	.datab(!Xd_0__inst_mult_8_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_36 ),
	.sharein(Xd_0__inst_mult_8_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_39 ),
	.cout(Xd_0__inst_mult_8_40 ),
	.shareout(Xd_0__inst_mult_8_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_9 (
// Equation(s):
// Xd_0__inst_mult_9_40  = SUM(( !Xd_0__inst_mult_9_6_q  $ (!Xd_0__inst_mult_9_7_q ) ) + ( Xd_0__inst_mult_9_38  ) + ( Xd_0__inst_mult_9_37  ))
// Xd_0__inst_mult_9_41  = CARRY(( !Xd_0__inst_mult_9_6_q  $ (!Xd_0__inst_mult_9_7_q ) ) + ( Xd_0__inst_mult_9_38  ) + ( Xd_0__inst_mult_9_37  ))
// Xd_0__inst_mult_9_42  = SHARE((Xd_0__inst_mult_9_6_q  & Xd_0__inst_mult_9_7_q ))

	.dataa(!Xd_0__inst_mult_9_6_q ),
	.datab(!Xd_0__inst_mult_9_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_37 ),
	.sharein(Xd_0__inst_mult_9_38 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_40 ),
	.cout(Xd_0__inst_mult_9_41 ),
	.shareout(Xd_0__inst_mult_9_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6 (
// Equation(s):
// Xd_0__inst_mult_6_38  = SUM(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_36  ) + ( Xd_0__inst_mult_6_35  ))
// Xd_0__inst_mult_6_39  = CARRY(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_36  ) + ( Xd_0__inst_mult_6_35  ))
// Xd_0__inst_mult_6_40  = SHARE((Xd_0__inst_mult_6_6_q  & Xd_0__inst_mult_6_7_q ))

	.dataa(!Xd_0__inst_mult_6_6_q ),
	.datab(!Xd_0__inst_mult_6_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_35 ),
	.sharein(Xd_0__inst_mult_6_36 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_38 ),
	.cout(Xd_0__inst_mult_6_39 ),
	.shareout(Xd_0__inst_mult_6_40 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7 (
// Equation(s):
// Xd_0__inst_mult_7_39  = SUM(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_7_40  = CARRY(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_7_41  = SHARE((Xd_0__inst_mult_7_6_q  & Xd_0__inst_mult_7_7_q ))

	.dataa(!Xd_0__inst_mult_7_6_q ),
	.datab(!Xd_0__inst_mult_7_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_36 ),
	.sharein(Xd_0__inst_mult_7_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_39 ),
	.cout(Xd_0__inst_mult_7_40 ),
	.shareout(Xd_0__inst_mult_7_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4 (
// Equation(s):
// Xd_0__inst_mult_4_38  = SUM(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_36  ) + ( Xd_0__inst_mult_4_35  ))
// Xd_0__inst_mult_4_39  = CARRY(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_36  ) + ( Xd_0__inst_mult_4_35  ))
// Xd_0__inst_mult_4_40  = SHARE((Xd_0__inst_mult_4_6_q  & Xd_0__inst_mult_4_7_q ))

	.dataa(!Xd_0__inst_mult_4_6_q ),
	.datab(!Xd_0__inst_mult_4_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_35 ),
	.sharein(Xd_0__inst_mult_4_36 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_38 ),
	.cout(Xd_0__inst_mult_4_39 ),
	.shareout(Xd_0__inst_mult_4_40 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5 (
// Equation(s):
// Xd_0__inst_mult_5_39  = SUM(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_5_40  = CARRY(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_5_41  = SHARE((Xd_0__inst_mult_5_6_q  & Xd_0__inst_mult_5_7_q ))

	.dataa(!Xd_0__inst_mult_5_6_q ),
	.datab(!Xd_0__inst_mult_5_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_36 ),
	.sharein(Xd_0__inst_mult_5_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_39 ),
	.cout(Xd_0__inst_mult_5_40 ),
	.shareout(Xd_0__inst_mult_5_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_16 (
// Equation(s):
// Xd_0__inst_mult_2_42  = SUM(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_43  = CARRY(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_44  = SHARE((Xd_0__inst_mult_2_6_q  & Xd_0__inst_mult_2_7_q ))

	.dataa(!Xd_0__inst_mult_2_6_q ),
	.datab(!Xd_0__inst_mult_2_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_40 ),
	.sharein(Xd_0__inst_mult_2_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_42 ),
	.cout(Xd_0__inst_mult_2_43 ),
	.shareout(Xd_0__inst_mult_2_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_16 (
// Equation(s):
// Xd_0__inst_mult_3_42  = SUM(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_mult_3_43  = CARRY(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_mult_3_44  = SHARE((Xd_0__inst_mult_3_6_q  & Xd_0__inst_mult_3_7_q ))

	.dataa(!Xd_0__inst_mult_3_6_q ),
	.datab(!Xd_0__inst_mult_3_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_40 ),
	.sharein(Xd_0__inst_mult_3_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_42 ),
	.cout(Xd_0__inst_mult_3_43 ),
	.shareout(Xd_0__inst_mult_3_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_16 (
// Equation(s):
// Xd_0__inst_mult_0_42  = SUM(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_41  ) + ( Xd_0__inst_mult_0_40  ))
// Xd_0__inst_mult_0_43  = CARRY(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_41  ) + ( Xd_0__inst_mult_0_40  ))
// Xd_0__inst_mult_0_44  = SHARE((Xd_0__inst_mult_0_6_q  & Xd_0__inst_mult_0_7_q ))

	.dataa(!Xd_0__inst_mult_0_6_q ),
	.datab(!Xd_0__inst_mult_0_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_40 ),
	.sharein(Xd_0__inst_mult_0_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_42 ),
	.cout(Xd_0__inst_mult_0_43 ),
	.shareout(Xd_0__inst_mult_0_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_16 (
// Equation(s):
// Xd_0__inst_mult_1_42  = SUM(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_1_43  = CARRY(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_1_44  = SHARE((Xd_0__inst_mult_1_6_q  & Xd_0__inst_mult_1_7_q ))

	.dataa(!Xd_0__inst_mult_1_6_q ),
	.datab(!Xd_0__inst_mult_1_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_40 ),
	.sharein(Xd_0__inst_mult_1_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_42 ),
	.cout(Xd_0__inst_mult_1_43 ),
	.shareout(Xd_0__inst_mult_1_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_28_19 (
// Equation(s):
// Xd_0__inst_mult_28_55  = SUM(( !Xd_0__inst_mult_28_6_q  $ (!Xd_0__inst_mult_28_7_q ) ) + ( Xd_0__inst_mult_28_53  ) + ( Xd_0__inst_mult_28_52  ))
// Xd_0__inst_mult_28_56  = CARRY(( !Xd_0__inst_mult_28_6_q  $ (!Xd_0__inst_mult_28_7_q ) ) + ( Xd_0__inst_mult_28_53  ) + ( Xd_0__inst_mult_28_52  ))
// Xd_0__inst_mult_28_57  = SHARE((Xd_0__inst_mult_28_6_q  & Xd_0__inst_mult_28_7_q ))

	.dataa(!Xd_0__inst_mult_28_6_q ),
	.datab(!Xd_0__inst_mult_28_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_52 ),
	.sharein(Xd_0__inst_mult_28_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_55 ),
	.cout(Xd_0__inst_mult_28_56 ),
	.shareout(Xd_0__inst_mult_28_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_29_17 (
// Equation(s):
// Xd_0__inst_mult_29_47  = SUM(( !Xd_0__inst_mult_29_6_q  $ (!Xd_0__inst_mult_29_7_q ) ) + ( Xd_0__inst_mult_29_45  ) + ( Xd_0__inst_mult_29_44  ))
// Xd_0__inst_mult_29_48  = CARRY(( !Xd_0__inst_mult_29_6_q  $ (!Xd_0__inst_mult_29_7_q ) ) + ( Xd_0__inst_mult_29_45  ) + ( Xd_0__inst_mult_29_44  ))
// Xd_0__inst_mult_29_49  = SHARE((Xd_0__inst_mult_29_6_q  & Xd_0__inst_mult_29_7_q ))

	.dataa(!Xd_0__inst_mult_29_6_q ),
	.datab(!Xd_0__inst_mult_29_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_44 ),
	.sharein(Xd_0__inst_mult_29_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_47 ),
	.cout(Xd_0__inst_mult_29_48 ),
	.shareout(Xd_0__inst_mult_29_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_26_19 (
// Equation(s):
// Xd_0__inst_mult_26_55  = SUM(( !Xd_0__inst_mult_26_6_q  $ (!Xd_0__inst_mult_26_7_q ) ) + ( Xd_0__inst_mult_26_53  ) + ( Xd_0__inst_mult_26_52  ))
// Xd_0__inst_mult_26_56  = CARRY(( !Xd_0__inst_mult_26_6_q  $ (!Xd_0__inst_mult_26_7_q ) ) + ( Xd_0__inst_mult_26_53  ) + ( Xd_0__inst_mult_26_52  ))
// Xd_0__inst_mult_26_57  = SHARE((Xd_0__inst_mult_26_6_q  & Xd_0__inst_mult_26_7_q ))

	.dataa(!Xd_0__inst_mult_26_6_q ),
	.datab(!Xd_0__inst_mult_26_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_52 ),
	.sharein(Xd_0__inst_mult_26_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_55 ),
	.cout(Xd_0__inst_mult_26_56 ),
	.shareout(Xd_0__inst_mult_26_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_27_17 (
// Equation(s):
// Xd_0__inst_mult_27_47  = SUM(( !Xd_0__inst_mult_27_6_q  $ (!Xd_0__inst_mult_27_7_q ) ) + ( Xd_0__inst_mult_27_45  ) + ( Xd_0__inst_mult_27_44  ))
// Xd_0__inst_mult_27_48  = CARRY(( !Xd_0__inst_mult_27_6_q  $ (!Xd_0__inst_mult_27_7_q ) ) + ( Xd_0__inst_mult_27_45  ) + ( Xd_0__inst_mult_27_44  ))
// Xd_0__inst_mult_27_49  = SHARE((Xd_0__inst_mult_27_6_q  & Xd_0__inst_mult_27_7_q ))

	.dataa(!Xd_0__inst_mult_27_6_q ),
	.datab(!Xd_0__inst_mult_27_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_44 ),
	.sharein(Xd_0__inst_mult_27_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_47 ),
	.cout(Xd_0__inst_mult_27_48 ),
	.shareout(Xd_0__inst_mult_27_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_24_19 (
// Equation(s):
// Xd_0__inst_mult_24_55  = SUM(( !Xd_0__inst_mult_24_6_q  $ (!Xd_0__inst_mult_24_7_q ) ) + ( Xd_0__inst_mult_24_53  ) + ( Xd_0__inst_mult_24_52  ))
// Xd_0__inst_mult_24_56  = CARRY(( !Xd_0__inst_mult_24_6_q  $ (!Xd_0__inst_mult_24_7_q ) ) + ( Xd_0__inst_mult_24_53  ) + ( Xd_0__inst_mult_24_52  ))
// Xd_0__inst_mult_24_57  = SHARE((Xd_0__inst_mult_24_6_q  & Xd_0__inst_mult_24_7_q ))

	.dataa(!Xd_0__inst_mult_24_6_q ),
	.datab(!Xd_0__inst_mult_24_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_52 ),
	.sharein(Xd_0__inst_mult_24_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_55 ),
	.cout(Xd_0__inst_mult_24_56 ),
	.shareout(Xd_0__inst_mult_24_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_25_17 (
// Equation(s):
// Xd_0__inst_mult_25_47  = SUM(( !Xd_0__inst_mult_25_6_q  $ (!Xd_0__inst_mult_25_7_q ) ) + ( Xd_0__inst_mult_25_45  ) + ( Xd_0__inst_mult_25_44  ))
// Xd_0__inst_mult_25_48  = CARRY(( !Xd_0__inst_mult_25_6_q  $ (!Xd_0__inst_mult_25_7_q ) ) + ( Xd_0__inst_mult_25_45  ) + ( Xd_0__inst_mult_25_44  ))
// Xd_0__inst_mult_25_49  = SHARE((Xd_0__inst_mult_25_6_q  & Xd_0__inst_mult_25_7_q ))

	.dataa(!Xd_0__inst_mult_25_6_q ),
	.datab(!Xd_0__inst_mult_25_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_44 ),
	.sharein(Xd_0__inst_mult_25_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_47 ),
	.cout(Xd_0__inst_mult_25_48 ),
	.shareout(Xd_0__inst_mult_25_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_22_19 (
// Equation(s):
// Xd_0__inst_mult_22_55  = SUM(( !Xd_0__inst_mult_22_6_q  $ (!Xd_0__inst_mult_22_7_q ) ) + ( Xd_0__inst_mult_22_53  ) + ( Xd_0__inst_mult_22_52  ))
// Xd_0__inst_mult_22_56  = CARRY(( !Xd_0__inst_mult_22_6_q  $ (!Xd_0__inst_mult_22_7_q ) ) + ( Xd_0__inst_mult_22_53  ) + ( Xd_0__inst_mult_22_52  ))
// Xd_0__inst_mult_22_57  = SHARE((Xd_0__inst_mult_22_6_q  & Xd_0__inst_mult_22_7_q ))

	.dataa(!Xd_0__inst_mult_22_6_q ),
	.datab(!Xd_0__inst_mult_22_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_52 ),
	.sharein(Xd_0__inst_mult_22_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_55 ),
	.cout(Xd_0__inst_mult_22_56 ),
	.shareout(Xd_0__inst_mult_22_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_23_19 (
// Equation(s):
// Xd_0__inst_mult_23_55  = SUM(( !Xd_0__inst_mult_23_6_q  $ (!Xd_0__inst_mult_23_7_q ) ) + ( Xd_0__inst_mult_23_53  ) + ( Xd_0__inst_mult_23_52  ))
// Xd_0__inst_mult_23_56  = CARRY(( !Xd_0__inst_mult_23_6_q  $ (!Xd_0__inst_mult_23_7_q ) ) + ( Xd_0__inst_mult_23_53  ) + ( Xd_0__inst_mult_23_52  ))
// Xd_0__inst_mult_23_57  = SHARE((Xd_0__inst_mult_23_6_q  & Xd_0__inst_mult_23_7_q ))

	.dataa(!Xd_0__inst_mult_23_6_q ),
	.datab(!Xd_0__inst_mult_23_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_52 ),
	.sharein(Xd_0__inst_mult_23_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_55 ),
	.cout(Xd_0__inst_mult_23_56 ),
	.shareout(Xd_0__inst_mult_23_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_20_19 (
// Equation(s):
// Xd_0__inst_mult_20_55  = SUM(( !Xd_0__inst_mult_20_6_q  $ (!Xd_0__inst_mult_20_7_q ) ) + ( Xd_0__inst_mult_20_53  ) + ( Xd_0__inst_mult_20_52  ))
// Xd_0__inst_mult_20_56  = CARRY(( !Xd_0__inst_mult_20_6_q  $ (!Xd_0__inst_mult_20_7_q ) ) + ( Xd_0__inst_mult_20_53  ) + ( Xd_0__inst_mult_20_52  ))
// Xd_0__inst_mult_20_57  = SHARE((Xd_0__inst_mult_20_6_q  & Xd_0__inst_mult_20_7_q ))

	.dataa(!Xd_0__inst_mult_20_6_q ),
	.datab(!Xd_0__inst_mult_20_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_52 ),
	.sharein(Xd_0__inst_mult_20_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_55 ),
	.cout(Xd_0__inst_mult_20_56 ),
	.shareout(Xd_0__inst_mult_20_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_21 (
// Equation(s):
// Xd_0__inst_mult_21_40  = SUM(( !Xd_0__inst_mult_21_6_q  $ (!Xd_0__inst_mult_21_7_q ) ) + ( Xd_0__inst_mult_21_38  ) + ( Xd_0__inst_mult_21_37  ))
// Xd_0__inst_mult_21_41  = CARRY(( !Xd_0__inst_mult_21_6_q  $ (!Xd_0__inst_mult_21_7_q ) ) + ( Xd_0__inst_mult_21_38  ) + ( Xd_0__inst_mult_21_37  ))
// Xd_0__inst_mult_21_42  = SHARE((Xd_0__inst_mult_21_6_q  & Xd_0__inst_mult_21_7_q ))

	.dataa(!Xd_0__inst_mult_21_6_q ),
	.datab(!Xd_0__inst_mult_21_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_37 ),
	.sharein(Xd_0__inst_mult_21_38 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_40 ),
	.cout(Xd_0__inst_mult_21_41 ),
	.shareout(Xd_0__inst_mult_21_42 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_18 (
// Equation(s):
// Xd_0__inst_mult_18_39  = SUM(( !Xd_0__inst_mult_18_6_q  $ (!Xd_0__inst_mult_18_7_q ) ) + ( Xd_0__inst_mult_18_37  ) + ( Xd_0__inst_mult_18_36  ))
// Xd_0__inst_mult_18_40  = CARRY(( !Xd_0__inst_mult_18_6_q  $ (!Xd_0__inst_mult_18_7_q ) ) + ( Xd_0__inst_mult_18_37  ) + ( Xd_0__inst_mult_18_36  ))
// Xd_0__inst_mult_18_41  = SHARE((Xd_0__inst_mult_18_6_q  & Xd_0__inst_mult_18_7_q ))

	.dataa(!Xd_0__inst_mult_18_6_q ),
	.datab(!Xd_0__inst_mult_18_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_36 ),
	.sharein(Xd_0__inst_mult_18_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_39 ),
	.cout(Xd_0__inst_mult_18_40 ),
	.shareout(Xd_0__inst_mult_18_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_19_18 (
// Equation(s):
// Xd_0__inst_mult_19_51  = SUM(( !Xd_0__inst_mult_19_6_q  $ (!Xd_0__inst_mult_19_7_q ) ) + ( Xd_0__inst_mult_19_49  ) + ( Xd_0__inst_mult_19_48  ))
// Xd_0__inst_mult_19_52  = CARRY(( !Xd_0__inst_mult_19_6_q  $ (!Xd_0__inst_mult_19_7_q ) ) + ( Xd_0__inst_mult_19_49  ) + ( Xd_0__inst_mult_19_48  ))
// Xd_0__inst_mult_19_53  = SHARE((Xd_0__inst_mult_19_6_q  & Xd_0__inst_mult_19_7_q ))

	.dataa(!Xd_0__inst_mult_19_6_q ),
	.datab(!Xd_0__inst_mult_19_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_48 ),
	.sharein(Xd_0__inst_mult_19_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_51 ),
	.cout(Xd_0__inst_mult_19_52 ),
	.shareout(Xd_0__inst_mult_19_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_16_16 (
// Equation(s):
// Xd_0__inst_mult_16_42  = SUM(( !Xd_0__inst_mult_16_8_q  $ (!Xd_0__inst_mult_16_9_q  $ (((Xd_0__inst_mult_16_4_q  & Xd_0__inst_mult_16_10_q )))) ) + ( Xd_0__inst_mult_16_41  ) + ( Xd_0__inst_mult_16_40  ))
// Xd_0__inst_mult_16_43  = CARRY(( !Xd_0__inst_mult_16_8_q  $ (!Xd_0__inst_mult_16_9_q  $ (((Xd_0__inst_mult_16_4_q  & Xd_0__inst_mult_16_10_q )))) ) + ( Xd_0__inst_mult_16_41  ) + ( Xd_0__inst_mult_16_40  ))
// Xd_0__inst_mult_16_44  = SHARE((!Xd_0__inst_mult_16_8_q  & (Xd_0__inst_mult_16_9_q  & (Xd_0__inst_mult_16_4_q  & Xd_0__inst_mult_16_10_q ))) # (Xd_0__inst_mult_16_8_q  & (((Xd_0__inst_mult_16_4_q  & Xd_0__inst_mult_16_10_q )) # (Xd_0__inst_mult_16_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_16_8_q ),
	.datab(!Xd_0__inst_mult_16_9_q ),
	.datac(!Xd_0__inst_mult_16_4_q ),
	.datad(!Xd_0__inst_mult_16_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_40 ),
	.sharein(Xd_0__inst_mult_16_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_42 ),
	.cout(Xd_0__inst_mult_16_43 ),
	.shareout(Xd_0__inst_mult_16_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_17_16 (
// Equation(s):
// Xd_0__inst_mult_17_43  = SUM(( !Xd_0__inst_mult_17_8_q  $ (!Xd_0__inst_mult_17_9_q  $ (((Xd_0__inst_mult_17_4_q  & Xd_0__inst_mult_17_10_q )))) ) + ( Xd_0__inst_mult_17_42  ) + ( Xd_0__inst_mult_17_41  ))
// Xd_0__inst_mult_17_44  = CARRY(( !Xd_0__inst_mult_17_8_q  $ (!Xd_0__inst_mult_17_9_q  $ (((Xd_0__inst_mult_17_4_q  & Xd_0__inst_mult_17_10_q )))) ) + ( Xd_0__inst_mult_17_42  ) + ( Xd_0__inst_mult_17_41  ))
// Xd_0__inst_mult_17_45  = SHARE((!Xd_0__inst_mult_17_8_q  & (Xd_0__inst_mult_17_9_q  & (Xd_0__inst_mult_17_4_q  & Xd_0__inst_mult_17_10_q ))) # (Xd_0__inst_mult_17_8_q  & (((Xd_0__inst_mult_17_4_q  & Xd_0__inst_mult_17_10_q )) # (Xd_0__inst_mult_17_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_17_8_q ),
	.datab(!Xd_0__inst_mult_17_9_q ),
	.datac(!Xd_0__inst_mult_17_4_q ),
	.datad(!Xd_0__inst_mult_17_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_41 ),
	.sharein(Xd_0__inst_mult_17_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_43 ),
	.cout(Xd_0__inst_mult_17_44 ),
	.shareout(Xd_0__inst_mult_17_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_14_16 (
// Equation(s):
// Xd_0__inst_mult_14_42  = SUM(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q  $ (((Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_10_q )))) ) + ( Xd_0__inst_mult_14_41  ) + ( Xd_0__inst_mult_14_40  ))
// Xd_0__inst_mult_14_43  = CARRY(( !Xd_0__inst_mult_14_8_q  $ (!Xd_0__inst_mult_14_9_q  $ (((Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_10_q )))) ) + ( Xd_0__inst_mult_14_41  ) + ( Xd_0__inst_mult_14_40  ))
// Xd_0__inst_mult_14_44  = SHARE((!Xd_0__inst_mult_14_8_q  & (Xd_0__inst_mult_14_9_q  & (Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_10_q ))) # (Xd_0__inst_mult_14_8_q  & (((Xd_0__inst_mult_14_4_q  & Xd_0__inst_mult_14_10_q )) # (Xd_0__inst_mult_14_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_14_8_q ),
	.datab(!Xd_0__inst_mult_14_9_q ),
	.datac(!Xd_0__inst_mult_14_4_q ),
	.datad(!Xd_0__inst_mult_14_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_40 ),
	.sharein(Xd_0__inst_mult_14_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_42 ),
	.cout(Xd_0__inst_mult_14_43 ),
	.shareout(Xd_0__inst_mult_14_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_15_16 (
// Equation(s):
// Xd_0__inst_mult_15_43  = SUM(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q  $ (((Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_10_q )))) ) + ( Xd_0__inst_mult_15_42  ) + ( Xd_0__inst_mult_15_41  ))
// Xd_0__inst_mult_15_44  = CARRY(( !Xd_0__inst_mult_15_8_q  $ (!Xd_0__inst_mult_15_9_q  $ (((Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_10_q )))) ) + ( Xd_0__inst_mult_15_42  ) + ( Xd_0__inst_mult_15_41  ))
// Xd_0__inst_mult_15_45  = SHARE((!Xd_0__inst_mult_15_8_q  & (Xd_0__inst_mult_15_9_q  & (Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_10_q ))) # (Xd_0__inst_mult_15_8_q  & (((Xd_0__inst_mult_15_4_q  & Xd_0__inst_mult_15_10_q )) # (Xd_0__inst_mult_15_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_15_8_q ),
	.datab(!Xd_0__inst_mult_15_9_q ),
	.datac(!Xd_0__inst_mult_15_4_q ),
	.datad(!Xd_0__inst_mult_15_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_41 ),
	.sharein(Xd_0__inst_mult_15_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_43 ),
	.cout(Xd_0__inst_mult_15_44 ),
	.shareout(Xd_0__inst_mult_15_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_12_16 (
// Equation(s):
// Xd_0__inst_mult_12_42  = SUM(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q  $ (((Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_10_q )))) ) + ( Xd_0__inst_mult_12_41  ) + ( Xd_0__inst_mult_12_40  ))
// Xd_0__inst_mult_12_43  = CARRY(( !Xd_0__inst_mult_12_8_q  $ (!Xd_0__inst_mult_12_9_q  $ (((Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_10_q )))) ) + ( Xd_0__inst_mult_12_41  ) + ( Xd_0__inst_mult_12_40  ))
// Xd_0__inst_mult_12_44  = SHARE((!Xd_0__inst_mult_12_8_q  & (Xd_0__inst_mult_12_9_q  & (Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_10_q ))) # (Xd_0__inst_mult_12_8_q  & (((Xd_0__inst_mult_12_4_q  & Xd_0__inst_mult_12_10_q )) # (Xd_0__inst_mult_12_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_12_8_q ),
	.datab(!Xd_0__inst_mult_12_9_q ),
	.datac(!Xd_0__inst_mult_12_4_q ),
	.datad(!Xd_0__inst_mult_12_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_40 ),
	.sharein(Xd_0__inst_mult_12_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_42 ),
	.cout(Xd_0__inst_mult_12_43 ),
	.shareout(Xd_0__inst_mult_12_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_13_16 (
// Equation(s):
// Xd_0__inst_mult_13_43  = SUM(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q  $ (((Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_10_q )))) ) + ( Xd_0__inst_mult_13_42  ) + ( Xd_0__inst_mult_13_41  ))
// Xd_0__inst_mult_13_44  = CARRY(( !Xd_0__inst_mult_13_8_q  $ (!Xd_0__inst_mult_13_9_q  $ (((Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_10_q )))) ) + ( Xd_0__inst_mult_13_42  ) + ( Xd_0__inst_mult_13_41  ))
// Xd_0__inst_mult_13_45  = SHARE((!Xd_0__inst_mult_13_8_q  & (Xd_0__inst_mult_13_9_q  & (Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_10_q ))) # (Xd_0__inst_mult_13_8_q  & (((Xd_0__inst_mult_13_4_q  & Xd_0__inst_mult_13_10_q )) # (Xd_0__inst_mult_13_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_13_8_q ),
	.datab(!Xd_0__inst_mult_13_9_q ),
	.datac(!Xd_0__inst_mult_13_4_q ),
	.datad(!Xd_0__inst_mult_13_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_41 ),
	.sharein(Xd_0__inst_mult_13_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_43 ),
	.cout(Xd_0__inst_mult_13_44 ),
	.shareout(Xd_0__inst_mult_13_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_10_16 (
// Equation(s):
// Xd_0__inst_mult_10_42  = SUM(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q  $ (((Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_10_q )))) ) + ( Xd_0__inst_mult_10_41  ) + ( Xd_0__inst_mult_10_40  ))
// Xd_0__inst_mult_10_43  = CARRY(( !Xd_0__inst_mult_10_8_q  $ (!Xd_0__inst_mult_10_9_q  $ (((Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_10_q )))) ) + ( Xd_0__inst_mult_10_41  ) + ( Xd_0__inst_mult_10_40  ))
// Xd_0__inst_mult_10_44  = SHARE((!Xd_0__inst_mult_10_8_q  & (Xd_0__inst_mult_10_9_q  & (Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_10_q ))) # (Xd_0__inst_mult_10_8_q  & (((Xd_0__inst_mult_10_4_q  & Xd_0__inst_mult_10_10_q )) # (Xd_0__inst_mult_10_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_10_8_q ),
	.datab(!Xd_0__inst_mult_10_9_q ),
	.datac(!Xd_0__inst_mult_10_4_q ),
	.datad(!Xd_0__inst_mult_10_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_40 ),
	.sharein(Xd_0__inst_mult_10_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_42 ),
	.cout(Xd_0__inst_mult_10_43 ),
	.shareout(Xd_0__inst_mult_10_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_11_18 (
// Equation(s):
// Xd_0__inst_mult_11_51  = SUM(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q  $ (((Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_10_q )))) ) + ( Xd_0__inst_mult_11_49  ) + ( Xd_0__inst_mult_11_48  ))
// Xd_0__inst_mult_11_52  = CARRY(( !Xd_0__inst_mult_11_8_q  $ (!Xd_0__inst_mult_11_9_q  $ (((Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_10_q )))) ) + ( Xd_0__inst_mult_11_49  ) + ( Xd_0__inst_mult_11_48  ))
// Xd_0__inst_mult_11_53  = SHARE((!Xd_0__inst_mult_11_8_q  & (Xd_0__inst_mult_11_9_q  & (Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_10_q ))) # (Xd_0__inst_mult_11_8_q  & (((Xd_0__inst_mult_11_4_q  & Xd_0__inst_mult_11_10_q )) # (Xd_0__inst_mult_11_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_11_8_q ),
	.datab(!Xd_0__inst_mult_11_9_q ),
	.datac(!Xd_0__inst_mult_11_4_q ),
	.datad(!Xd_0__inst_mult_11_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_48 ),
	.sharein(Xd_0__inst_mult_11_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_51 ),
	.cout(Xd_0__inst_mult_11_52 ),
	.shareout(Xd_0__inst_mult_11_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_8_16 (
// Equation(s):
// Xd_0__inst_mult_8_42  = SUM(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q  $ (((Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_10_q )))) ) + ( Xd_0__inst_mult_8_41  ) + ( Xd_0__inst_mult_8_40  ))
// Xd_0__inst_mult_8_43  = CARRY(( !Xd_0__inst_mult_8_8_q  $ (!Xd_0__inst_mult_8_9_q  $ (((Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_10_q )))) ) + ( Xd_0__inst_mult_8_41  ) + ( Xd_0__inst_mult_8_40  ))
// Xd_0__inst_mult_8_44  = SHARE((!Xd_0__inst_mult_8_8_q  & (Xd_0__inst_mult_8_9_q  & (Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_10_q ))) # (Xd_0__inst_mult_8_8_q  & (((Xd_0__inst_mult_8_4_q  & Xd_0__inst_mult_8_10_q )) # (Xd_0__inst_mult_8_9_q ))))

	.dataa(!Xd_0__inst_mult_8_8_q ),
	.datab(!Xd_0__inst_mult_8_9_q ),
	.datac(!Xd_0__inst_mult_8_4_q ),
	.datad(!Xd_0__inst_mult_8_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_40 ),
	.sharein(Xd_0__inst_mult_8_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_42 ),
	.cout(Xd_0__inst_mult_8_43 ),
	.shareout(Xd_0__inst_mult_8_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_9_16 (
// Equation(s):
// Xd_0__inst_mult_9_43  = SUM(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q  $ (((Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_10_q )))) ) + ( Xd_0__inst_mult_9_42  ) + ( Xd_0__inst_mult_9_41  ))
// Xd_0__inst_mult_9_44  = CARRY(( !Xd_0__inst_mult_9_8_q  $ (!Xd_0__inst_mult_9_9_q  $ (((Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_10_q )))) ) + ( Xd_0__inst_mult_9_42  ) + ( Xd_0__inst_mult_9_41  ))
// Xd_0__inst_mult_9_45  = SHARE((!Xd_0__inst_mult_9_8_q  & (Xd_0__inst_mult_9_9_q  & (Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_10_q ))) # (Xd_0__inst_mult_9_8_q  & (((Xd_0__inst_mult_9_4_q  & Xd_0__inst_mult_9_10_q )) # (Xd_0__inst_mult_9_9_q ))))

	.dataa(!Xd_0__inst_mult_9_8_q ),
	.datab(!Xd_0__inst_mult_9_9_q ),
	.datac(!Xd_0__inst_mult_9_4_q ),
	.datad(!Xd_0__inst_mult_9_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_41 ),
	.sharein(Xd_0__inst_mult_9_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_43 ),
	.cout(Xd_0__inst_mult_9_44 ),
	.shareout(Xd_0__inst_mult_9_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_16 (
// Equation(s):
// Xd_0__inst_mult_6_41  = SUM(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q  $ (((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_10_q )))) ) + ( Xd_0__inst_mult_6_40  ) + ( Xd_0__inst_mult_6_39  ))
// Xd_0__inst_mult_6_42  = CARRY(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q  $ (((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_10_q )))) ) + ( Xd_0__inst_mult_6_40  ) + ( Xd_0__inst_mult_6_39  ))
// Xd_0__inst_mult_6_43  = SHARE((!Xd_0__inst_mult_6_8_q  & (Xd_0__inst_mult_6_9_q  & (Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_10_q ))) # (Xd_0__inst_mult_6_8_q  & (((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_10_q )) # (Xd_0__inst_mult_6_9_q ))))

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(!Xd_0__inst_mult_6_4_q ),
	.datad(!Xd_0__inst_mult_6_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_39 ),
	.sharein(Xd_0__inst_mult_6_40 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_41 ),
	.cout(Xd_0__inst_mult_6_42 ),
	.shareout(Xd_0__inst_mult_6_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_16 (
// Equation(s):
// Xd_0__inst_mult_7_42  = SUM(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q  $ (((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_10_q )))) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_7_43  = CARRY(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q  $ (((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_10_q )))) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_7_44  = SHARE((!Xd_0__inst_mult_7_8_q  & (Xd_0__inst_mult_7_9_q  & (Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_10_q ))) # (Xd_0__inst_mult_7_8_q  & (((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_10_q )) # (Xd_0__inst_mult_7_9_q ))))

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(!Xd_0__inst_mult_7_4_q ),
	.datad(!Xd_0__inst_mult_7_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_40 ),
	.sharein(Xd_0__inst_mult_7_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_42 ),
	.cout(Xd_0__inst_mult_7_43 ),
	.shareout(Xd_0__inst_mult_7_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_16 (
// Equation(s):
// Xd_0__inst_mult_4_41  = SUM(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q  $ (((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_10_q )))) ) + ( Xd_0__inst_mult_4_40  ) + ( Xd_0__inst_mult_4_39  ))
// Xd_0__inst_mult_4_42  = CARRY(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q  $ (((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_10_q )))) ) + ( Xd_0__inst_mult_4_40  ) + ( Xd_0__inst_mult_4_39  ))
// Xd_0__inst_mult_4_43  = SHARE((!Xd_0__inst_mult_4_8_q  & (Xd_0__inst_mult_4_9_q  & (Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_10_q ))) # (Xd_0__inst_mult_4_8_q  & (((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_10_q )) # (Xd_0__inst_mult_4_9_q ))))

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(!Xd_0__inst_mult_4_4_q ),
	.datad(!Xd_0__inst_mult_4_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_39 ),
	.sharein(Xd_0__inst_mult_4_40 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_41 ),
	.cout(Xd_0__inst_mult_4_42 ),
	.shareout(Xd_0__inst_mult_4_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_16 (
// Equation(s):
// Xd_0__inst_mult_5_42  = SUM(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q  $ (((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_10_q )))) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_5_43  = CARRY(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q  $ (((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_10_q )))) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_5_44  = SHARE((!Xd_0__inst_mult_5_8_q  & (Xd_0__inst_mult_5_9_q  & (Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_10_q ))) # (Xd_0__inst_mult_5_8_q  & (((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_10_q )) # (Xd_0__inst_mult_5_9_q ))))

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(!Xd_0__inst_mult_5_4_q ),
	.datad(!Xd_0__inst_mult_5_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_40 ),
	.sharein(Xd_0__inst_mult_5_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_42 ),
	.cout(Xd_0__inst_mult_5_43 ),
	.shareout(Xd_0__inst_mult_5_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_17 (
// Equation(s):
// Xd_0__inst_mult_2_46  = SUM(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q  $ (((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_10_q )))) ) + ( Xd_0__inst_mult_2_44  ) + ( Xd_0__inst_mult_2_43  ))
// Xd_0__inst_mult_2_47  = CARRY(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q  $ (((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_10_q )))) ) + ( Xd_0__inst_mult_2_44  ) + ( Xd_0__inst_mult_2_43  ))
// Xd_0__inst_mult_2_48  = SHARE((!Xd_0__inst_mult_2_8_q  & (Xd_0__inst_mult_2_9_q  & (Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_10_q ))) # (Xd_0__inst_mult_2_8_q  & (((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_10_q )) # (Xd_0__inst_mult_2_9_q ))))

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(!Xd_0__inst_mult_2_4_q ),
	.datad(!Xd_0__inst_mult_2_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_43 ),
	.sharein(Xd_0__inst_mult_2_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_46 ),
	.cout(Xd_0__inst_mult_2_47 ),
	.shareout(Xd_0__inst_mult_2_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_17 (
// Equation(s):
// Xd_0__inst_mult_3_46  = SUM(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q  $ (((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_10_q )))) ) + ( Xd_0__inst_mult_3_44  ) + ( Xd_0__inst_mult_3_43  ))
// Xd_0__inst_mult_3_47  = CARRY(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q  $ (((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_10_q )))) ) + ( Xd_0__inst_mult_3_44  ) + ( Xd_0__inst_mult_3_43  ))
// Xd_0__inst_mult_3_48  = SHARE((!Xd_0__inst_mult_3_8_q  & (Xd_0__inst_mult_3_9_q  & (Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_10_q ))) # (Xd_0__inst_mult_3_8_q  & (((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_10_q )) # (Xd_0__inst_mult_3_9_q ))))

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(!Xd_0__inst_mult_3_4_q ),
	.datad(!Xd_0__inst_mult_3_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_43 ),
	.sharein(Xd_0__inst_mult_3_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_46 ),
	.cout(Xd_0__inst_mult_3_47 ),
	.shareout(Xd_0__inst_mult_3_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_17 (
// Equation(s):
// Xd_0__inst_mult_0_46  = SUM(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q  $ (((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_10_q )))) ) + ( Xd_0__inst_mult_0_44  ) + ( Xd_0__inst_mult_0_43  ))
// Xd_0__inst_mult_0_47  = CARRY(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q  $ (((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_10_q )))) ) + ( Xd_0__inst_mult_0_44  ) + ( Xd_0__inst_mult_0_43  ))
// Xd_0__inst_mult_0_48  = SHARE((!Xd_0__inst_mult_0_8_q  & (Xd_0__inst_mult_0_9_q  & (Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_10_q ))) # (Xd_0__inst_mult_0_8_q  & (((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_10_q )) # (Xd_0__inst_mult_0_9_q ))))

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(!Xd_0__inst_mult_0_4_q ),
	.datad(!Xd_0__inst_mult_0_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_43 ),
	.sharein(Xd_0__inst_mult_0_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_46 ),
	.cout(Xd_0__inst_mult_0_47 ),
	.shareout(Xd_0__inst_mult_0_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_17 (
// Equation(s):
// Xd_0__inst_mult_1_46  = SUM(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q  $ (((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_10_q )))) ) + ( Xd_0__inst_mult_1_44  ) + ( Xd_0__inst_mult_1_43  ))
// Xd_0__inst_mult_1_47  = CARRY(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q  $ (((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_10_q )))) ) + ( Xd_0__inst_mult_1_44  ) + ( Xd_0__inst_mult_1_43  ))
// Xd_0__inst_mult_1_48  = SHARE((!Xd_0__inst_mult_1_8_q  & (Xd_0__inst_mult_1_9_q  & (Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_10_q ))) # (Xd_0__inst_mult_1_8_q  & (((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_10_q )) # (Xd_0__inst_mult_1_9_q ))))

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(!Xd_0__inst_mult_1_4_q ),
	.datad(!Xd_0__inst_mult_1_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_43 ),
	.sharein(Xd_0__inst_mult_1_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_46 ),
	.cout(Xd_0__inst_mult_1_47 ),
	.shareout(Xd_0__inst_mult_1_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_28_20 (
// Equation(s):
// Xd_0__inst_mult_28_59  = SUM(( !Xd_0__inst_mult_28_8_q  $ (!Xd_0__inst_mult_28_9_q  $ (((Xd_0__inst_mult_28_4_q  & Xd_0__inst_mult_28_10_q )))) ) + ( Xd_0__inst_mult_28_57  ) + ( Xd_0__inst_mult_28_56  ))
// Xd_0__inst_mult_28_60  = CARRY(( !Xd_0__inst_mult_28_8_q  $ (!Xd_0__inst_mult_28_9_q  $ (((Xd_0__inst_mult_28_4_q  & Xd_0__inst_mult_28_10_q )))) ) + ( Xd_0__inst_mult_28_57  ) + ( Xd_0__inst_mult_28_56  ))
// Xd_0__inst_mult_28_61  = SHARE((!Xd_0__inst_mult_28_8_q  & (Xd_0__inst_mult_28_9_q  & (Xd_0__inst_mult_28_4_q  & Xd_0__inst_mult_28_10_q ))) # (Xd_0__inst_mult_28_8_q  & (((Xd_0__inst_mult_28_4_q  & Xd_0__inst_mult_28_10_q )) # (Xd_0__inst_mult_28_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_28_8_q ),
	.datab(!Xd_0__inst_mult_28_9_q ),
	.datac(!Xd_0__inst_mult_28_4_q ),
	.datad(!Xd_0__inst_mult_28_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_56 ),
	.sharein(Xd_0__inst_mult_28_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_59 ),
	.cout(Xd_0__inst_mult_28_60 ),
	.shareout(Xd_0__inst_mult_28_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_29_18 (
// Equation(s):
// Xd_0__inst_mult_29_51  = SUM(( !Xd_0__inst_mult_29_8_q  $ (!Xd_0__inst_mult_29_9_q  $ (((Xd_0__inst_mult_29_4_q  & Xd_0__inst_mult_29_10_q )))) ) + ( Xd_0__inst_mult_29_49  ) + ( Xd_0__inst_mult_29_48  ))
// Xd_0__inst_mult_29_52  = CARRY(( !Xd_0__inst_mult_29_8_q  $ (!Xd_0__inst_mult_29_9_q  $ (((Xd_0__inst_mult_29_4_q  & Xd_0__inst_mult_29_10_q )))) ) + ( Xd_0__inst_mult_29_49  ) + ( Xd_0__inst_mult_29_48  ))
// Xd_0__inst_mult_29_53  = SHARE((!Xd_0__inst_mult_29_8_q  & (Xd_0__inst_mult_29_9_q  & (Xd_0__inst_mult_29_4_q  & Xd_0__inst_mult_29_10_q ))) # (Xd_0__inst_mult_29_8_q  & (((Xd_0__inst_mult_29_4_q  & Xd_0__inst_mult_29_10_q )) # (Xd_0__inst_mult_29_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_29_8_q ),
	.datab(!Xd_0__inst_mult_29_9_q ),
	.datac(!Xd_0__inst_mult_29_4_q ),
	.datad(!Xd_0__inst_mult_29_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_48 ),
	.sharein(Xd_0__inst_mult_29_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_51 ),
	.cout(Xd_0__inst_mult_29_52 ),
	.shareout(Xd_0__inst_mult_29_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_26_20 (
// Equation(s):
// Xd_0__inst_mult_26_59  = SUM(( !Xd_0__inst_mult_26_8_q  $ (!Xd_0__inst_mult_26_9_q  $ (((Xd_0__inst_mult_26_4_q  & Xd_0__inst_mult_26_10_q )))) ) + ( Xd_0__inst_mult_26_57  ) + ( Xd_0__inst_mult_26_56  ))
// Xd_0__inst_mult_26_60  = CARRY(( !Xd_0__inst_mult_26_8_q  $ (!Xd_0__inst_mult_26_9_q  $ (((Xd_0__inst_mult_26_4_q  & Xd_0__inst_mult_26_10_q )))) ) + ( Xd_0__inst_mult_26_57  ) + ( Xd_0__inst_mult_26_56  ))
// Xd_0__inst_mult_26_61  = SHARE((!Xd_0__inst_mult_26_8_q  & (Xd_0__inst_mult_26_9_q  & (Xd_0__inst_mult_26_4_q  & Xd_0__inst_mult_26_10_q ))) # (Xd_0__inst_mult_26_8_q  & (((Xd_0__inst_mult_26_4_q  & Xd_0__inst_mult_26_10_q )) # (Xd_0__inst_mult_26_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_26_8_q ),
	.datab(!Xd_0__inst_mult_26_9_q ),
	.datac(!Xd_0__inst_mult_26_4_q ),
	.datad(!Xd_0__inst_mult_26_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_56 ),
	.sharein(Xd_0__inst_mult_26_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_59 ),
	.cout(Xd_0__inst_mult_26_60 ),
	.shareout(Xd_0__inst_mult_26_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_27_18 (
// Equation(s):
// Xd_0__inst_mult_27_51  = SUM(( !Xd_0__inst_mult_27_8_q  $ (!Xd_0__inst_mult_27_9_q  $ (((Xd_0__inst_mult_27_4_q  & Xd_0__inst_mult_27_10_q )))) ) + ( Xd_0__inst_mult_27_49  ) + ( Xd_0__inst_mult_27_48  ))
// Xd_0__inst_mult_27_52  = CARRY(( !Xd_0__inst_mult_27_8_q  $ (!Xd_0__inst_mult_27_9_q  $ (((Xd_0__inst_mult_27_4_q  & Xd_0__inst_mult_27_10_q )))) ) + ( Xd_0__inst_mult_27_49  ) + ( Xd_0__inst_mult_27_48  ))
// Xd_0__inst_mult_27_53  = SHARE((!Xd_0__inst_mult_27_8_q  & (Xd_0__inst_mult_27_9_q  & (Xd_0__inst_mult_27_4_q  & Xd_0__inst_mult_27_10_q ))) # (Xd_0__inst_mult_27_8_q  & (((Xd_0__inst_mult_27_4_q  & Xd_0__inst_mult_27_10_q )) # (Xd_0__inst_mult_27_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_27_8_q ),
	.datab(!Xd_0__inst_mult_27_9_q ),
	.datac(!Xd_0__inst_mult_27_4_q ),
	.datad(!Xd_0__inst_mult_27_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_48 ),
	.sharein(Xd_0__inst_mult_27_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_51 ),
	.cout(Xd_0__inst_mult_27_52 ),
	.shareout(Xd_0__inst_mult_27_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_24_20 (
// Equation(s):
// Xd_0__inst_mult_24_59  = SUM(( !Xd_0__inst_mult_24_8_q  $ (!Xd_0__inst_mult_24_9_q  $ (((Xd_0__inst_mult_24_4_q  & Xd_0__inst_mult_24_10_q )))) ) + ( Xd_0__inst_mult_24_57  ) + ( Xd_0__inst_mult_24_56  ))
// Xd_0__inst_mult_24_60  = CARRY(( !Xd_0__inst_mult_24_8_q  $ (!Xd_0__inst_mult_24_9_q  $ (((Xd_0__inst_mult_24_4_q  & Xd_0__inst_mult_24_10_q )))) ) + ( Xd_0__inst_mult_24_57  ) + ( Xd_0__inst_mult_24_56  ))
// Xd_0__inst_mult_24_61  = SHARE((!Xd_0__inst_mult_24_8_q  & (Xd_0__inst_mult_24_9_q  & (Xd_0__inst_mult_24_4_q  & Xd_0__inst_mult_24_10_q ))) # (Xd_0__inst_mult_24_8_q  & (((Xd_0__inst_mult_24_4_q  & Xd_0__inst_mult_24_10_q )) # (Xd_0__inst_mult_24_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_24_8_q ),
	.datab(!Xd_0__inst_mult_24_9_q ),
	.datac(!Xd_0__inst_mult_24_4_q ),
	.datad(!Xd_0__inst_mult_24_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_56 ),
	.sharein(Xd_0__inst_mult_24_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_59 ),
	.cout(Xd_0__inst_mult_24_60 ),
	.shareout(Xd_0__inst_mult_24_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_25_18 (
// Equation(s):
// Xd_0__inst_mult_25_51  = SUM(( !Xd_0__inst_mult_25_8_q  $ (!Xd_0__inst_mult_25_9_q  $ (((Xd_0__inst_mult_25_4_q  & Xd_0__inst_mult_25_10_q )))) ) + ( Xd_0__inst_mult_25_49  ) + ( Xd_0__inst_mult_25_48  ))
// Xd_0__inst_mult_25_52  = CARRY(( !Xd_0__inst_mult_25_8_q  $ (!Xd_0__inst_mult_25_9_q  $ (((Xd_0__inst_mult_25_4_q  & Xd_0__inst_mult_25_10_q )))) ) + ( Xd_0__inst_mult_25_49  ) + ( Xd_0__inst_mult_25_48  ))
// Xd_0__inst_mult_25_53  = SHARE((!Xd_0__inst_mult_25_8_q  & (Xd_0__inst_mult_25_9_q  & (Xd_0__inst_mult_25_4_q  & Xd_0__inst_mult_25_10_q ))) # (Xd_0__inst_mult_25_8_q  & (((Xd_0__inst_mult_25_4_q  & Xd_0__inst_mult_25_10_q )) # (Xd_0__inst_mult_25_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_25_8_q ),
	.datab(!Xd_0__inst_mult_25_9_q ),
	.datac(!Xd_0__inst_mult_25_4_q ),
	.datad(!Xd_0__inst_mult_25_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_48 ),
	.sharein(Xd_0__inst_mult_25_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_51 ),
	.cout(Xd_0__inst_mult_25_52 ),
	.shareout(Xd_0__inst_mult_25_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_22_20 (
// Equation(s):
// Xd_0__inst_mult_22_59  = SUM(( !Xd_0__inst_mult_22_8_q  $ (!Xd_0__inst_mult_22_9_q  $ (((Xd_0__inst_mult_22_4_q  & Xd_0__inst_mult_22_10_q )))) ) + ( Xd_0__inst_mult_22_57  ) + ( Xd_0__inst_mult_22_56  ))
// Xd_0__inst_mult_22_60  = CARRY(( !Xd_0__inst_mult_22_8_q  $ (!Xd_0__inst_mult_22_9_q  $ (((Xd_0__inst_mult_22_4_q  & Xd_0__inst_mult_22_10_q )))) ) + ( Xd_0__inst_mult_22_57  ) + ( Xd_0__inst_mult_22_56  ))
// Xd_0__inst_mult_22_61  = SHARE((!Xd_0__inst_mult_22_8_q  & (Xd_0__inst_mult_22_9_q  & (Xd_0__inst_mult_22_4_q  & Xd_0__inst_mult_22_10_q ))) # (Xd_0__inst_mult_22_8_q  & (((Xd_0__inst_mult_22_4_q  & Xd_0__inst_mult_22_10_q )) # (Xd_0__inst_mult_22_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_22_8_q ),
	.datab(!Xd_0__inst_mult_22_9_q ),
	.datac(!Xd_0__inst_mult_22_4_q ),
	.datad(!Xd_0__inst_mult_22_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_56 ),
	.sharein(Xd_0__inst_mult_22_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_59 ),
	.cout(Xd_0__inst_mult_22_60 ),
	.shareout(Xd_0__inst_mult_22_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_23_20 (
// Equation(s):
// Xd_0__inst_mult_23_59  = SUM(( !Xd_0__inst_mult_23_8_q  $ (!Xd_0__inst_mult_23_9_q  $ (((Xd_0__inst_mult_23_4_q  & Xd_0__inst_mult_23_10_q )))) ) + ( Xd_0__inst_mult_23_57  ) + ( Xd_0__inst_mult_23_56  ))
// Xd_0__inst_mult_23_60  = CARRY(( !Xd_0__inst_mult_23_8_q  $ (!Xd_0__inst_mult_23_9_q  $ (((Xd_0__inst_mult_23_4_q  & Xd_0__inst_mult_23_10_q )))) ) + ( Xd_0__inst_mult_23_57  ) + ( Xd_0__inst_mult_23_56  ))
// Xd_0__inst_mult_23_61  = SHARE((!Xd_0__inst_mult_23_8_q  & (Xd_0__inst_mult_23_9_q  & (Xd_0__inst_mult_23_4_q  & Xd_0__inst_mult_23_10_q ))) # (Xd_0__inst_mult_23_8_q  & (((Xd_0__inst_mult_23_4_q  & Xd_0__inst_mult_23_10_q )) # (Xd_0__inst_mult_23_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_23_8_q ),
	.datab(!Xd_0__inst_mult_23_9_q ),
	.datac(!Xd_0__inst_mult_23_4_q ),
	.datad(!Xd_0__inst_mult_23_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_56 ),
	.sharein(Xd_0__inst_mult_23_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_59 ),
	.cout(Xd_0__inst_mult_23_60 ),
	.shareout(Xd_0__inst_mult_23_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_20_20 (
// Equation(s):
// Xd_0__inst_mult_20_59  = SUM(( !Xd_0__inst_mult_20_8_q  $ (!Xd_0__inst_mult_20_9_q  $ (((Xd_0__inst_mult_20_4_q  & Xd_0__inst_mult_20_10_q )))) ) + ( Xd_0__inst_mult_20_57  ) + ( Xd_0__inst_mult_20_56  ))
// Xd_0__inst_mult_20_60  = CARRY(( !Xd_0__inst_mult_20_8_q  $ (!Xd_0__inst_mult_20_9_q  $ (((Xd_0__inst_mult_20_4_q  & Xd_0__inst_mult_20_10_q )))) ) + ( Xd_0__inst_mult_20_57  ) + ( Xd_0__inst_mult_20_56  ))
// Xd_0__inst_mult_20_61  = SHARE((!Xd_0__inst_mult_20_8_q  & (Xd_0__inst_mult_20_9_q  & (Xd_0__inst_mult_20_4_q  & Xd_0__inst_mult_20_10_q ))) # (Xd_0__inst_mult_20_8_q  & (((Xd_0__inst_mult_20_4_q  & Xd_0__inst_mult_20_10_q )) # (Xd_0__inst_mult_20_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_20_8_q ),
	.datab(!Xd_0__inst_mult_20_9_q ),
	.datac(!Xd_0__inst_mult_20_4_q ),
	.datad(!Xd_0__inst_mult_20_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_56 ),
	.sharein(Xd_0__inst_mult_20_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_59 ),
	.cout(Xd_0__inst_mult_20_60 ),
	.shareout(Xd_0__inst_mult_20_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_21_16 (
// Equation(s):
// Xd_0__inst_mult_21_43  = SUM(( !Xd_0__inst_mult_21_8_q  $ (!Xd_0__inst_mult_21_9_q  $ (((Xd_0__inst_mult_21_4_q  & Xd_0__inst_mult_21_10_q )))) ) + ( Xd_0__inst_mult_21_42  ) + ( Xd_0__inst_mult_21_41  ))
// Xd_0__inst_mult_21_44  = CARRY(( !Xd_0__inst_mult_21_8_q  $ (!Xd_0__inst_mult_21_9_q  $ (((Xd_0__inst_mult_21_4_q  & Xd_0__inst_mult_21_10_q )))) ) + ( Xd_0__inst_mult_21_42  ) + ( Xd_0__inst_mult_21_41  ))
// Xd_0__inst_mult_21_45  = SHARE((!Xd_0__inst_mult_21_8_q  & (Xd_0__inst_mult_21_9_q  & (Xd_0__inst_mult_21_4_q  & Xd_0__inst_mult_21_10_q ))) # (Xd_0__inst_mult_21_8_q  & (((Xd_0__inst_mult_21_4_q  & Xd_0__inst_mult_21_10_q )) # (Xd_0__inst_mult_21_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_21_8_q ),
	.datab(!Xd_0__inst_mult_21_9_q ),
	.datac(!Xd_0__inst_mult_21_4_q ),
	.datad(!Xd_0__inst_mult_21_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_41 ),
	.sharein(Xd_0__inst_mult_21_42 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_43 ),
	.cout(Xd_0__inst_mult_21_44 ),
	.shareout(Xd_0__inst_mult_21_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_18_16 (
// Equation(s):
// Xd_0__inst_mult_18_42  = SUM(( !Xd_0__inst_mult_18_8_q  $ (!Xd_0__inst_mult_18_9_q  $ (((Xd_0__inst_mult_18_4_q  & Xd_0__inst_mult_18_10_q )))) ) + ( Xd_0__inst_mult_18_41  ) + ( Xd_0__inst_mult_18_40  ))
// Xd_0__inst_mult_18_43  = CARRY(( !Xd_0__inst_mult_18_8_q  $ (!Xd_0__inst_mult_18_9_q  $ (((Xd_0__inst_mult_18_4_q  & Xd_0__inst_mult_18_10_q )))) ) + ( Xd_0__inst_mult_18_41  ) + ( Xd_0__inst_mult_18_40  ))
// Xd_0__inst_mult_18_44  = SHARE((!Xd_0__inst_mult_18_8_q  & (Xd_0__inst_mult_18_9_q  & (Xd_0__inst_mult_18_4_q  & Xd_0__inst_mult_18_10_q ))) # (Xd_0__inst_mult_18_8_q  & (((Xd_0__inst_mult_18_4_q  & Xd_0__inst_mult_18_10_q )) # (Xd_0__inst_mult_18_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_18_8_q ),
	.datab(!Xd_0__inst_mult_18_9_q ),
	.datac(!Xd_0__inst_mult_18_4_q ),
	.datad(!Xd_0__inst_mult_18_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_40 ),
	.sharein(Xd_0__inst_mult_18_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_42 ),
	.cout(Xd_0__inst_mult_18_43 ),
	.shareout(Xd_0__inst_mult_18_44 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_19_19 (
// Equation(s):
// Xd_0__inst_mult_19_55  = SUM(( !Xd_0__inst_mult_19_8_q  $ (!Xd_0__inst_mult_19_9_q  $ (((Xd_0__inst_mult_19_4_q  & Xd_0__inst_mult_19_10_q )))) ) + ( Xd_0__inst_mult_19_53  ) + ( Xd_0__inst_mult_19_52  ))
// Xd_0__inst_mult_19_56  = CARRY(( !Xd_0__inst_mult_19_8_q  $ (!Xd_0__inst_mult_19_9_q  $ (((Xd_0__inst_mult_19_4_q  & Xd_0__inst_mult_19_10_q )))) ) + ( Xd_0__inst_mult_19_53  ) + ( Xd_0__inst_mult_19_52  ))
// Xd_0__inst_mult_19_57  = SHARE((!Xd_0__inst_mult_19_8_q  & (Xd_0__inst_mult_19_9_q  & (Xd_0__inst_mult_19_4_q  & Xd_0__inst_mult_19_10_q ))) # (Xd_0__inst_mult_19_8_q  & (((Xd_0__inst_mult_19_4_q  & Xd_0__inst_mult_19_10_q )) # (Xd_0__inst_mult_19_9_q 
// ))))

	.dataa(!Xd_0__inst_mult_19_8_q ),
	.datab(!Xd_0__inst_mult_19_9_q ),
	.datac(!Xd_0__inst_mult_19_4_q ),
	.datad(!Xd_0__inst_mult_19_10_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_52 ),
	.sharein(Xd_0__inst_mult_19_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_55 ),
	.cout(Xd_0__inst_mult_19_56 ),
	.shareout(Xd_0__inst_mult_19_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_16_17 (
// Equation(s):
// Xd_0__inst_mult_16_46  = SUM(( !Xd_0__inst_mult_16_12_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_11_q ))) ) + ( Xd_0__inst_mult_16_44  ) + ( Xd_0__inst_mult_16_43  ))
// Xd_0__inst_mult_16_47  = CARRY(( !Xd_0__inst_mult_16_12_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_11_q ))) ) + ( Xd_0__inst_mult_16_44  ) + ( Xd_0__inst_mult_16_43  ))
// Xd_0__inst_mult_16_48  = SHARE((Xd_0__inst_mult_16_4_q  & (Xd_0__inst_mult_16_11_q  & Xd_0__inst_mult_16_12_q )))

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_11_q ),
	.datac(!Xd_0__inst_mult_16_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_43 ),
	.sharein(Xd_0__inst_mult_16_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_46 ),
	.cout(Xd_0__inst_mult_16_47 ),
	.shareout(Xd_0__inst_mult_16_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_17_17 (
// Equation(s):
// Xd_0__inst_mult_17_47  = SUM(( !Xd_0__inst_mult_17_12_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_11_q ))) ) + ( Xd_0__inst_mult_17_45  ) + ( Xd_0__inst_mult_17_44  ))
// Xd_0__inst_mult_17_48  = CARRY(( !Xd_0__inst_mult_17_12_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_11_q ))) ) + ( Xd_0__inst_mult_17_45  ) + ( Xd_0__inst_mult_17_44  ))
// Xd_0__inst_mult_17_49  = SHARE((Xd_0__inst_mult_17_4_q  & (Xd_0__inst_mult_17_11_q  & Xd_0__inst_mult_17_12_q )))

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_11_q ),
	.datac(!Xd_0__inst_mult_17_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_44 ),
	.sharein(Xd_0__inst_mult_17_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_47 ),
	.cout(Xd_0__inst_mult_17_48 ),
	.shareout(Xd_0__inst_mult_17_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_17 (
// Equation(s):
// Xd_0__inst_mult_14_46  = SUM(( !Xd_0__inst_mult_14_12_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_11_q ))) ) + ( Xd_0__inst_mult_14_44  ) + ( Xd_0__inst_mult_14_43  ))
// Xd_0__inst_mult_14_47  = CARRY(( !Xd_0__inst_mult_14_12_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_11_q ))) ) + ( Xd_0__inst_mult_14_44  ) + ( Xd_0__inst_mult_14_43  ))
// Xd_0__inst_mult_14_48  = SHARE((Xd_0__inst_mult_14_4_q  & (Xd_0__inst_mult_14_11_q  & Xd_0__inst_mult_14_12_q )))

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_11_q ),
	.datac(!Xd_0__inst_mult_14_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_43 ),
	.sharein(Xd_0__inst_mult_14_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_46 ),
	.cout(Xd_0__inst_mult_14_47 ),
	.shareout(Xd_0__inst_mult_14_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_17 (
// Equation(s):
// Xd_0__inst_mult_15_47  = SUM(( !Xd_0__inst_mult_15_12_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_11_q ))) ) + ( Xd_0__inst_mult_15_45  ) + ( Xd_0__inst_mult_15_44  ))
// Xd_0__inst_mult_15_48  = CARRY(( !Xd_0__inst_mult_15_12_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_11_q ))) ) + ( Xd_0__inst_mult_15_45  ) + ( Xd_0__inst_mult_15_44  ))
// Xd_0__inst_mult_15_49  = SHARE((Xd_0__inst_mult_15_4_q  & (Xd_0__inst_mult_15_11_q  & Xd_0__inst_mult_15_12_q )))

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_11_q ),
	.datac(!Xd_0__inst_mult_15_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_44 ),
	.sharein(Xd_0__inst_mult_15_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_47 ),
	.cout(Xd_0__inst_mult_15_48 ),
	.shareout(Xd_0__inst_mult_15_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_17 (
// Equation(s):
// Xd_0__inst_mult_12_46  = SUM(( !Xd_0__inst_mult_12_12_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_11_q ))) ) + ( Xd_0__inst_mult_12_44  ) + ( Xd_0__inst_mult_12_43  ))
// Xd_0__inst_mult_12_47  = CARRY(( !Xd_0__inst_mult_12_12_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_11_q ))) ) + ( Xd_0__inst_mult_12_44  ) + ( Xd_0__inst_mult_12_43  ))
// Xd_0__inst_mult_12_48  = SHARE((Xd_0__inst_mult_12_4_q  & (Xd_0__inst_mult_12_11_q  & Xd_0__inst_mult_12_12_q )))

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_11_q ),
	.datac(!Xd_0__inst_mult_12_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_43 ),
	.sharein(Xd_0__inst_mult_12_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_46 ),
	.cout(Xd_0__inst_mult_12_47 ),
	.shareout(Xd_0__inst_mult_12_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_17 (
// Equation(s):
// Xd_0__inst_mult_13_47  = SUM(( !Xd_0__inst_mult_13_12_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_11_q ))) ) + ( Xd_0__inst_mult_13_45  ) + ( Xd_0__inst_mult_13_44  ))
// Xd_0__inst_mult_13_48  = CARRY(( !Xd_0__inst_mult_13_12_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_11_q ))) ) + ( Xd_0__inst_mult_13_45  ) + ( Xd_0__inst_mult_13_44  ))
// Xd_0__inst_mult_13_49  = SHARE((Xd_0__inst_mult_13_4_q  & (Xd_0__inst_mult_13_11_q  & Xd_0__inst_mult_13_12_q )))

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_11_q ),
	.datac(!Xd_0__inst_mult_13_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_44 ),
	.sharein(Xd_0__inst_mult_13_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_47 ),
	.cout(Xd_0__inst_mult_13_48 ),
	.shareout(Xd_0__inst_mult_13_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_17 (
// Equation(s):
// Xd_0__inst_mult_10_46  = SUM(( !Xd_0__inst_mult_10_12_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_11_q ))) ) + ( Xd_0__inst_mult_10_44  ) + ( Xd_0__inst_mult_10_43  ))
// Xd_0__inst_mult_10_47  = CARRY(( !Xd_0__inst_mult_10_12_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_11_q ))) ) + ( Xd_0__inst_mult_10_44  ) + ( Xd_0__inst_mult_10_43  ))
// Xd_0__inst_mult_10_48  = SHARE((Xd_0__inst_mult_10_4_q  & (Xd_0__inst_mult_10_11_q  & Xd_0__inst_mult_10_12_q )))

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_11_q ),
	.datac(!Xd_0__inst_mult_10_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_43 ),
	.sharein(Xd_0__inst_mult_10_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_46 ),
	.cout(Xd_0__inst_mult_10_47 ),
	.shareout(Xd_0__inst_mult_10_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_19 (
// Equation(s):
// Xd_0__inst_mult_11_55  = SUM(( !Xd_0__inst_mult_11_12_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_11_q ))) ) + ( Xd_0__inst_mult_11_53  ) + ( Xd_0__inst_mult_11_52  ))
// Xd_0__inst_mult_11_56  = CARRY(( !Xd_0__inst_mult_11_12_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_11_q ))) ) + ( Xd_0__inst_mult_11_53  ) + ( Xd_0__inst_mult_11_52  ))
// Xd_0__inst_mult_11_57  = SHARE((Xd_0__inst_mult_11_4_q  & (Xd_0__inst_mult_11_11_q  & Xd_0__inst_mult_11_12_q )))

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_11_q ),
	.datac(!Xd_0__inst_mult_11_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_52 ),
	.sharein(Xd_0__inst_mult_11_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_55 ),
	.cout(Xd_0__inst_mult_11_56 ),
	.shareout(Xd_0__inst_mult_11_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_17 (
// Equation(s):
// Xd_0__inst_mult_8_46  = SUM(( !Xd_0__inst_mult_8_12_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_11_q ))) ) + ( Xd_0__inst_mult_8_44  ) + ( Xd_0__inst_mult_8_43  ))
// Xd_0__inst_mult_8_47  = CARRY(( !Xd_0__inst_mult_8_12_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_11_q ))) ) + ( Xd_0__inst_mult_8_44  ) + ( Xd_0__inst_mult_8_43  ))
// Xd_0__inst_mult_8_48  = SHARE((Xd_0__inst_mult_8_4_q  & (Xd_0__inst_mult_8_11_q  & Xd_0__inst_mult_8_12_q )))

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_11_q ),
	.datac(!Xd_0__inst_mult_8_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_43 ),
	.sharein(Xd_0__inst_mult_8_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_46 ),
	.cout(Xd_0__inst_mult_8_47 ),
	.shareout(Xd_0__inst_mult_8_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_17 (
// Equation(s):
// Xd_0__inst_mult_9_47  = SUM(( !Xd_0__inst_mult_9_12_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_11_q ))) ) + ( Xd_0__inst_mult_9_45  ) + ( Xd_0__inst_mult_9_44  ))
// Xd_0__inst_mult_9_48  = CARRY(( !Xd_0__inst_mult_9_12_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_11_q ))) ) + ( Xd_0__inst_mult_9_45  ) + ( Xd_0__inst_mult_9_44  ))
// Xd_0__inst_mult_9_49  = SHARE((Xd_0__inst_mult_9_4_q  & (Xd_0__inst_mult_9_11_q  & Xd_0__inst_mult_9_12_q )))

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_11_q ),
	.datac(!Xd_0__inst_mult_9_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_44 ),
	.sharein(Xd_0__inst_mult_9_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_47 ),
	.cout(Xd_0__inst_mult_9_48 ),
	.shareout(Xd_0__inst_mult_9_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_17 (
// Equation(s):
// Xd_0__inst_mult_6_45  = SUM(( !Xd_0__inst_mult_6_12_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_11_q ))) ) + ( Xd_0__inst_mult_6_43  ) + ( Xd_0__inst_mult_6_42  ))
// Xd_0__inst_mult_6_46  = CARRY(( !Xd_0__inst_mult_6_12_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_11_q ))) ) + ( Xd_0__inst_mult_6_43  ) + ( Xd_0__inst_mult_6_42  ))
// Xd_0__inst_mult_6_47  = SHARE((Xd_0__inst_mult_6_4_q  & (Xd_0__inst_mult_6_11_q  & Xd_0__inst_mult_6_12_q )))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(!Xd_0__inst_mult_6_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_42 ),
	.sharein(Xd_0__inst_mult_6_43 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_45 ),
	.cout(Xd_0__inst_mult_6_46 ),
	.shareout(Xd_0__inst_mult_6_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_17 (
// Equation(s):
// Xd_0__inst_mult_7_46  = SUM(( !Xd_0__inst_mult_7_12_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_11_q ))) ) + ( Xd_0__inst_mult_7_44  ) + ( Xd_0__inst_mult_7_43  ))
// Xd_0__inst_mult_7_47  = CARRY(( !Xd_0__inst_mult_7_12_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_11_q ))) ) + ( Xd_0__inst_mult_7_44  ) + ( Xd_0__inst_mult_7_43  ))
// Xd_0__inst_mult_7_48  = SHARE((Xd_0__inst_mult_7_4_q  & (Xd_0__inst_mult_7_11_q  & Xd_0__inst_mult_7_12_q )))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(!Xd_0__inst_mult_7_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_43 ),
	.sharein(Xd_0__inst_mult_7_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_46 ),
	.cout(Xd_0__inst_mult_7_47 ),
	.shareout(Xd_0__inst_mult_7_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_17 (
// Equation(s):
// Xd_0__inst_mult_4_45  = SUM(( !Xd_0__inst_mult_4_12_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_11_q ))) ) + ( Xd_0__inst_mult_4_43  ) + ( Xd_0__inst_mult_4_42  ))
// Xd_0__inst_mult_4_46  = CARRY(( !Xd_0__inst_mult_4_12_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_11_q ))) ) + ( Xd_0__inst_mult_4_43  ) + ( Xd_0__inst_mult_4_42  ))
// Xd_0__inst_mult_4_47  = SHARE((Xd_0__inst_mult_4_4_q  & (Xd_0__inst_mult_4_11_q  & Xd_0__inst_mult_4_12_q )))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(!Xd_0__inst_mult_4_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_42 ),
	.sharein(Xd_0__inst_mult_4_43 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_45 ),
	.cout(Xd_0__inst_mult_4_46 ),
	.shareout(Xd_0__inst_mult_4_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_17 (
// Equation(s):
// Xd_0__inst_mult_5_46  = SUM(( !Xd_0__inst_mult_5_12_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_11_q ))) ) + ( Xd_0__inst_mult_5_44  ) + ( Xd_0__inst_mult_5_43  ))
// Xd_0__inst_mult_5_47  = CARRY(( !Xd_0__inst_mult_5_12_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_11_q ))) ) + ( Xd_0__inst_mult_5_44  ) + ( Xd_0__inst_mult_5_43  ))
// Xd_0__inst_mult_5_48  = SHARE((Xd_0__inst_mult_5_4_q  & (Xd_0__inst_mult_5_11_q  & Xd_0__inst_mult_5_12_q )))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(!Xd_0__inst_mult_5_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_43 ),
	.sharein(Xd_0__inst_mult_5_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_46 ),
	.cout(Xd_0__inst_mult_5_47 ),
	.shareout(Xd_0__inst_mult_5_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_18 (
// Equation(s):
// Xd_0__inst_mult_2_50  = SUM(( !Xd_0__inst_mult_2_12_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_11_q ))) ) + ( Xd_0__inst_mult_2_48  ) + ( Xd_0__inst_mult_2_47  ))
// Xd_0__inst_mult_2_51  = CARRY(( !Xd_0__inst_mult_2_12_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_11_q ))) ) + ( Xd_0__inst_mult_2_48  ) + ( Xd_0__inst_mult_2_47  ))
// Xd_0__inst_mult_2_52  = SHARE((Xd_0__inst_mult_2_4_q  & (Xd_0__inst_mult_2_11_q  & Xd_0__inst_mult_2_12_q )))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(!Xd_0__inst_mult_2_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_47 ),
	.sharein(Xd_0__inst_mult_2_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_50 ),
	.cout(Xd_0__inst_mult_2_51 ),
	.shareout(Xd_0__inst_mult_2_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_18 (
// Equation(s):
// Xd_0__inst_mult_3_50  = SUM(( !Xd_0__inst_mult_3_12_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_11_q ))) ) + ( Xd_0__inst_mult_3_48  ) + ( Xd_0__inst_mult_3_47  ))
// Xd_0__inst_mult_3_51  = CARRY(( !Xd_0__inst_mult_3_12_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_11_q ))) ) + ( Xd_0__inst_mult_3_48  ) + ( Xd_0__inst_mult_3_47  ))
// Xd_0__inst_mult_3_52  = SHARE((Xd_0__inst_mult_3_4_q  & (Xd_0__inst_mult_3_11_q  & Xd_0__inst_mult_3_12_q )))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(!Xd_0__inst_mult_3_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_47 ),
	.sharein(Xd_0__inst_mult_3_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_50 ),
	.cout(Xd_0__inst_mult_3_51 ),
	.shareout(Xd_0__inst_mult_3_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_18 (
// Equation(s):
// Xd_0__inst_mult_0_50  = SUM(( !Xd_0__inst_mult_0_12_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_11_q ))) ) + ( Xd_0__inst_mult_0_48  ) + ( Xd_0__inst_mult_0_47  ))
// Xd_0__inst_mult_0_51  = CARRY(( !Xd_0__inst_mult_0_12_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_11_q ))) ) + ( Xd_0__inst_mult_0_48  ) + ( Xd_0__inst_mult_0_47  ))
// Xd_0__inst_mult_0_52  = SHARE((Xd_0__inst_mult_0_4_q  & (Xd_0__inst_mult_0_11_q  & Xd_0__inst_mult_0_12_q )))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(!Xd_0__inst_mult_0_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_47 ),
	.sharein(Xd_0__inst_mult_0_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_50 ),
	.cout(Xd_0__inst_mult_0_51 ),
	.shareout(Xd_0__inst_mult_0_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_18 (
// Equation(s):
// Xd_0__inst_mult_1_50  = SUM(( !Xd_0__inst_mult_1_12_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_11_q ))) ) + ( Xd_0__inst_mult_1_48  ) + ( Xd_0__inst_mult_1_47  ))
// Xd_0__inst_mult_1_51  = CARRY(( !Xd_0__inst_mult_1_12_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_11_q ))) ) + ( Xd_0__inst_mult_1_48  ) + ( Xd_0__inst_mult_1_47  ))
// Xd_0__inst_mult_1_52  = SHARE((Xd_0__inst_mult_1_4_q  & (Xd_0__inst_mult_1_11_q  & Xd_0__inst_mult_1_12_q )))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(!Xd_0__inst_mult_1_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_47 ),
	.sharein(Xd_0__inst_mult_1_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_50 ),
	.cout(Xd_0__inst_mult_1_51 ),
	.shareout(Xd_0__inst_mult_1_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_28_21 (
// Equation(s):
// Xd_0__inst_mult_28_63  = SUM(( !Xd_0__inst_mult_28_12_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_11_q ))) ) + ( Xd_0__inst_mult_28_61  ) + ( Xd_0__inst_mult_28_60  ))
// Xd_0__inst_mult_28_64  = CARRY(( !Xd_0__inst_mult_28_12_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_11_q ))) ) + ( Xd_0__inst_mult_28_61  ) + ( Xd_0__inst_mult_28_60  ))
// Xd_0__inst_mult_28_65  = SHARE((Xd_0__inst_mult_28_4_q  & (Xd_0__inst_mult_28_11_q  & Xd_0__inst_mult_28_12_q )))

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_11_q ),
	.datac(!Xd_0__inst_mult_28_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_60 ),
	.sharein(Xd_0__inst_mult_28_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_63 ),
	.cout(Xd_0__inst_mult_28_64 ),
	.shareout(Xd_0__inst_mult_28_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_29_19 (
// Equation(s):
// Xd_0__inst_mult_29_55  = SUM(( !Xd_0__inst_mult_29_12_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_11_q ))) ) + ( Xd_0__inst_mult_29_53  ) + ( Xd_0__inst_mult_29_52  ))
// Xd_0__inst_mult_29_56  = CARRY(( !Xd_0__inst_mult_29_12_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_11_q ))) ) + ( Xd_0__inst_mult_29_53  ) + ( Xd_0__inst_mult_29_52  ))
// Xd_0__inst_mult_29_57  = SHARE((Xd_0__inst_mult_29_4_q  & (Xd_0__inst_mult_29_11_q  & Xd_0__inst_mult_29_12_q )))

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_11_q ),
	.datac(!Xd_0__inst_mult_29_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_52 ),
	.sharein(Xd_0__inst_mult_29_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_55 ),
	.cout(Xd_0__inst_mult_29_56 ),
	.shareout(Xd_0__inst_mult_29_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_26_21 (
// Equation(s):
// Xd_0__inst_mult_26_63  = SUM(( !Xd_0__inst_mult_26_12_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_11_q ))) ) + ( Xd_0__inst_mult_26_61  ) + ( Xd_0__inst_mult_26_60  ))
// Xd_0__inst_mult_26_64  = CARRY(( !Xd_0__inst_mult_26_12_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_11_q ))) ) + ( Xd_0__inst_mult_26_61  ) + ( Xd_0__inst_mult_26_60  ))
// Xd_0__inst_mult_26_65  = SHARE((Xd_0__inst_mult_26_4_q  & (Xd_0__inst_mult_26_11_q  & Xd_0__inst_mult_26_12_q )))

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_11_q ),
	.datac(!Xd_0__inst_mult_26_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_60 ),
	.sharein(Xd_0__inst_mult_26_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_63 ),
	.cout(Xd_0__inst_mult_26_64 ),
	.shareout(Xd_0__inst_mult_26_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_27_19 (
// Equation(s):
// Xd_0__inst_mult_27_55  = SUM(( !Xd_0__inst_mult_27_12_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_11_q ))) ) + ( Xd_0__inst_mult_27_53  ) + ( Xd_0__inst_mult_27_52  ))
// Xd_0__inst_mult_27_56  = CARRY(( !Xd_0__inst_mult_27_12_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_11_q ))) ) + ( Xd_0__inst_mult_27_53  ) + ( Xd_0__inst_mult_27_52  ))
// Xd_0__inst_mult_27_57  = SHARE((Xd_0__inst_mult_27_4_q  & (Xd_0__inst_mult_27_11_q  & Xd_0__inst_mult_27_12_q )))

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_11_q ),
	.datac(!Xd_0__inst_mult_27_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_52 ),
	.sharein(Xd_0__inst_mult_27_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_55 ),
	.cout(Xd_0__inst_mult_27_56 ),
	.shareout(Xd_0__inst_mult_27_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_24_21 (
// Equation(s):
// Xd_0__inst_mult_24_63  = SUM(( !Xd_0__inst_mult_24_12_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_11_q ))) ) + ( Xd_0__inst_mult_24_61  ) + ( Xd_0__inst_mult_24_60  ))
// Xd_0__inst_mult_24_64  = CARRY(( !Xd_0__inst_mult_24_12_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_11_q ))) ) + ( Xd_0__inst_mult_24_61  ) + ( Xd_0__inst_mult_24_60  ))
// Xd_0__inst_mult_24_65  = SHARE((Xd_0__inst_mult_24_4_q  & (Xd_0__inst_mult_24_11_q  & Xd_0__inst_mult_24_12_q )))

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_11_q ),
	.datac(!Xd_0__inst_mult_24_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_60 ),
	.sharein(Xd_0__inst_mult_24_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_63 ),
	.cout(Xd_0__inst_mult_24_64 ),
	.shareout(Xd_0__inst_mult_24_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_25_19 (
// Equation(s):
// Xd_0__inst_mult_25_55  = SUM(( !Xd_0__inst_mult_25_12_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_11_q ))) ) + ( Xd_0__inst_mult_25_53  ) + ( Xd_0__inst_mult_25_52  ))
// Xd_0__inst_mult_25_56  = CARRY(( !Xd_0__inst_mult_25_12_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_11_q ))) ) + ( Xd_0__inst_mult_25_53  ) + ( Xd_0__inst_mult_25_52  ))
// Xd_0__inst_mult_25_57  = SHARE((Xd_0__inst_mult_25_4_q  & (Xd_0__inst_mult_25_11_q  & Xd_0__inst_mult_25_12_q )))

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_11_q ),
	.datac(!Xd_0__inst_mult_25_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_52 ),
	.sharein(Xd_0__inst_mult_25_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_55 ),
	.cout(Xd_0__inst_mult_25_56 ),
	.shareout(Xd_0__inst_mult_25_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_22_21 (
// Equation(s):
// Xd_0__inst_mult_22_63  = SUM(( !Xd_0__inst_mult_22_12_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_11_q ))) ) + ( Xd_0__inst_mult_22_61  ) + ( Xd_0__inst_mult_22_60  ))
// Xd_0__inst_mult_22_64  = CARRY(( !Xd_0__inst_mult_22_12_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_11_q ))) ) + ( Xd_0__inst_mult_22_61  ) + ( Xd_0__inst_mult_22_60  ))
// Xd_0__inst_mult_22_65  = SHARE((Xd_0__inst_mult_22_4_q  & (Xd_0__inst_mult_22_11_q  & Xd_0__inst_mult_22_12_q )))

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_11_q ),
	.datac(!Xd_0__inst_mult_22_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_60 ),
	.sharein(Xd_0__inst_mult_22_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_63 ),
	.cout(Xd_0__inst_mult_22_64 ),
	.shareout(Xd_0__inst_mult_22_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_23_21 (
// Equation(s):
// Xd_0__inst_mult_23_63  = SUM(( !Xd_0__inst_mult_23_12_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_11_q ))) ) + ( Xd_0__inst_mult_23_61  ) + ( Xd_0__inst_mult_23_60  ))
// Xd_0__inst_mult_23_64  = CARRY(( !Xd_0__inst_mult_23_12_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_11_q ))) ) + ( Xd_0__inst_mult_23_61  ) + ( Xd_0__inst_mult_23_60  ))
// Xd_0__inst_mult_23_65  = SHARE((Xd_0__inst_mult_23_4_q  & (Xd_0__inst_mult_23_11_q  & Xd_0__inst_mult_23_12_q )))

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_11_q ),
	.datac(!Xd_0__inst_mult_23_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_60 ),
	.sharein(Xd_0__inst_mult_23_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_63 ),
	.cout(Xd_0__inst_mult_23_64 ),
	.shareout(Xd_0__inst_mult_23_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_20_21 (
// Equation(s):
// Xd_0__inst_mult_20_63  = SUM(( !Xd_0__inst_mult_20_12_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_11_q ))) ) + ( Xd_0__inst_mult_20_61  ) + ( Xd_0__inst_mult_20_60  ))
// Xd_0__inst_mult_20_64  = CARRY(( !Xd_0__inst_mult_20_12_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_11_q ))) ) + ( Xd_0__inst_mult_20_61  ) + ( Xd_0__inst_mult_20_60  ))
// Xd_0__inst_mult_20_65  = SHARE((Xd_0__inst_mult_20_4_q  & (Xd_0__inst_mult_20_11_q  & Xd_0__inst_mult_20_12_q )))

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_11_q ),
	.datac(!Xd_0__inst_mult_20_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_60 ),
	.sharein(Xd_0__inst_mult_20_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_63 ),
	.cout(Xd_0__inst_mult_20_64 ),
	.shareout(Xd_0__inst_mult_20_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_21_17 (
// Equation(s):
// Xd_0__inst_mult_21_47  = SUM(( !Xd_0__inst_mult_21_12_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_11_q ))) ) + ( Xd_0__inst_mult_21_45  ) + ( Xd_0__inst_mult_21_44  ))
// Xd_0__inst_mult_21_48  = CARRY(( !Xd_0__inst_mult_21_12_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_11_q ))) ) + ( Xd_0__inst_mult_21_45  ) + ( Xd_0__inst_mult_21_44  ))
// Xd_0__inst_mult_21_49  = SHARE((Xd_0__inst_mult_21_4_q  & (Xd_0__inst_mult_21_11_q  & Xd_0__inst_mult_21_12_q )))

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_11_q ),
	.datac(!Xd_0__inst_mult_21_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_44 ),
	.sharein(Xd_0__inst_mult_21_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_47 ),
	.cout(Xd_0__inst_mult_21_48 ),
	.shareout(Xd_0__inst_mult_21_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_18_17 (
// Equation(s):
// Xd_0__inst_mult_18_46  = SUM(( !Xd_0__inst_mult_18_12_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_11_q ))) ) + ( Xd_0__inst_mult_18_44  ) + ( Xd_0__inst_mult_18_43  ))
// Xd_0__inst_mult_18_47  = CARRY(( !Xd_0__inst_mult_18_12_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_11_q ))) ) + ( Xd_0__inst_mult_18_44  ) + ( Xd_0__inst_mult_18_43  ))
// Xd_0__inst_mult_18_48  = SHARE((Xd_0__inst_mult_18_4_q  & (Xd_0__inst_mult_18_11_q  & Xd_0__inst_mult_18_12_q )))

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_11_q ),
	.datac(!Xd_0__inst_mult_18_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_43 ),
	.sharein(Xd_0__inst_mult_18_44 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_46 ),
	.cout(Xd_0__inst_mult_18_47 ),
	.shareout(Xd_0__inst_mult_18_48 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_19_20 (
// Equation(s):
// Xd_0__inst_mult_19_59  = SUM(( !Xd_0__inst_mult_19_12_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_11_q ))) ) + ( Xd_0__inst_mult_19_57  ) + ( Xd_0__inst_mult_19_56  ))
// Xd_0__inst_mult_19_60  = CARRY(( !Xd_0__inst_mult_19_12_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_11_q ))) ) + ( Xd_0__inst_mult_19_57  ) + ( Xd_0__inst_mult_19_56  ))
// Xd_0__inst_mult_19_61  = SHARE((Xd_0__inst_mult_19_4_q  & (Xd_0__inst_mult_19_11_q  & Xd_0__inst_mult_19_12_q )))

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_11_q ),
	.datac(!Xd_0__inst_mult_19_12_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_56 ),
	.sharein(Xd_0__inst_mult_19_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_59 ),
	.cout(Xd_0__inst_mult_19_60 ),
	.shareout(Xd_0__inst_mult_19_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_16_18 (
// Equation(s):
// Xd_0__inst_mult_16_50  = SUM(( !Xd_0__inst_mult_16_13_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_0_q ))) ) + ( Xd_0__inst_mult_16_48  ) + ( Xd_0__inst_mult_16_47  ))
// Xd_0__inst_mult_16_51  = CARRY(( !Xd_0__inst_mult_16_13_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_0_q ))) ) + ( Xd_0__inst_mult_16_48  ) + ( Xd_0__inst_mult_16_47  ))
// Xd_0__inst_mult_16_52  = SHARE((Xd_0__inst_mult_16_4_q  & (Xd_0__inst_mult_16_0_q  & Xd_0__inst_mult_16_13_q )))

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_0_q ),
	.datac(!Xd_0__inst_mult_16_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_47 ),
	.sharein(Xd_0__inst_mult_16_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_50 ),
	.cout(Xd_0__inst_mult_16_51 ),
	.shareout(Xd_0__inst_mult_16_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_17_18 (
// Equation(s):
// Xd_0__inst_mult_17_51  = SUM(( !Xd_0__inst_mult_17_13_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_0_q ))) ) + ( Xd_0__inst_mult_17_49  ) + ( Xd_0__inst_mult_17_48  ))
// Xd_0__inst_mult_17_52  = CARRY(( !Xd_0__inst_mult_17_13_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_0_q ))) ) + ( Xd_0__inst_mult_17_49  ) + ( Xd_0__inst_mult_17_48  ))
// Xd_0__inst_mult_17_53  = SHARE((Xd_0__inst_mult_17_4_q  & (Xd_0__inst_mult_17_0_q  & Xd_0__inst_mult_17_13_q )))

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_0_q ),
	.datac(!Xd_0__inst_mult_17_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_48 ),
	.sharein(Xd_0__inst_mult_17_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_51 ),
	.cout(Xd_0__inst_mult_17_52 ),
	.shareout(Xd_0__inst_mult_17_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_18 (
// Equation(s):
// Xd_0__inst_mult_14_50  = SUM(( !Xd_0__inst_mult_14_13_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_0_q ))) ) + ( Xd_0__inst_mult_14_48  ) + ( Xd_0__inst_mult_14_47  ))
// Xd_0__inst_mult_14_51  = CARRY(( !Xd_0__inst_mult_14_13_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_0_q ))) ) + ( Xd_0__inst_mult_14_48  ) + ( Xd_0__inst_mult_14_47  ))
// Xd_0__inst_mult_14_52  = SHARE((Xd_0__inst_mult_14_4_q  & (Xd_0__inst_mult_14_0_q  & Xd_0__inst_mult_14_13_q )))

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_0_q ),
	.datac(!Xd_0__inst_mult_14_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_47 ),
	.sharein(Xd_0__inst_mult_14_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_50 ),
	.cout(Xd_0__inst_mult_14_51 ),
	.shareout(Xd_0__inst_mult_14_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_18 (
// Equation(s):
// Xd_0__inst_mult_15_51  = SUM(( !Xd_0__inst_mult_15_13_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_0_q ))) ) + ( Xd_0__inst_mult_15_49  ) + ( Xd_0__inst_mult_15_48  ))
// Xd_0__inst_mult_15_52  = CARRY(( !Xd_0__inst_mult_15_13_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_0_q ))) ) + ( Xd_0__inst_mult_15_49  ) + ( Xd_0__inst_mult_15_48  ))
// Xd_0__inst_mult_15_53  = SHARE((Xd_0__inst_mult_15_4_q  & (Xd_0__inst_mult_15_0_q  & Xd_0__inst_mult_15_13_q )))

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_0_q ),
	.datac(!Xd_0__inst_mult_15_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_48 ),
	.sharein(Xd_0__inst_mult_15_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_51 ),
	.cout(Xd_0__inst_mult_15_52 ),
	.shareout(Xd_0__inst_mult_15_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_18 (
// Equation(s):
// Xd_0__inst_mult_12_50  = SUM(( !Xd_0__inst_mult_12_13_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_0_q ))) ) + ( Xd_0__inst_mult_12_48  ) + ( Xd_0__inst_mult_12_47  ))
// Xd_0__inst_mult_12_51  = CARRY(( !Xd_0__inst_mult_12_13_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_0_q ))) ) + ( Xd_0__inst_mult_12_48  ) + ( Xd_0__inst_mult_12_47  ))
// Xd_0__inst_mult_12_52  = SHARE((Xd_0__inst_mult_12_4_q  & (Xd_0__inst_mult_12_0_q  & Xd_0__inst_mult_12_13_q )))

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_0_q ),
	.datac(!Xd_0__inst_mult_12_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_47 ),
	.sharein(Xd_0__inst_mult_12_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_50 ),
	.cout(Xd_0__inst_mult_12_51 ),
	.shareout(Xd_0__inst_mult_12_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_18 (
// Equation(s):
// Xd_0__inst_mult_13_51  = SUM(( !Xd_0__inst_mult_13_13_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_0_q ))) ) + ( Xd_0__inst_mult_13_49  ) + ( Xd_0__inst_mult_13_48  ))
// Xd_0__inst_mult_13_52  = CARRY(( !Xd_0__inst_mult_13_13_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_0_q ))) ) + ( Xd_0__inst_mult_13_49  ) + ( Xd_0__inst_mult_13_48  ))
// Xd_0__inst_mult_13_53  = SHARE((Xd_0__inst_mult_13_4_q  & (Xd_0__inst_mult_13_0_q  & Xd_0__inst_mult_13_13_q )))

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_0_q ),
	.datac(!Xd_0__inst_mult_13_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_48 ),
	.sharein(Xd_0__inst_mult_13_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_51 ),
	.cout(Xd_0__inst_mult_13_52 ),
	.shareout(Xd_0__inst_mult_13_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_18 (
// Equation(s):
// Xd_0__inst_mult_10_50  = SUM(( !Xd_0__inst_mult_10_13_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_0_q ))) ) + ( Xd_0__inst_mult_10_48  ) + ( Xd_0__inst_mult_10_47  ))
// Xd_0__inst_mult_10_51  = CARRY(( !Xd_0__inst_mult_10_13_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_0_q ))) ) + ( Xd_0__inst_mult_10_48  ) + ( Xd_0__inst_mult_10_47  ))
// Xd_0__inst_mult_10_52  = SHARE((Xd_0__inst_mult_10_4_q  & (Xd_0__inst_mult_10_0_q  & Xd_0__inst_mult_10_13_q )))

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_0_q ),
	.datac(!Xd_0__inst_mult_10_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_47 ),
	.sharein(Xd_0__inst_mult_10_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_50 ),
	.cout(Xd_0__inst_mult_10_51 ),
	.shareout(Xd_0__inst_mult_10_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_20 (
// Equation(s):
// Xd_0__inst_mult_11_59  = SUM(( !Xd_0__inst_mult_11_13_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_0_q ))) ) + ( Xd_0__inst_mult_11_57  ) + ( Xd_0__inst_mult_11_56  ))
// Xd_0__inst_mult_11_60  = CARRY(( !Xd_0__inst_mult_11_13_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_0_q ))) ) + ( Xd_0__inst_mult_11_57  ) + ( Xd_0__inst_mult_11_56  ))
// Xd_0__inst_mult_11_61  = SHARE((Xd_0__inst_mult_11_4_q  & (Xd_0__inst_mult_11_0_q  & Xd_0__inst_mult_11_13_q )))

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_0_q ),
	.datac(!Xd_0__inst_mult_11_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_56 ),
	.sharein(Xd_0__inst_mult_11_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_59 ),
	.cout(Xd_0__inst_mult_11_60 ),
	.shareout(Xd_0__inst_mult_11_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_18 (
// Equation(s):
// Xd_0__inst_mult_8_50  = SUM(( !Xd_0__inst_mult_8_13_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_0_q ))) ) + ( Xd_0__inst_mult_8_48  ) + ( Xd_0__inst_mult_8_47  ))
// Xd_0__inst_mult_8_51  = CARRY(( !Xd_0__inst_mult_8_13_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_0_q ))) ) + ( Xd_0__inst_mult_8_48  ) + ( Xd_0__inst_mult_8_47  ))
// Xd_0__inst_mult_8_52  = SHARE((Xd_0__inst_mult_8_4_q  & (Xd_0__inst_mult_8_0_q  & Xd_0__inst_mult_8_13_q )))

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_0_q ),
	.datac(!Xd_0__inst_mult_8_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_47 ),
	.sharein(Xd_0__inst_mult_8_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_50 ),
	.cout(Xd_0__inst_mult_8_51 ),
	.shareout(Xd_0__inst_mult_8_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_18 (
// Equation(s):
// Xd_0__inst_mult_9_51  = SUM(( !Xd_0__inst_mult_9_13_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_0_q ))) ) + ( Xd_0__inst_mult_9_49  ) + ( Xd_0__inst_mult_9_48  ))
// Xd_0__inst_mult_9_52  = CARRY(( !Xd_0__inst_mult_9_13_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_0_q ))) ) + ( Xd_0__inst_mult_9_49  ) + ( Xd_0__inst_mult_9_48  ))
// Xd_0__inst_mult_9_53  = SHARE((Xd_0__inst_mult_9_4_q  & (Xd_0__inst_mult_9_0_q  & Xd_0__inst_mult_9_13_q )))

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_0_q ),
	.datac(!Xd_0__inst_mult_9_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_48 ),
	.sharein(Xd_0__inst_mult_9_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_51 ),
	.cout(Xd_0__inst_mult_9_52 ),
	.shareout(Xd_0__inst_mult_9_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_18 (
// Equation(s):
// Xd_0__inst_mult_6_49  = SUM(( !Xd_0__inst_mult_6_13_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_0_q ))) ) + ( Xd_0__inst_mult_6_47  ) + ( Xd_0__inst_mult_6_46  ))
// Xd_0__inst_mult_6_50  = CARRY(( !Xd_0__inst_mult_6_13_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_0_q ))) ) + ( Xd_0__inst_mult_6_47  ) + ( Xd_0__inst_mult_6_46  ))
// Xd_0__inst_mult_6_51  = SHARE((Xd_0__inst_mult_6_4_q  & (Xd_0__inst_mult_6_0_q  & Xd_0__inst_mult_6_13_q )))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_0_q ),
	.datac(!Xd_0__inst_mult_6_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_46 ),
	.sharein(Xd_0__inst_mult_6_47 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_49 ),
	.cout(Xd_0__inst_mult_6_50 ),
	.shareout(Xd_0__inst_mult_6_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_18 (
// Equation(s):
// Xd_0__inst_mult_7_50  = SUM(( !Xd_0__inst_mult_7_13_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_0_q ))) ) + ( Xd_0__inst_mult_7_48  ) + ( Xd_0__inst_mult_7_47  ))
// Xd_0__inst_mult_7_51  = CARRY(( !Xd_0__inst_mult_7_13_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_0_q ))) ) + ( Xd_0__inst_mult_7_48  ) + ( Xd_0__inst_mult_7_47  ))
// Xd_0__inst_mult_7_52  = SHARE((Xd_0__inst_mult_7_4_q  & (Xd_0__inst_mult_7_0_q  & Xd_0__inst_mult_7_13_q )))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_0_q ),
	.datac(!Xd_0__inst_mult_7_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_47 ),
	.sharein(Xd_0__inst_mult_7_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_50 ),
	.cout(Xd_0__inst_mult_7_51 ),
	.shareout(Xd_0__inst_mult_7_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_18 (
// Equation(s):
// Xd_0__inst_mult_4_49  = SUM(( !Xd_0__inst_mult_4_13_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_0_q ))) ) + ( Xd_0__inst_mult_4_47  ) + ( Xd_0__inst_mult_4_46  ))
// Xd_0__inst_mult_4_50  = CARRY(( !Xd_0__inst_mult_4_13_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_0_q ))) ) + ( Xd_0__inst_mult_4_47  ) + ( Xd_0__inst_mult_4_46  ))
// Xd_0__inst_mult_4_51  = SHARE((Xd_0__inst_mult_4_4_q  & (Xd_0__inst_mult_4_0_q  & Xd_0__inst_mult_4_13_q )))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_0_q ),
	.datac(!Xd_0__inst_mult_4_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_46 ),
	.sharein(Xd_0__inst_mult_4_47 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_49 ),
	.cout(Xd_0__inst_mult_4_50 ),
	.shareout(Xd_0__inst_mult_4_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_18 (
// Equation(s):
// Xd_0__inst_mult_5_50  = SUM(( !Xd_0__inst_mult_5_13_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_0_q ))) ) + ( Xd_0__inst_mult_5_48  ) + ( Xd_0__inst_mult_5_47  ))
// Xd_0__inst_mult_5_51  = CARRY(( !Xd_0__inst_mult_5_13_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_0_q ))) ) + ( Xd_0__inst_mult_5_48  ) + ( Xd_0__inst_mult_5_47  ))
// Xd_0__inst_mult_5_52  = SHARE((Xd_0__inst_mult_5_4_q  & (Xd_0__inst_mult_5_0_q  & Xd_0__inst_mult_5_13_q )))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_0_q ),
	.datac(!Xd_0__inst_mult_5_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_47 ),
	.sharein(Xd_0__inst_mult_5_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_50 ),
	.cout(Xd_0__inst_mult_5_51 ),
	.shareout(Xd_0__inst_mult_5_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_19 (
// Equation(s):
// Xd_0__inst_mult_2_54  = SUM(( !Xd_0__inst_mult_2_13_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_0_q ))) ) + ( Xd_0__inst_mult_2_52  ) + ( Xd_0__inst_mult_2_51  ))
// Xd_0__inst_mult_2_55  = CARRY(( !Xd_0__inst_mult_2_13_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_0_q ))) ) + ( Xd_0__inst_mult_2_52  ) + ( Xd_0__inst_mult_2_51  ))
// Xd_0__inst_mult_2_56  = SHARE((Xd_0__inst_mult_2_4_q  & (Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_13_q )))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_0_q ),
	.datac(!Xd_0__inst_mult_2_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_51 ),
	.sharein(Xd_0__inst_mult_2_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_54 ),
	.cout(Xd_0__inst_mult_2_55 ),
	.shareout(Xd_0__inst_mult_2_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_19 (
// Equation(s):
// Xd_0__inst_mult_3_54  = SUM(( !Xd_0__inst_mult_3_13_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_0_q ))) ) + ( Xd_0__inst_mult_3_52  ) + ( Xd_0__inst_mult_3_51  ))
// Xd_0__inst_mult_3_55  = CARRY(( !Xd_0__inst_mult_3_13_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_0_q ))) ) + ( Xd_0__inst_mult_3_52  ) + ( Xd_0__inst_mult_3_51  ))
// Xd_0__inst_mult_3_56  = SHARE((Xd_0__inst_mult_3_4_q  & (Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_13_q )))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_0_q ),
	.datac(!Xd_0__inst_mult_3_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_51 ),
	.sharein(Xd_0__inst_mult_3_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_54 ),
	.cout(Xd_0__inst_mult_3_55 ),
	.shareout(Xd_0__inst_mult_3_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_19 (
// Equation(s):
// Xd_0__inst_mult_0_54  = SUM(( !Xd_0__inst_mult_0_13_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_0_q ))) ) + ( Xd_0__inst_mult_0_52  ) + ( Xd_0__inst_mult_0_51  ))
// Xd_0__inst_mult_0_55  = CARRY(( !Xd_0__inst_mult_0_13_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_0_q ))) ) + ( Xd_0__inst_mult_0_52  ) + ( Xd_0__inst_mult_0_51  ))
// Xd_0__inst_mult_0_56  = SHARE((Xd_0__inst_mult_0_4_q  & (Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_13_q )))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_0_q ),
	.datac(!Xd_0__inst_mult_0_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_51 ),
	.sharein(Xd_0__inst_mult_0_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_54 ),
	.cout(Xd_0__inst_mult_0_55 ),
	.shareout(Xd_0__inst_mult_0_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_19 (
// Equation(s):
// Xd_0__inst_mult_1_54  = SUM(( !Xd_0__inst_mult_1_13_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_0_q ))) ) + ( Xd_0__inst_mult_1_52  ) + ( Xd_0__inst_mult_1_51  ))
// Xd_0__inst_mult_1_55  = CARRY(( !Xd_0__inst_mult_1_13_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_0_q ))) ) + ( Xd_0__inst_mult_1_52  ) + ( Xd_0__inst_mult_1_51  ))
// Xd_0__inst_mult_1_56  = SHARE((Xd_0__inst_mult_1_4_q  & (Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_13_q )))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_0_q ),
	.datac(!Xd_0__inst_mult_1_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_51 ),
	.sharein(Xd_0__inst_mult_1_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_54 ),
	.cout(Xd_0__inst_mult_1_55 ),
	.shareout(Xd_0__inst_mult_1_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_28_22 (
// Equation(s):
// Xd_0__inst_mult_28_67  = SUM(( !Xd_0__inst_mult_28_13_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_0_q ))) ) + ( Xd_0__inst_mult_28_65  ) + ( Xd_0__inst_mult_28_64  ))
// Xd_0__inst_mult_28_68  = CARRY(( !Xd_0__inst_mult_28_13_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_0_q ))) ) + ( Xd_0__inst_mult_28_65  ) + ( Xd_0__inst_mult_28_64  ))
// Xd_0__inst_mult_28_69  = SHARE((Xd_0__inst_mult_28_4_q  & (Xd_0__inst_mult_28_0_q  & Xd_0__inst_mult_28_13_q )))

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_0_q ),
	.datac(!Xd_0__inst_mult_28_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_64 ),
	.sharein(Xd_0__inst_mult_28_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_67 ),
	.cout(Xd_0__inst_mult_28_68 ),
	.shareout(Xd_0__inst_mult_28_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_29_20 (
// Equation(s):
// Xd_0__inst_mult_29_59  = SUM(( !Xd_0__inst_mult_29_13_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_0_q ))) ) + ( Xd_0__inst_mult_29_57  ) + ( Xd_0__inst_mult_29_56  ))
// Xd_0__inst_mult_29_60  = CARRY(( !Xd_0__inst_mult_29_13_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_0_q ))) ) + ( Xd_0__inst_mult_29_57  ) + ( Xd_0__inst_mult_29_56  ))
// Xd_0__inst_mult_29_61  = SHARE((Xd_0__inst_mult_29_4_q  & (Xd_0__inst_mult_29_0_q  & Xd_0__inst_mult_29_13_q )))

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_0_q ),
	.datac(!Xd_0__inst_mult_29_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_56 ),
	.sharein(Xd_0__inst_mult_29_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_59 ),
	.cout(Xd_0__inst_mult_29_60 ),
	.shareout(Xd_0__inst_mult_29_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_26_22 (
// Equation(s):
// Xd_0__inst_mult_26_67  = SUM(( !Xd_0__inst_mult_26_13_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_0_q ))) ) + ( Xd_0__inst_mult_26_65  ) + ( Xd_0__inst_mult_26_64  ))
// Xd_0__inst_mult_26_68  = CARRY(( !Xd_0__inst_mult_26_13_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_0_q ))) ) + ( Xd_0__inst_mult_26_65  ) + ( Xd_0__inst_mult_26_64  ))
// Xd_0__inst_mult_26_69  = SHARE((Xd_0__inst_mult_26_4_q  & (Xd_0__inst_mult_26_0_q  & Xd_0__inst_mult_26_13_q )))

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_0_q ),
	.datac(!Xd_0__inst_mult_26_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_64 ),
	.sharein(Xd_0__inst_mult_26_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_67 ),
	.cout(Xd_0__inst_mult_26_68 ),
	.shareout(Xd_0__inst_mult_26_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_27_20 (
// Equation(s):
// Xd_0__inst_mult_27_59  = SUM(( !Xd_0__inst_mult_27_13_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_0_q ))) ) + ( Xd_0__inst_mult_27_57  ) + ( Xd_0__inst_mult_27_56  ))
// Xd_0__inst_mult_27_60  = CARRY(( !Xd_0__inst_mult_27_13_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_0_q ))) ) + ( Xd_0__inst_mult_27_57  ) + ( Xd_0__inst_mult_27_56  ))
// Xd_0__inst_mult_27_61  = SHARE((Xd_0__inst_mult_27_4_q  & (Xd_0__inst_mult_27_0_q  & Xd_0__inst_mult_27_13_q )))

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_0_q ),
	.datac(!Xd_0__inst_mult_27_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_56 ),
	.sharein(Xd_0__inst_mult_27_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_59 ),
	.cout(Xd_0__inst_mult_27_60 ),
	.shareout(Xd_0__inst_mult_27_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_24_22 (
// Equation(s):
// Xd_0__inst_mult_24_67  = SUM(( !Xd_0__inst_mult_24_13_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_0_q ))) ) + ( Xd_0__inst_mult_24_65  ) + ( Xd_0__inst_mult_24_64  ))
// Xd_0__inst_mult_24_68  = CARRY(( !Xd_0__inst_mult_24_13_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_0_q ))) ) + ( Xd_0__inst_mult_24_65  ) + ( Xd_0__inst_mult_24_64  ))
// Xd_0__inst_mult_24_69  = SHARE((Xd_0__inst_mult_24_4_q  & (Xd_0__inst_mult_24_0_q  & Xd_0__inst_mult_24_13_q )))

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_0_q ),
	.datac(!Xd_0__inst_mult_24_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_64 ),
	.sharein(Xd_0__inst_mult_24_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_67 ),
	.cout(Xd_0__inst_mult_24_68 ),
	.shareout(Xd_0__inst_mult_24_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_25_20 (
// Equation(s):
// Xd_0__inst_mult_25_59  = SUM(( !Xd_0__inst_mult_25_13_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_0_q ))) ) + ( Xd_0__inst_mult_25_57  ) + ( Xd_0__inst_mult_25_56  ))
// Xd_0__inst_mult_25_60  = CARRY(( !Xd_0__inst_mult_25_13_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_0_q ))) ) + ( Xd_0__inst_mult_25_57  ) + ( Xd_0__inst_mult_25_56  ))
// Xd_0__inst_mult_25_61  = SHARE((Xd_0__inst_mult_25_4_q  & (Xd_0__inst_mult_25_0_q  & Xd_0__inst_mult_25_13_q )))

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_0_q ),
	.datac(!Xd_0__inst_mult_25_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_56 ),
	.sharein(Xd_0__inst_mult_25_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_59 ),
	.cout(Xd_0__inst_mult_25_60 ),
	.shareout(Xd_0__inst_mult_25_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_22_22 (
// Equation(s):
// Xd_0__inst_mult_22_67  = SUM(( !Xd_0__inst_mult_22_13_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_0_q ))) ) + ( Xd_0__inst_mult_22_65  ) + ( Xd_0__inst_mult_22_64  ))
// Xd_0__inst_mult_22_68  = CARRY(( !Xd_0__inst_mult_22_13_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_0_q ))) ) + ( Xd_0__inst_mult_22_65  ) + ( Xd_0__inst_mult_22_64  ))
// Xd_0__inst_mult_22_69  = SHARE((Xd_0__inst_mult_22_4_q  & (Xd_0__inst_mult_22_0_q  & Xd_0__inst_mult_22_13_q )))

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_0_q ),
	.datac(!Xd_0__inst_mult_22_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_64 ),
	.sharein(Xd_0__inst_mult_22_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_67 ),
	.cout(Xd_0__inst_mult_22_68 ),
	.shareout(Xd_0__inst_mult_22_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_23_22 (
// Equation(s):
// Xd_0__inst_mult_23_67  = SUM(( !Xd_0__inst_mult_23_13_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_0_q ))) ) + ( Xd_0__inst_mult_23_65  ) + ( Xd_0__inst_mult_23_64  ))
// Xd_0__inst_mult_23_68  = CARRY(( !Xd_0__inst_mult_23_13_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_0_q ))) ) + ( Xd_0__inst_mult_23_65  ) + ( Xd_0__inst_mult_23_64  ))
// Xd_0__inst_mult_23_69  = SHARE((Xd_0__inst_mult_23_4_q  & (Xd_0__inst_mult_23_0_q  & Xd_0__inst_mult_23_13_q )))

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_0_q ),
	.datac(!Xd_0__inst_mult_23_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_64 ),
	.sharein(Xd_0__inst_mult_23_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_67 ),
	.cout(Xd_0__inst_mult_23_68 ),
	.shareout(Xd_0__inst_mult_23_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_20_22 (
// Equation(s):
// Xd_0__inst_mult_20_67  = SUM(( !Xd_0__inst_mult_20_13_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_0_q ))) ) + ( Xd_0__inst_mult_20_65  ) + ( Xd_0__inst_mult_20_64  ))
// Xd_0__inst_mult_20_68  = CARRY(( !Xd_0__inst_mult_20_13_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_0_q ))) ) + ( Xd_0__inst_mult_20_65  ) + ( Xd_0__inst_mult_20_64  ))
// Xd_0__inst_mult_20_69  = SHARE((Xd_0__inst_mult_20_4_q  & (Xd_0__inst_mult_20_0_q  & Xd_0__inst_mult_20_13_q )))

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_0_q ),
	.datac(!Xd_0__inst_mult_20_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_64 ),
	.sharein(Xd_0__inst_mult_20_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_67 ),
	.cout(Xd_0__inst_mult_20_68 ),
	.shareout(Xd_0__inst_mult_20_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_21_18 (
// Equation(s):
// Xd_0__inst_mult_21_51  = SUM(( !Xd_0__inst_mult_21_13_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_0_q ))) ) + ( Xd_0__inst_mult_21_49  ) + ( Xd_0__inst_mult_21_48  ))
// Xd_0__inst_mult_21_52  = CARRY(( !Xd_0__inst_mult_21_13_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_0_q ))) ) + ( Xd_0__inst_mult_21_49  ) + ( Xd_0__inst_mult_21_48  ))
// Xd_0__inst_mult_21_53  = SHARE((Xd_0__inst_mult_21_4_q  & (Xd_0__inst_mult_21_0_q  & Xd_0__inst_mult_21_13_q )))

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_0_q ),
	.datac(!Xd_0__inst_mult_21_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_48 ),
	.sharein(Xd_0__inst_mult_21_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_51 ),
	.cout(Xd_0__inst_mult_21_52 ),
	.shareout(Xd_0__inst_mult_21_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_18_18 (
// Equation(s):
// Xd_0__inst_mult_18_50  = SUM(( !Xd_0__inst_mult_18_13_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_0_q ))) ) + ( Xd_0__inst_mult_18_48  ) + ( Xd_0__inst_mult_18_47  ))
// Xd_0__inst_mult_18_51  = CARRY(( !Xd_0__inst_mult_18_13_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_0_q ))) ) + ( Xd_0__inst_mult_18_48  ) + ( Xd_0__inst_mult_18_47  ))
// Xd_0__inst_mult_18_52  = SHARE((Xd_0__inst_mult_18_4_q  & (Xd_0__inst_mult_18_0_q  & Xd_0__inst_mult_18_13_q )))

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_0_q ),
	.datac(!Xd_0__inst_mult_18_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_47 ),
	.sharein(Xd_0__inst_mult_18_48 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_50 ),
	.cout(Xd_0__inst_mult_18_51 ),
	.shareout(Xd_0__inst_mult_18_52 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_19_21 (
// Equation(s):
// Xd_0__inst_mult_19_63  = SUM(( !Xd_0__inst_mult_19_13_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_0_q ))) ) + ( Xd_0__inst_mult_19_61  ) + ( Xd_0__inst_mult_19_60  ))
// Xd_0__inst_mult_19_64  = CARRY(( !Xd_0__inst_mult_19_13_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_0_q ))) ) + ( Xd_0__inst_mult_19_61  ) + ( Xd_0__inst_mult_19_60  ))
// Xd_0__inst_mult_19_65  = SHARE((Xd_0__inst_mult_19_4_q  & (Xd_0__inst_mult_19_0_q  & Xd_0__inst_mult_19_13_q )))

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_0_q ),
	.datac(!Xd_0__inst_mult_19_13_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_60 ),
	.sharein(Xd_0__inst_mult_19_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_63 ),
	.cout(Xd_0__inst_mult_19_64 ),
	.shareout(Xd_0__inst_mult_19_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_16_19 (
// Equation(s):
// Xd_0__inst_mult_16_54  = SUM(( !Xd_0__inst_mult_16_15_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_14_q ))) ) + ( Xd_0__inst_mult_16_52  ) + ( Xd_0__inst_mult_16_51  ))
// Xd_0__inst_mult_16_55  = CARRY(( !Xd_0__inst_mult_16_15_q  $ (((!Xd_0__inst_mult_16_4_q ) # (!Xd_0__inst_mult_16_14_q ))) ) + ( Xd_0__inst_mult_16_52  ) + ( Xd_0__inst_mult_16_51  ))
// Xd_0__inst_mult_16_56  = SHARE((Xd_0__inst_mult_16_4_q  & (Xd_0__inst_mult_16_14_q  & Xd_0__inst_mult_16_15_q )))

	.dataa(!Xd_0__inst_mult_16_4_q ),
	.datab(!Xd_0__inst_mult_16_14_q ),
	.datac(!Xd_0__inst_mult_16_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_51 ),
	.sharein(Xd_0__inst_mult_16_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_54 ),
	.cout(Xd_0__inst_mult_16_55 ),
	.shareout(Xd_0__inst_mult_16_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_17_19 (
// Equation(s):
// Xd_0__inst_mult_17_55  = SUM(( !Xd_0__inst_mult_17_15_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_14_q ))) ) + ( Xd_0__inst_mult_17_53  ) + ( Xd_0__inst_mult_17_52  ))
// Xd_0__inst_mult_17_56  = CARRY(( !Xd_0__inst_mult_17_15_q  $ (((!Xd_0__inst_mult_17_4_q ) # (!Xd_0__inst_mult_17_14_q ))) ) + ( Xd_0__inst_mult_17_53  ) + ( Xd_0__inst_mult_17_52  ))
// Xd_0__inst_mult_17_57  = SHARE((Xd_0__inst_mult_17_4_q  & (Xd_0__inst_mult_17_14_q  & Xd_0__inst_mult_17_15_q )))

	.dataa(!Xd_0__inst_mult_17_4_q ),
	.datab(!Xd_0__inst_mult_17_14_q ),
	.datac(!Xd_0__inst_mult_17_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_52 ),
	.sharein(Xd_0__inst_mult_17_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_55 ),
	.cout(Xd_0__inst_mult_17_56 ),
	.shareout(Xd_0__inst_mult_17_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_14_19 (
// Equation(s):
// Xd_0__inst_mult_14_54  = SUM(( !Xd_0__inst_mult_14_15_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_14_q ))) ) + ( Xd_0__inst_mult_14_52  ) + ( Xd_0__inst_mult_14_51  ))
// Xd_0__inst_mult_14_55  = CARRY(( !Xd_0__inst_mult_14_15_q  $ (((!Xd_0__inst_mult_14_4_q ) # (!Xd_0__inst_mult_14_14_q ))) ) + ( Xd_0__inst_mult_14_52  ) + ( Xd_0__inst_mult_14_51  ))
// Xd_0__inst_mult_14_56  = SHARE((Xd_0__inst_mult_14_4_q  & (Xd_0__inst_mult_14_14_q  & Xd_0__inst_mult_14_15_q )))

	.dataa(!Xd_0__inst_mult_14_4_q ),
	.datab(!Xd_0__inst_mult_14_14_q ),
	.datac(!Xd_0__inst_mult_14_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_51 ),
	.sharein(Xd_0__inst_mult_14_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_54 ),
	.cout(Xd_0__inst_mult_14_55 ),
	.shareout(Xd_0__inst_mult_14_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_15_19 (
// Equation(s):
// Xd_0__inst_mult_15_55  = SUM(( !Xd_0__inst_mult_15_15_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_14_q ))) ) + ( Xd_0__inst_mult_15_53  ) + ( Xd_0__inst_mult_15_52  ))
// Xd_0__inst_mult_15_56  = CARRY(( !Xd_0__inst_mult_15_15_q  $ (((!Xd_0__inst_mult_15_4_q ) # (!Xd_0__inst_mult_15_14_q ))) ) + ( Xd_0__inst_mult_15_53  ) + ( Xd_0__inst_mult_15_52  ))
// Xd_0__inst_mult_15_57  = SHARE((Xd_0__inst_mult_15_4_q  & (Xd_0__inst_mult_15_14_q  & Xd_0__inst_mult_15_15_q )))

	.dataa(!Xd_0__inst_mult_15_4_q ),
	.datab(!Xd_0__inst_mult_15_14_q ),
	.datac(!Xd_0__inst_mult_15_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_52 ),
	.sharein(Xd_0__inst_mult_15_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_55 ),
	.cout(Xd_0__inst_mult_15_56 ),
	.shareout(Xd_0__inst_mult_15_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_12_19 (
// Equation(s):
// Xd_0__inst_mult_12_54  = SUM(( !Xd_0__inst_mult_12_15_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_14_q ))) ) + ( Xd_0__inst_mult_12_52  ) + ( Xd_0__inst_mult_12_51  ))
// Xd_0__inst_mult_12_55  = CARRY(( !Xd_0__inst_mult_12_15_q  $ (((!Xd_0__inst_mult_12_4_q ) # (!Xd_0__inst_mult_12_14_q ))) ) + ( Xd_0__inst_mult_12_52  ) + ( Xd_0__inst_mult_12_51  ))
// Xd_0__inst_mult_12_56  = SHARE((Xd_0__inst_mult_12_4_q  & (Xd_0__inst_mult_12_14_q  & Xd_0__inst_mult_12_15_q )))

	.dataa(!Xd_0__inst_mult_12_4_q ),
	.datab(!Xd_0__inst_mult_12_14_q ),
	.datac(!Xd_0__inst_mult_12_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_51 ),
	.sharein(Xd_0__inst_mult_12_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_54 ),
	.cout(Xd_0__inst_mult_12_55 ),
	.shareout(Xd_0__inst_mult_12_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_13_19 (
// Equation(s):
// Xd_0__inst_mult_13_55  = SUM(( !Xd_0__inst_mult_13_15_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_14_q ))) ) + ( Xd_0__inst_mult_13_53  ) + ( Xd_0__inst_mult_13_52  ))
// Xd_0__inst_mult_13_56  = CARRY(( !Xd_0__inst_mult_13_15_q  $ (((!Xd_0__inst_mult_13_4_q ) # (!Xd_0__inst_mult_13_14_q ))) ) + ( Xd_0__inst_mult_13_53  ) + ( Xd_0__inst_mult_13_52  ))
// Xd_0__inst_mult_13_57  = SHARE((Xd_0__inst_mult_13_4_q  & (Xd_0__inst_mult_13_14_q  & Xd_0__inst_mult_13_15_q )))

	.dataa(!Xd_0__inst_mult_13_4_q ),
	.datab(!Xd_0__inst_mult_13_14_q ),
	.datac(!Xd_0__inst_mult_13_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_52 ),
	.sharein(Xd_0__inst_mult_13_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_55 ),
	.cout(Xd_0__inst_mult_13_56 ),
	.shareout(Xd_0__inst_mult_13_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_10_19 (
// Equation(s):
// Xd_0__inst_mult_10_54  = SUM(( !Xd_0__inst_mult_10_15_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_14_q ))) ) + ( Xd_0__inst_mult_10_52  ) + ( Xd_0__inst_mult_10_51  ))
// Xd_0__inst_mult_10_55  = CARRY(( !Xd_0__inst_mult_10_15_q  $ (((!Xd_0__inst_mult_10_4_q ) # (!Xd_0__inst_mult_10_14_q ))) ) + ( Xd_0__inst_mult_10_52  ) + ( Xd_0__inst_mult_10_51  ))
// Xd_0__inst_mult_10_56  = SHARE((Xd_0__inst_mult_10_4_q  & (Xd_0__inst_mult_10_14_q  & Xd_0__inst_mult_10_15_q )))

	.dataa(!Xd_0__inst_mult_10_4_q ),
	.datab(!Xd_0__inst_mult_10_14_q ),
	.datac(!Xd_0__inst_mult_10_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_51 ),
	.sharein(Xd_0__inst_mult_10_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_54 ),
	.cout(Xd_0__inst_mult_10_55 ),
	.shareout(Xd_0__inst_mult_10_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_11_21 (
// Equation(s):
// Xd_0__inst_mult_11_63  = SUM(( !Xd_0__inst_mult_11_15_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_14_q ))) ) + ( Xd_0__inst_mult_11_61  ) + ( Xd_0__inst_mult_11_60  ))
// Xd_0__inst_mult_11_64  = CARRY(( !Xd_0__inst_mult_11_15_q  $ (((!Xd_0__inst_mult_11_4_q ) # (!Xd_0__inst_mult_11_14_q ))) ) + ( Xd_0__inst_mult_11_61  ) + ( Xd_0__inst_mult_11_60  ))
// Xd_0__inst_mult_11_65  = SHARE((Xd_0__inst_mult_11_4_q  & (Xd_0__inst_mult_11_14_q  & Xd_0__inst_mult_11_15_q )))

	.dataa(!Xd_0__inst_mult_11_4_q ),
	.datab(!Xd_0__inst_mult_11_14_q ),
	.datac(!Xd_0__inst_mult_11_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_60 ),
	.sharein(Xd_0__inst_mult_11_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_63 ),
	.cout(Xd_0__inst_mult_11_64 ),
	.shareout(Xd_0__inst_mult_11_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_8_19 (
// Equation(s):
// Xd_0__inst_mult_8_54  = SUM(( !Xd_0__inst_mult_8_15_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_14_q ))) ) + ( Xd_0__inst_mult_8_52  ) + ( Xd_0__inst_mult_8_51  ))
// Xd_0__inst_mult_8_55  = CARRY(( !Xd_0__inst_mult_8_15_q  $ (((!Xd_0__inst_mult_8_4_q ) # (!Xd_0__inst_mult_8_14_q ))) ) + ( Xd_0__inst_mult_8_52  ) + ( Xd_0__inst_mult_8_51  ))
// Xd_0__inst_mult_8_56  = SHARE((Xd_0__inst_mult_8_4_q  & (Xd_0__inst_mult_8_14_q  & Xd_0__inst_mult_8_15_q )))

	.dataa(!Xd_0__inst_mult_8_4_q ),
	.datab(!Xd_0__inst_mult_8_14_q ),
	.datac(!Xd_0__inst_mult_8_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_51 ),
	.sharein(Xd_0__inst_mult_8_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_54 ),
	.cout(Xd_0__inst_mult_8_55 ),
	.shareout(Xd_0__inst_mult_8_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_9_19 (
// Equation(s):
// Xd_0__inst_mult_9_55  = SUM(( !Xd_0__inst_mult_9_15_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_14_q ))) ) + ( Xd_0__inst_mult_9_53  ) + ( Xd_0__inst_mult_9_52  ))
// Xd_0__inst_mult_9_56  = CARRY(( !Xd_0__inst_mult_9_15_q  $ (((!Xd_0__inst_mult_9_4_q ) # (!Xd_0__inst_mult_9_14_q ))) ) + ( Xd_0__inst_mult_9_53  ) + ( Xd_0__inst_mult_9_52  ))
// Xd_0__inst_mult_9_57  = SHARE((Xd_0__inst_mult_9_4_q  & (Xd_0__inst_mult_9_14_q  & Xd_0__inst_mult_9_15_q )))

	.dataa(!Xd_0__inst_mult_9_4_q ),
	.datab(!Xd_0__inst_mult_9_14_q ),
	.datac(!Xd_0__inst_mult_9_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_52 ),
	.sharein(Xd_0__inst_mult_9_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_55 ),
	.cout(Xd_0__inst_mult_9_56 ),
	.shareout(Xd_0__inst_mult_9_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_19 (
// Equation(s):
// Xd_0__inst_mult_6_53  = SUM(( !Xd_0__inst_mult_6_15_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_14_q ))) ) + ( Xd_0__inst_mult_6_51  ) + ( Xd_0__inst_mult_6_50  ))
// Xd_0__inst_mult_6_54  = CARRY(( !Xd_0__inst_mult_6_15_q  $ (((!Xd_0__inst_mult_6_4_q ) # (!Xd_0__inst_mult_6_14_q ))) ) + ( Xd_0__inst_mult_6_51  ) + ( Xd_0__inst_mult_6_50  ))
// Xd_0__inst_mult_6_55  = SHARE((Xd_0__inst_mult_6_4_q  & (Xd_0__inst_mult_6_14_q  & Xd_0__inst_mult_6_15_q )))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_14_q ),
	.datac(!Xd_0__inst_mult_6_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_50 ),
	.sharein(Xd_0__inst_mult_6_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_53 ),
	.cout(Xd_0__inst_mult_6_54 ),
	.shareout(Xd_0__inst_mult_6_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_19 (
// Equation(s):
// Xd_0__inst_mult_7_54  = SUM(( !Xd_0__inst_mult_7_15_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_14_q ))) ) + ( Xd_0__inst_mult_7_52  ) + ( Xd_0__inst_mult_7_51  ))
// Xd_0__inst_mult_7_55  = CARRY(( !Xd_0__inst_mult_7_15_q  $ (((!Xd_0__inst_mult_7_4_q ) # (!Xd_0__inst_mult_7_14_q ))) ) + ( Xd_0__inst_mult_7_52  ) + ( Xd_0__inst_mult_7_51  ))
// Xd_0__inst_mult_7_56  = SHARE((Xd_0__inst_mult_7_4_q  & (Xd_0__inst_mult_7_14_q  & Xd_0__inst_mult_7_15_q )))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_14_q ),
	.datac(!Xd_0__inst_mult_7_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_51 ),
	.sharein(Xd_0__inst_mult_7_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_54 ),
	.cout(Xd_0__inst_mult_7_55 ),
	.shareout(Xd_0__inst_mult_7_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_19 (
// Equation(s):
// Xd_0__inst_mult_4_53  = SUM(( !Xd_0__inst_mult_4_15_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_14_q ))) ) + ( Xd_0__inst_mult_4_51  ) + ( Xd_0__inst_mult_4_50  ))
// Xd_0__inst_mult_4_54  = CARRY(( !Xd_0__inst_mult_4_15_q  $ (((!Xd_0__inst_mult_4_4_q ) # (!Xd_0__inst_mult_4_14_q ))) ) + ( Xd_0__inst_mult_4_51  ) + ( Xd_0__inst_mult_4_50  ))
// Xd_0__inst_mult_4_55  = SHARE((Xd_0__inst_mult_4_4_q  & (Xd_0__inst_mult_4_14_q  & Xd_0__inst_mult_4_15_q )))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_14_q ),
	.datac(!Xd_0__inst_mult_4_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_50 ),
	.sharein(Xd_0__inst_mult_4_51 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_53 ),
	.cout(Xd_0__inst_mult_4_54 ),
	.shareout(Xd_0__inst_mult_4_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_19 (
// Equation(s):
// Xd_0__inst_mult_5_54  = SUM(( !Xd_0__inst_mult_5_15_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_14_q ))) ) + ( Xd_0__inst_mult_5_52  ) + ( Xd_0__inst_mult_5_51  ))
// Xd_0__inst_mult_5_55  = CARRY(( !Xd_0__inst_mult_5_15_q  $ (((!Xd_0__inst_mult_5_4_q ) # (!Xd_0__inst_mult_5_14_q ))) ) + ( Xd_0__inst_mult_5_52  ) + ( Xd_0__inst_mult_5_51  ))
// Xd_0__inst_mult_5_56  = SHARE((Xd_0__inst_mult_5_4_q  & (Xd_0__inst_mult_5_14_q  & Xd_0__inst_mult_5_15_q )))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_14_q ),
	.datac(!Xd_0__inst_mult_5_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_51 ),
	.sharein(Xd_0__inst_mult_5_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_54 ),
	.cout(Xd_0__inst_mult_5_55 ),
	.shareout(Xd_0__inst_mult_5_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_20 (
// Equation(s):
// Xd_0__inst_mult_2_58  = SUM(( !Xd_0__inst_mult_2_15_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_14_q ))) ) + ( Xd_0__inst_mult_2_56  ) + ( Xd_0__inst_mult_2_55  ))
// Xd_0__inst_mult_2_59  = CARRY(( !Xd_0__inst_mult_2_15_q  $ (((!Xd_0__inst_mult_2_4_q ) # (!Xd_0__inst_mult_2_14_q ))) ) + ( Xd_0__inst_mult_2_56  ) + ( Xd_0__inst_mult_2_55  ))
// Xd_0__inst_mult_2_60  = SHARE((Xd_0__inst_mult_2_4_q  & (Xd_0__inst_mult_2_14_q  & Xd_0__inst_mult_2_15_q )))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_14_q ),
	.datac(!Xd_0__inst_mult_2_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_55 ),
	.sharein(Xd_0__inst_mult_2_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_58 ),
	.cout(Xd_0__inst_mult_2_59 ),
	.shareout(Xd_0__inst_mult_2_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_20 (
// Equation(s):
// Xd_0__inst_mult_3_58  = SUM(( !Xd_0__inst_mult_3_15_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_14_q ))) ) + ( Xd_0__inst_mult_3_56  ) + ( Xd_0__inst_mult_3_55  ))
// Xd_0__inst_mult_3_59  = CARRY(( !Xd_0__inst_mult_3_15_q  $ (((!Xd_0__inst_mult_3_4_q ) # (!Xd_0__inst_mult_3_14_q ))) ) + ( Xd_0__inst_mult_3_56  ) + ( Xd_0__inst_mult_3_55  ))
// Xd_0__inst_mult_3_60  = SHARE((Xd_0__inst_mult_3_4_q  & (Xd_0__inst_mult_3_14_q  & Xd_0__inst_mult_3_15_q )))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_14_q ),
	.datac(!Xd_0__inst_mult_3_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_55 ),
	.sharein(Xd_0__inst_mult_3_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_58 ),
	.cout(Xd_0__inst_mult_3_59 ),
	.shareout(Xd_0__inst_mult_3_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_20 (
// Equation(s):
// Xd_0__inst_mult_0_58  = SUM(( !Xd_0__inst_mult_0_15_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_14_q ))) ) + ( Xd_0__inst_mult_0_56  ) + ( Xd_0__inst_mult_0_55  ))
// Xd_0__inst_mult_0_59  = CARRY(( !Xd_0__inst_mult_0_15_q  $ (((!Xd_0__inst_mult_0_4_q ) # (!Xd_0__inst_mult_0_14_q ))) ) + ( Xd_0__inst_mult_0_56  ) + ( Xd_0__inst_mult_0_55  ))
// Xd_0__inst_mult_0_60  = SHARE((Xd_0__inst_mult_0_4_q  & (Xd_0__inst_mult_0_14_q  & Xd_0__inst_mult_0_15_q )))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_14_q ),
	.datac(!Xd_0__inst_mult_0_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_55 ),
	.sharein(Xd_0__inst_mult_0_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_58 ),
	.cout(Xd_0__inst_mult_0_59 ),
	.shareout(Xd_0__inst_mult_0_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_20 (
// Equation(s):
// Xd_0__inst_mult_1_58  = SUM(( !Xd_0__inst_mult_1_15_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_14_q ))) ) + ( Xd_0__inst_mult_1_56  ) + ( Xd_0__inst_mult_1_55  ))
// Xd_0__inst_mult_1_59  = CARRY(( !Xd_0__inst_mult_1_15_q  $ (((!Xd_0__inst_mult_1_4_q ) # (!Xd_0__inst_mult_1_14_q ))) ) + ( Xd_0__inst_mult_1_56  ) + ( Xd_0__inst_mult_1_55  ))
// Xd_0__inst_mult_1_60  = SHARE((Xd_0__inst_mult_1_4_q  & (Xd_0__inst_mult_1_14_q  & Xd_0__inst_mult_1_15_q )))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_14_q ),
	.datac(!Xd_0__inst_mult_1_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_55 ),
	.sharein(Xd_0__inst_mult_1_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_58 ),
	.cout(Xd_0__inst_mult_1_59 ),
	.shareout(Xd_0__inst_mult_1_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_28_23 (
// Equation(s):
// Xd_0__inst_mult_28_71  = SUM(( !Xd_0__inst_mult_28_15_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_14_q ))) ) + ( Xd_0__inst_mult_28_69  ) + ( Xd_0__inst_mult_28_68  ))
// Xd_0__inst_mult_28_72  = CARRY(( !Xd_0__inst_mult_28_15_q  $ (((!Xd_0__inst_mult_28_4_q ) # (!Xd_0__inst_mult_28_14_q ))) ) + ( Xd_0__inst_mult_28_69  ) + ( Xd_0__inst_mult_28_68  ))
// Xd_0__inst_mult_28_73  = SHARE((Xd_0__inst_mult_28_4_q  & (Xd_0__inst_mult_28_14_q  & Xd_0__inst_mult_28_15_q )))

	.dataa(!Xd_0__inst_mult_28_4_q ),
	.datab(!Xd_0__inst_mult_28_14_q ),
	.datac(!Xd_0__inst_mult_28_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_68 ),
	.sharein(Xd_0__inst_mult_28_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_71 ),
	.cout(Xd_0__inst_mult_28_72 ),
	.shareout(Xd_0__inst_mult_28_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_29_21 (
// Equation(s):
// Xd_0__inst_mult_29_63  = SUM(( !Xd_0__inst_mult_29_15_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_14_q ))) ) + ( Xd_0__inst_mult_29_61  ) + ( Xd_0__inst_mult_29_60  ))
// Xd_0__inst_mult_29_64  = CARRY(( !Xd_0__inst_mult_29_15_q  $ (((!Xd_0__inst_mult_29_4_q ) # (!Xd_0__inst_mult_29_14_q ))) ) + ( Xd_0__inst_mult_29_61  ) + ( Xd_0__inst_mult_29_60  ))
// Xd_0__inst_mult_29_65  = SHARE((Xd_0__inst_mult_29_4_q  & (Xd_0__inst_mult_29_14_q  & Xd_0__inst_mult_29_15_q )))

	.dataa(!Xd_0__inst_mult_29_4_q ),
	.datab(!Xd_0__inst_mult_29_14_q ),
	.datac(!Xd_0__inst_mult_29_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_60 ),
	.sharein(Xd_0__inst_mult_29_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_63 ),
	.cout(Xd_0__inst_mult_29_64 ),
	.shareout(Xd_0__inst_mult_29_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_26_23 (
// Equation(s):
// Xd_0__inst_mult_26_71  = SUM(( !Xd_0__inst_mult_26_15_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_14_q ))) ) + ( Xd_0__inst_mult_26_69  ) + ( Xd_0__inst_mult_26_68  ))
// Xd_0__inst_mult_26_72  = CARRY(( !Xd_0__inst_mult_26_15_q  $ (((!Xd_0__inst_mult_26_4_q ) # (!Xd_0__inst_mult_26_14_q ))) ) + ( Xd_0__inst_mult_26_69  ) + ( Xd_0__inst_mult_26_68  ))
// Xd_0__inst_mult_26_73  = SHARE((Xd_0__inst_mult_26_4_q  & (Xd_0__inst_mult_26_14_q  & Xd_0__inst_mult_26_15_q )))

	.dataa(!Xd_0__inst_mult_26_4_q ),
	.datab(!Xd_0__inst_mult_26_14_q ),
	.datac(!Xd_0__inst_mult_26_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_68 ),
	.sharein(Xd_0__inst_mult_26_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_71 ),
	.cout(Xd_0__inst_mult_26_72 ),
	.shareout(Xd_0__inst_mult_26_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_27_21 (
// Equation(s):
// Xd_0__inst_mult_27_63  = SUM(( !Xd_0__inst_mult_27_15_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_14_q ))) ) + ( Xd_0__inst_mult_27_61  ) + ( Xd_0__inst_mult_27_60  ))
// Xd_0__inst_mult_27_64  = CARRY(( !Xd_0__inst_mult_27_15_q  $ (((!Xd_0__inst_mult_27_4_q ) # (!Xd_0__inst_mult_27_14_q ))) ) + ( Xd_0__inst_mult_27_61  ) + ( Xd_0__inst_mult_27_60  ))
// Xd_0__inst_mult_27_65  = SHARE((Xd_0__inst_mult_27_4_q  & (Xd_0__inst_mult_27_14_q  & Xd_0__inst_mult_27_15_q )))

	.dataa(!Xd_0__inst_mult_27_4_q ),
	.datab(!Xd_0__inst_mult_27_14_q ),
	.datac(!Xd_0__inst_mult_27_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_60 ),
	.sharein(Xd_0__inst_mult_27_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_63 ),
	.cout(Xd_0__inst_mult_27_64 ),
	.shareout(Xd_0__inst_mult_27_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_24_23 (
// Equation(s):
// Xd_0__inst_mult_24_71  = SUM(( !Xd_0__inst_mult_24_15_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_14_q ))) ) + ( Xd_0__inst_mult_24_69  ) + ( Xd_0__inst_mult_24_68  ))
// Xd_0__inst_mult_24_72  = CARRY(( !Xd_0__inst_mult_24_15_q  $ (((!Xd_0__inst_mult_24_4_q ) # (!Xd_0__inst_mult_24_14_q ))) ) + ( Xd_0__inst_mult_24_69  ) + ( Xd_0__inst_mult_24_68  ))
// Xd_0__inst_mult_24_73  = SHARE((Xd_0__inst_mult_24_4_q  & (Xd_0__inst_mult_24_14_q  & Xd_0__inst_mult_24_15_q )))

	.dataa(!Xd_0__inst_mult_24_4_q ),
	.datab(!Xd_0__inst_mult_24_14_q ),
	.datac(!Xd_0__inst_mult_24_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_68 ),
	.sharein(Xd_0__inst_mult_24_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_71 ),
	.cout(Xd_0__inst_mult_24_72 ),
	.shareout(Xd_0__inst_mult_24_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_25_21 (
// Equation(s):
// Xd_0__inst_mult_25_63  = SUM(( !Xd_0__inst_mult_25_15_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_14_q ))) ) + ( Xd_0__inst_mult_25_61  ) + ( Xd_0__inst_mult_25_60  ))
// Xd_0__inst_mult_25_64  = CARRY(( !Xd_0__inst_mult_25_15_q  $ (((!Xd_0__inst_mult_25_4_q ) # (!Xd_0__inst_mult_25_14_q ))) ) + ( Xd_0__inst_mult_25_61  ) + ( Xd_0__inst_mult_25_60  ))
// Xd_0__inst_mult_25_65  = SHARE((Xd_0__inst_mult_25_4_q  & (Xd_0__inst_mult_25_14_q  & Xd_0__inst_mult_25_15_q )))

	.dataa(!Xd_0__inst_mult_25_4_q ),
	.datab(!Xd_0__inst_mult_25_14_q ),
	.datac(!Xd_0__inst_mult_25_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_60 ),
	.sharein(Xd_0__inst_mult_25_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_63 ),
	.cout(Xd_0__inst_mult_25_64 ),
	.shareout(Xd_0__inst_mult_25_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_22_23 (
// Equation(s):
// Xd_0__inst_mult_22_71  = SUM(( !Xd_0__inst_mult_22_15_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_14_q ))) ) + ( Xd_0__inst_mult_22_69  ) + ( Xd_0__inst_mult_22_68  ))
// Xd_0__inst_mult_22_72  = CARRY(( !Xd_0__inst_mult_22_15_q  $ (((!Xd_0__inst_mult_22_4_q ) # (!Xd_0__inst_mult_22_14_q ))) ) + ( Xd_0__inst_mult_22_69  ) + ( Xd_0__inst_mult_22_68  ))
// Xd_0__inst_mult_22_73  = SHARE((Xd_0__inst_mult_22_4_q  & (Xd_0__inst_mult_22_14_q  & Xd_0__inst_mult_22_15_q )))

	.dataa(!Xd_0__inst_mult_22_4_q ),
	.datab(!Xd_0__inst_mult_22_14_q ),
	.datac(!Xd_0__inst_mult_22_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_68 ),
	.sharein(Xd_0__inst_mult_22_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_71 ),
	.cout(Xd_0__inst_mult_22_72 ),
	.shareout(Xd_0__inst_mult_22_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_23_23 (
// Equation(s):
// Xd_0__inst_mult_23_71  = SUM(( !Xd_0__inst_mult_23_15_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_14_q ))) ) + ( Xd_0__inst_mult_23_69  ) + ( Xd_0__inst_mult_23_68  ))
// Xd_0__inst_mult_23_72  = CARRY(( !Xd_0__inst_mult_23_15_q  $ (((!Xd_0__inst_mult_23_4_q ) # (!Xd_0__inst_mult_23_14_q ))) ) + ( Xd_0__inst_mult_23_69  ) + ( Xd_0__inst_mult_23_68  ))
// Xd_0__inst_mult_23_73  = SHARE((Xd_0__inst_mult_23_4_q  & (Xd_0__inst_mult_23_14_q  & Xd_0__inst_mult_23_15_q )))

	.dataa(!Xd_0__inst_mult_23_4_q ),
	.datab(!Xd_0__inst_mult_23_14_q ),
	.datac(!Xd_0__inst_mult_23_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_68 ),
	.sharein(Xd_0__inst_mult_23_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_71 ),
	.cout(Xd_0__inst_mult_23_72 ),
	.shareout(Xd_0__inst_mult_23_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_20_23 (
// Equation(s):
// Xd_0__inst_mult_20_71  = SUM(( !Xd_0__inst_mult_20_15_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_14_q ))) ) + ( Xd_0__inst_mult_20_69  ) + ( Xd_0__inst_mult_20_68  ))
// Xd_0__inst_mult_20_72  = CARRY(( !Xd_0__inst_mult_20_15_q  $ (((!Xd_0__inst_mult_20_4_q ) # (!Xd_0__inst_mult_20_14_q ))) ) + ( Xd_0__inst_mult_20_69  ) + ( Xd_0__inst_mult_20_68  ))
// Xd_0__inst_mult_20_73  = SHARE((Xd_0__inst_mult_20_4_q  & (Xd_0__inst_mult_20_14_q  & Xd_0__inst_mult_20_15_q )))

	.dataa(!Xd_0__inst_mult_20_4_q ),
	.datab(!Xd_0__inst_mult_20_14_q ),
	.datac(!Xd_0__inst_mult_20_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_68 ),
	.sharein(Xd_0__inst_mult_20_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_71 ),
	.cout(Xd_0__inst_mult_20_72 ),
	.shareout(Xd_0__inst_mult_20_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_21_19 (
// Equation(s):
// Xd_0__inst_mult_21_55  = SUM(( !Xd_0__inst_mult_21_15_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_14_q ))) ) + ( Xd_0__inst_mult_21_53  ) + ( Xd_0__inst_mult_21_52  ))
// Xd_0__inst_mult_21_56  = CARRY(( !Xd_0__inst_mult_21_15_q  $ (((!Xd_0__inst_mult_21_4_q ) # (!Xd_0__inst_mult_21_14_q ))) ) + ( Xd_0__inst_mult_21_53  ) + ( Xd_0__inst_mult_21_52  ))
// Xd_0__inst_mult_21_57  = SHARE((Xd_0__inst_mult_21_4_q  & (Xd_0__inst_mult_21_14_q  & Xd_0__inst_mult_21_15_q )))

	.dataa(!Xd_0__inst_mult_21_4_q ),
	.datab(!Xd_0__inst_mult_21_14_q ),
	.datac(!Xd_0__inst_mult_21_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_52 ),
	.sharein(Xd_0__inst_mult_21_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_55 ),
	.cout(Xd_0__inst_mult_21_56 ),
	.shareout(Xd_0__inst_mult_21_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_18_19 (
// Equation(s):
// Xd_0__inst_mult_18_54  = SUM(( !Xd_0__inst_mult_18_15_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_14_q ))) ) + ( Xd_0__inst_mult_18_52  ) + ( Xd_0__inst_mult_18_51  ))
// Xd_0__inst_mult_18_55  = CARRY(( !Xd_0__inst_mult_18_15_q  $ (((!Xd_0__inst_mult_18_4_q ) # (!Xd_0__inst_mult_18_14_q ))) ) + ( Xd_0__inst_mult_18_52  ) + ( Xd_0__inst_mult_18_51  ))
// Xd_0__inst_mult_18_56  = SHARE((Xd_0__inst_mult_18_4_q  & (Xd_0__inst_mult_18_14_q  & Xd_0__inst_mult_18_15_q )))

	.dataa(!Xd_0__inst_mult_18_4_q ),
	.datab(!Xd_0__inst_mult_18_14_q ),
	.datac(!Xd_0__inst_mult_18_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_51 ),
	.sharein(Xd_0__inst_mult_18_52 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_54 ),
	.cout(Xd_0__inst_mult_18_55 ),
	.shareout(Xd_0__inst_mult_18_56 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_19_22 (
// Equation(s):
// Xd_0__inst_mult_19_67  = SUM(( !Xd_0__inst_mult_19_15_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_14_q ))) ) + ( Xd_0__inst_mult_19_65  ) + ( Xd_0__inst_mult_19_64  ))
// Xd_0__inst_mult_19_68  = CARRY(( !Xd_0__inst_mult_19_15_q  $ (((!Xd_0__inst_mult_19_4_q ) # (!Xd_0__inst_mult_19_14_q ))) ) + ( Xd_0__inst_mult_19_65  ) + ( Xd_0__inst_mult_19_64  ))
// Xd_0__inst_mult_19_69  = SHARE((Xd_0__inst_mult_19_4_q  & (Xd_0__inst_mult_19_14_q  & Xd_0__inst_mult_19_15_q )))

	.dataa(!Xd_0__inst_mult_19_4_q ),
	.datab(!Xd_0__inst_mult_19_14_q ),
	.datac(!Xd_0__inst_mult_19_15_q ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_64 ),
	.sharein(Xd_0__inst_mult_19_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_67 ),
	.cout(Xd_0__inst_mult_19_68 ),
	.shareout(Xd_0__inst_mult_19_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_20 (
// Equation(s):
// Xd_0__inst_mult_17_59  = SUM(( GND ) + ( Xd_0__inst_mult_16_56  ) + ( Xd_0__inst_mult_16_55  ))
// Xd_0__inst_mult_17_60  = CARRY(( GND ) + ( Xd_0__inst_mult_16_56  ) + ( Xd_0__inst_mult_16_55  ))
// Xd_0__inst_mult_17_61  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_17_0_q ),
	.datab(!Xd_0__inst_mult_17_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_55 ),
	.sharein(Xd_0__inst_mult_16_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_59 ),
	.cout(Xd_0__inst_mult_17_60 ),
	.shareout(Xd_0__inst_mult_17_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_21 (
// Equation(s):
// Xd_0__inst_mult_17_63  = SUM(( GND ) + ( Xd_0__inst_mult_17_57  ) + ( Xd_0__inst_mult_17_56  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_56 ),
	.sharein(Xd_0__inst_mult_17_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_20 (
// Equation(s):
// Xd_0__inst_mult_15_59  = SUM(( GND ) + ( Xd_0__inst_mult_14_56  ) + ( Xd_0__inst_mult_14_55  ))
// Xd_0__inst_mult_15_60  = CARRY(( GND ) + ( Xd_0__inst_mult_14_56  ) + ( Xd_0__inst_mult_14_55  ))
// Xd_0__inst_mult_15_61  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_55 ),
	.sharein(Xd_0__inst_mult_14_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_59 ),
	.cout(Xd_0__inst_mult_15_60 ),
	.shareout(Xd_0__inst_mult_15_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_21 (
// Equation(s):
// Xd_0__inst_mult_15_63  = SUM(( GND ) + ( Xd_0__inst_mult_15_57  ) + ( Xd_0__inst_mult_15_56  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_56 ),
	.sharein(Xd_0__inst_mult_15_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_20 (
// Equation(s):
// Xd_0__inst_mult_13_59  = SUM(( GND ) + ( Xd_0__inst_mult_12_56  ) + ( Xd_0__inst_mult_12_55  ))
// Xd_0__inst_mult_13_60  = CARRY(( GND ) + ( Xd_0__inst_mult_12_56  ) + ( Xd_0__inst_mult_12_55  ))
// Xd_0__inst_mult_13_61  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_55 ),
	.sharein(Xd_0__inst_mult_12_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_59 ),
	.cout(Xd_0__inst_mult_13_60 ),
	.shareout(Xd_0__inst_mult_13_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_21 (
// Equation(s):
// Xd_0__inst_mult_13_63  = SUM(( GND ) + ( Xd_0__inst_mult_13_57  ) + ( Xd_0__inst_mult_13_56  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_56 ),
	.sharein(Xd_0__inst_mult_13_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_20 (
// Equation(s):
// Xd_0__inst_mult_21_59  = SUM(( GND ) + ( Xd_0__inst_mult_10_56  ) + ( Xd_0__inst_mult_10_55  ))
// Xd_0__inst_mult_21_60  = CARRY(( GND ) + ( Xd_0__inst_mult_10_56  ) + ( Xd_0__inst_mult_10_55  ))
// Xd_0__inst_mult_21_61  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_21_0_q ),
	.datab(!Xd_0__inst_mult_21_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_55 ),
	.sharein(Xd_0__inst_mult_10_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_59 ),
	.cout(Xd_0__inst_mult_21_60 ),
	.shareout(Xd_0__inst_mult_21_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_22 (
// Equation(s):
// Xd_0__inst_mult_11_67  = SUM(( GND ) + ( Xd_0__inst_mult_11_65  ) + ( Xd_0__inst_mult_11_64  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_64 ),
	.sharein(Xd_0__inst_mult_11_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_67 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_20 (
// Equation(s):
// Xd_0__inst_mult_9_59  = SUM(( GND ) + ( Xd_0__inst_mult_8_56  ) + ( Xd_0__inst_mult_8_55  ))
// Xd_0__inst_mult_9_60  = CARRY(( GND ) + ( Xd_0__inst_mult_8_56  ) + ( Xd_0__inst_mult_8_55  ))
// Xd_0__inst_mult_9_61  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_55 ),
	.sharein(Xd_0__inst_mult_8_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_59 ),
	.cout(Xd_0__inst_mult_9_60 ),
	.shareout(Xd_0__inst_mult_9_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_21 (
// Equation(s):
// Xd_0__inst_mult_9_63  = SUM(( GND ) + ( Xd_0__inst_mult_9_57  ) + ( Xd_0__inst_mult_9_56  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_56 ),
	.sharein(Xd_0__inst_mult_9_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_20 (
// Equation(s):
// Xd_0__inst_mult_7_58  = SUM(( GND ) + ( Xd_0__inst_mult_6_55  ) + ( Xd_0__inst_mult_6_54  ))
// Xd_0__inst_mult_7_59  = CARRY(( GND ) + ( Xd_0__inst_mult_6_55  ) + ( Xd_0__inst_mult_6_54  ))
// Xd_0__inst_mult_7_60  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_54 ),
	.sharein(Xd_0__inst_mult_6_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_58 ),
	.cout(Xd_0__inst_mult_7_59 ),
	.shareout(Xd_0__inst_mult_7_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_21 (
// Equation(s):
// Xd_0__inst_mult_7_62  = SUM(( GND ) + ( Xd_0__inst_mult_7_56  ) + ( Xd_0__inst_mult_7_55  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_55 ),
	.sharein(Xd_0__inst_mult_7_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_20 (
// Equation(s):
// Xd_0__inst_mult_5_58  = SUM(( GND ) + ( Xd_0__inst_mult_4_55  ) + ( Xd_0__inst_mult_4_54  ))
// Xd_0__inst_mult_5_59  = CARRY(( GND ) + ( Xd_0__inst_mult_4_55  ) + ( Xd_0__inst_mult_4_54  ))
// Xd_0__inst_mult_5_60  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_54 ),
	.sharein(Xd_0__inst_mult_4_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_58 ),
	.cout(Xd_0__inst_mult_5_59 ),
	.shareout(Xd_0__inst_mult_5_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_21 (
// Equation(s):
// Xd_0__inst_mult_5_62  = SUM(( GND ) + ( Xd_0__inst_mult_5_56  ) + ( Xd_0__inst_mult_5_55  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_55 ),
	.sharein(Xd_0__inst_mult_5_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_21 (
// Equation(s):
// Xd_0__inst_mult_2_62  = SUM(( GND ) + ( Xd_0__inst_mult_2_60  ) + ( Xd_0__inst_mult_2_59  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_59 ),
	.sharein(Xd_0__inst_mult_2_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_21 (
// Equation(s):
// Xd_0__inst_mult_3_62  = SUM(( GND ) + ( Xd_0__inst_mult_3_60  ) + ( Xd_0__inst_mult_3_59  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_59 ),
	.sharein(Xd_0__inst_mult_3_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_21 (
// Equation(s):
// Xd_0__inst_mult_0_62  = SUM(( GND ) + ( Xd_0__inst_mult_0_60  ) + ( Xd_0__inst_mult_0_59  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_59 ),
	.sharein(Xd_0__inst_mult_0_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_21 (
// Equation(s):
// Xd_0__inst_mult_1_62  = SUM(( GND ) + ( Xd_0__inst_mult_1_60  ) + ( Xd_0__inst_mult_1_59  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_59 ),
	.sharein(Xd_0__inst_mult_1_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_62 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_24 (
// Equation(s):
// Xd_0__inst_mult_28_75  = SUM(( GND ) + ( Xd_0__inst_mult_28_73  ) + ( Xd_0__inst_mult_28_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_72 ),
	.sharein(Xd_0__inst_mult_28_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_22 (
// Equation(s):
// Xd_0__inst_mult_29_67  = SUM(( GND ) + ( Xd_0__inst_mult_29_65  ) + ( Xd_0__inst_mult_29_64  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_64 ),
	.sharein(Xd_0__inst_mult_29_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_67 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_24 (
// Equation(s):
// Xd_0__inst_mult_26_75  = SUM(( GND ) + ( Xd_0__inst_mult_26_73  ) + ( Xd_0__inst_mult_26_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_72 ),
	.sharein(Xd_0__inst_mult_26_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_22 (
// Equation(s):
// Xd_0__inst_mult_27_67  = SUM(( GND ) + ( Xd_0__inst_mult_27_65  ) + ( Xd_0__inst_mult_27_64  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_64 ),
	.sharein(Xd_0__inst_mult_27_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_67 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_24 (
// Equation(s):
// Xd_0__inst_mult_24_75  = SUM(( GND ) + ( Xd_0__inst_mult_24_73  ) + ( Xd_0__inst_mult_24_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_72 ),
	.sharein(Xd_0__inst_mult_24_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_22 (
// Equation(s):
// Xd_0__inst_mult_25_67  = SUM(( GND ) + ( Xd_0__inst_mult_25_65  ) + ( Xd_0__inst_mult_25_64  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_64 ),
	.sharein(Xd_0__inst_mult_25_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_67 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_24 (
// Equation(s):
// Xd_0__inst_mult_22_75  = SUM(( GND ) + ( Xd_0__inst_mult_22_73  ) + ( Xd_0__inst_mult_22_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_72 ),
	.sharein(Xd_0__inst_mult_22_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_24 (
// Equation(s):
// Xd_0__inst_mult_23_75  = SUM(( GND ) + ( Xd_0__inst_mult_23_73  ) + ( Xd_0__inst_mult_23_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_72 ),
	.sharein(Xd_0__inst_mult_23_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_24 (
// Equation(s):
// Xd_0__inst_mult_20_75  = SUM(( GND ) + ( Xd_0__inst_mult_20_73  ) + ( Xd_0__inst_mult_20_72  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_72 ),
	.sharein(Xd_0__inst_mult_20_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_21 (
// Equation(s):
// Xd_0__inst_mult_21_63  = SUM(( GND ) + ( Xd_0__inst_mult_21_57  ) + ( Xd_0__inst_mult_21_56  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_56 ),
	.sharein(Xd_0__inst_mult_21_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_63 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_23 (
// Equation(s):
// Xd_0__inst_mult_19_71  = SUM(( GND ) + ( Xd_0__inst_mult_18_56  ) + ( Xd_0__inst_mult_18_55  ))
// Xd_0__inst_mult_19_72  = CARRY(( GND ) + ( Xd_0__inst_mult_18_56  ) + ( Xd_0__inst_mult_18_55  ))
// Xd_0__inst_mult_19_73  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_19_0_q ),
	.datab(!Xd_0__inst_mult_19_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_55 ),
	.sharein(Xd_0__inst_mult_18_56 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_71 ),
	.cout(Xd_0__inst_mult_19_72 ),
	.shareout(Xd_0__inst_mult_19_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_24 (
// Equation(s):
// Xd_0__inst_mult_19_75  = SUM(( GND ) + ( Xd_0__inst_mult_19_69  ) + ( Xd_0__inst_mult_19_68  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_68 ),
	.sharein(Xd_0__inst_mult_19_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_75 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_20 (
// Equation(s):
// Xd_0__inst_mult_16_58  = SUM(( (din_a[96] & din_b[96]) ) + ( Xd_0__inst_mult_22_97  ) + ( Xd_0__inst_mult_22_96  ))
// Xd_0__inst_mult_16_59  = CARRY(( (din_a[96] & din_b[96]) ) + ( Xd_0__inst_mult_22_97  ) + ( Xd_0__inst_mult_22_96  ))
// Xd_0__inst_mult_16_60  = SHARE((din_b[96] & din_a[97]))

	.dataa(!din_a[96]),
	.datab(!din_b[96]),
	.datac(!din_a[97]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_96 ),
	.sharein(Xd_0__inst_mult_22_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_58 ),
	.cout(Xd_0__inst_mult_16_59 ),
	.shareout(Xd_0__inst_mult_16_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_22 (
// Equation(s):
// Xd_0__inst_mult_17_67  = SUM(( (din_a[102] & din_b[102]) ) + ( Xd_0__inst_i17_119  ) + ( Xd_0__inst_i17_118  ))
// Xd_0__inst_mult_17_68  = CARRY(( (din_a[102] & din_b[102]) ) + ( Xd_0__inst_i17_119  ) + ( Xd_0__inst_i17_118  ))
// Xd_0__inst_mult_17_69  = SHARE((din_b[102] & din_a[103]))

	.dataa(!din_a[102]),
	.datab(!din_b[102]),
	.datac(!din_a[103]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_118 ),
	.sharein(Xd_0__inst_i17_119 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_67 ),
	.cout(Xd_0__inst_mult_17_68 ),
	.shareout(Xd_0__inst_mult_17_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_21 (
// Equation(s):
// Xd_0__inst_i17_21_sumout  = SUM(( !din_a[101] $ (!din_b[101]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_22  = CARRY(( !din_a[101] $ (!din_b[101]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_23  = SHARE(GND)

	.dataa(!din_a[101]),
	.datab(!din_b[101]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_21_sumout ),
	.cout(Xd_0__inst_i17_22 ),
	.shareout(Xd_0__inst_i17_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_20 (
// Equation(s):
// Xd_0__inst_mult_14_58  = SUM(( (din_a[84] & din_b[84]) ) + ( Xd_0__inst_mult_15_85  ) + ( Xd_0__inst_mult_15_84  ))
// Xd_0__inst_mult_14_59  = CARRY(( (din_a[84] & din_b[84]) ) + ( Xd_0__inst_mult_15_85  ) + ( Xd_0__inst_mult_15_84  ))
// Xd_0__inst_mult_14_60  = SHARE((din_b[84] & din_a[85]))

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(!din_a[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_84 ),
	.sharein(Xd_0__inst_mult_15_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_58 ),
	.cout(Xd_0__inst_mult_14_59 ),
	.shareout(Xd_0__inst_mult_14_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_22 (
// Equation(s):
// Xd_0__inst_mult_15_67  = SUM(( (din_a[90] & din_b[90]) ) + ( Xd_0__inst_i17_95  ) + ( Xd_0__inst_i17_94  ))
// Xd_0__inst_mult_15_68  = CARRY(( (din_a[90] & din_b[90]) ) + ( Xd_0__inst_i17_95  ) + ( Xd_0__inst_i17_94  ))
// Xd_0__inst_mult_15_69  = SHARE((din_b[90] & din_a[91]))

	.dataa(!din_a[90]),
	.datab(!din_b[90]),
	.datac(!din_a[91]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_94 ),
	.sharein(Xd_0__inst_i17_95 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_67 ),
	.cout(Xd_0__inst_mult_15_68 ),
	.shareout(Xd_0__inst_mult_15_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_25 (
// Equation(s):
// Xd_0__inst_i17_25_sumout  = SUM(( !din_a[89] $ (!din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_26  = CARRY(( !din_a[89] $ (!din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_27  = SHARE(GND)

	.dataa(!din_a[89]),
	.datab(!din_b[89]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_25_sumout ),
	.cout(Xd_0__inst_i17_26 ),
	.shareout(Xd_0__inst_i17_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_29 (
// Equation(s):
// Xd_0__inst_i17_29_sumout  = SUM(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i17_27  ) + ( Xd_0__inst_i17_26  ))
// Xd_0__inst_i17_30  = CARRY(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i17_27  ) + ( Xd_0__inst_i17_26  ))
// Xd_0__inst_i17_31  = SHARE(GND)

	.dataa(!din_a[95]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_26 ),
	.sharein(Xd_0__inst_i17_27 ),
	.combout(),
	.sumout(Xd_0__inst_i17_29_sumout ),
	.cout(Xd_0__inst_i17_30 ),
	.shareout(Xd_0__inst_i17_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_20 (
// Equation(s):
// Xd_0__inst_mult_12_58  = SUM(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_59  = CARRY(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_60  = SHARE((din_b[72] & din_a[73]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_a[73]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_12_58 ),
	.cout(Xd_0__inst_mult_12_59 ),
	.shareout(Xd_0__inst_mult_12_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_22 (
// Equation(s):
// Xd_0__inst_mult_13_67  = SUM(( (din_a[78] & din_b[78]) ) + ( Xd_0__inst_mult_29_93  ) + ( Xd_0__inst_mult_29_92  ))
// Xd_0__inst_mult_13_68  = CARRY(( (din_a[78] & din_b[78]) ) + ( Xd_0__inst_mult_29_93  ) + ( Xd_0__inst_mult_29_92  ))
// Xd_0__inst_mult_13_69  = SHARE((din_b[78] & din_a[79]))

	.dataa(!din_a[78]),
	.datab(!din_b[78]),
	.datac(!din_a[79]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_92 ),
	.sharein(Xd_0__inst_mult_29_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_67 ),
	.cout(Xd_0__inst_mult_13_68 ),
	.shareout(Xd_0__inst_mult_13_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_33 (
// Equation(s):
// Xd_0__inst_i17_33_sumout  = SUM(( !din_a[77] $ (!din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_34  = CARRY(( !din_a[77] $ (!din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_35  = SHARE(GND)

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_33_sumout ),
	.cout(Xd_0__inst_i17_34 ),
	.shareout(Xd_0__inst_i17_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_37 (
// Equation(s):
// Xd_0__inst_i17_37_sumout  = SUM(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i17_35  ) + ( Xd_0__inst_i17_34  ))
// Xd_0__inst_i17_38  = CARRY(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i17_35  ) + ( Xd_0__inst_i17_34  ))
// Xd_0__inst_i17_39  = SHARE(GND)

	.dataa(!din_a[83]),
	.datab(!din_b[83]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_34 ),
	.sharein(Xd_0__inst_i17_35 ),
	.combout(),
	.sumout(Xd_0__inst_i17_37_sumout ),
	.cout(Xd_0__inst_i17_38 ),
	.shareout(Xd_0__inst_i17_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_23 (
// Equation(s):
// Xd_0__inst_mult_29_71  = SUM(( (!din_a[178] & (((din_a[177] & din_b[175])))) # (din_a[178] & (!din_b[174] $ (((!din_a[177]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_29_97  ) + ( Xd_0__inst_mult_29_96  ))
// Xd_0__inst_mult_29_72  = CARRY(( (!din_a[178] & (((din_a[177] & din_b[175])))) # (din_a[178] & (!din_b[174] $ (((!din_a[177]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_29_97  ) + ( Xd_0__inst_mult_29_96  ))
// Xd_0__inst_mult_29_73  = SHARE((din_a[178] & (din_b[174] & (din_a[177] & din_b[175]))))

	.dataa(!din_a[178]),
	.datab(!din_b[174]),
	.datac(!din_a[177]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_96 ),
	.sharein(Xd_0__inst_mult_29_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_71 ),
	.cout(Xd_0__inst_mult_29_72 ),
	.shareout(Xd_0__inst_mult_29_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_20 (
// Equation(s):
// Xd_0__inst_mult_10_58  = SUM(( (din_a[60] & din_b[60]) ) + ( Xd_0__inst_mult_11_93  ) + ( Xd_0__inst_mult_11_92  ))
// Xd_0__inst_mult_10_59  = CARRY(( (din_a[60] & din_b[60]) ) + ( Xd_0__inst_mult_11_93  ) + ( Xd_0__inst_mult_11_92  ))
// Xd_0__inst_mult_10_60  = SHARE((din_b[60] & din_a[61]))

	.dataa(!din_a[60]),
	.datab(!din_b[60]),
	.datac(!din_a[61]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_92 ),
	.sharein(Xd_0__inst_mult_11_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_58 ),
	.cout(Xd_0__inst_mult_10_59 ),
	.shareout(Xd_0__inst_mult_10_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_23 (
// Equation(s):
// Xd_0__inst_mult_11_71  = SUM(( (din_a[66] & din_b[66]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_72  = CARRY(( (din_a[66] & din_b[66]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_73  = SHARE((din_b[66] & din_a[67]))

	.dataa(!din_a[66]),
	.datab(!din_b[66]),
	.datac(!din_a[67]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_11_71 ),
	.cout(Xd_0__inst_mult_11_72 ),
	.shareout(Xd_0__inst_mult_11_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_41 (
// Equation(s):
// Xd_0__inst_i17_41_sumout  = SUM(( !din_a[65] $ (!din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_42  = CARRY(( !din_a[65] $ (!din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_43  = SHARE(GND)

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_41_sumout ),
	.cout(Xd_0__inst_i17_42 ),
	.shareout(Xd_0__inst_i17_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_20 (
// Equation(s):
// Xd_0__inst_mult_8_58  = SUM(( (din_a[48] & din_b[48]) ) + ( Xd_0__inst_i17_31  ) + ( Xd_0__inst_i17_30  ))
// Xd_0__inst_mult_8_59  = CARRY(( (din_a[48] & din_b[48]) ) + ( Xd_0__inst_i17_31  ) + ( Xd_0__inst_i17_30  ))
// Xd_0__inst_mult_8_60  = SHARE((din_b[48] & din_a[49]))

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(!din_a[49]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_30 ),
	.sharein(Xd_0__inst_i17_31 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_58 ),
	.cout(Xd_0__inst_mult_8_59 ),
	.shareout(Xd_0__inst_mult_8_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_22 (
// Equation(s):
// Xd_0__inst_mult_9_67  = SUM(( (din_a[54] & din_b[54]) ) + ( Xd_0__inst_i17_63  ) + ( Xd_0__inst_i17_62  ))
// Xd_0__inst_mult_9_68  = CARRY(( (din_a[54] & din_b[54]) ) + ( Xd_0__inst_i17_63  ) + ( Xd_0__inst_i17_62  ))
// Xd_0__inst_mult_9_69  = SHARE((din_b[54] & din_a[55]))

	.dataa(!din_a[54]),
	.datab(!din_b[54]),
	.datac(!din_a[55]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_62 ),
	.sharein(Xd_0__inst_i17_63 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_67 ),
	.cout(Xd_0__inst_mult_9_68 ),
	.shareout(Xd_0__inst_mult_9_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_45 (
// Equation(s):
// Xd_0__inst_i17_45_sumout  = SUM(( !din_a[53] $ (!din_b[53]) ) + ( Xd_0__inst_i17_51  ) + ( Xd_0__inst_i17_50  ))
// Xd_0__inst_i17_46  = CARRY(( !din_a[53] $ (!din_b[53]) ) + ( Xd_0__inst_i17_51  ) + ( Xd_0__inst_i17_50  ))
// Xd_0__inst_i17_47  = SHARE(GND)

	.dataa(!din_a[53]),
	.datab(!din_b[53]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_50 ),
	.sharein(Xd_0__inst_i17_51 ),
	.combout(),
	.sumout(Xd_0__inst_i17_45_sumout ),
	.cout(Xd_0__inst_i17_46 ),
	.shareout(Xd_0__inst_i17_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_49 (
// Equation(s):
// Xd_0__inst_i17_49_sumout  = SUM(( !din_a[59] $ (!din_b[59]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_50  = CARRY(( !din_a[59] $ (!din_b[59]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_51  = SHARE(GND)

	.dataa(!din_a[59]),
	.datab(!din_b[59]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_49_sumout ),
	.cout(Xd_0__inst_i17_50 ),
	.shareout(Xd_0__inst_i17_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_20 (
// Equation(s):
// Xd_0__inst_mult_6_57  = SUM(( (din_a[36] & din_b[36]) ) + ( Xd_0__inst_mult_9_85  ) + ( Xd_0__inst_mult_9_84  ))
// Xd_0__inst_mult_6_58  = CARRY(( (din_a[36] & din_b[36]) ) + ( Xd_0__inst_mult_9_85  ) + ( Xd_0__inst_mult_9_84  ))
// Xd_0__inst_mult_6_59  = SHARE((din_b[36] & din_a[37]))

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(!din_a[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_84 ),
	.sharein(Xd_0__inst_mult_9_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_57 ),
	.cout(Xd_0__inst_mult_6_58 ),
	.shareout(Xd_0__inst_mult_6_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_22 (
// Equation(s):
// Xd_0__inst_mult_7_66  = SUM(( (din_a[42] & din_b[42]) ) + ( Xd_0__inst_i17_55  ) + ( Xd_0__inst_i17_54  ))
// Xd_0__inst_mult_7_67  = CARRY(( (din_a[42] & din_b[42]) ) + ( Xd_0__inst_i17_55  ) + ( Xd_0__inst_i17_54  ))
// Xd_0__inst_mult_7_68  = SHARE((din_b[42] & din_a[43]))

	.dataa(!din_a[42]),
	.datab(!din_b[42]),
	.datac(!din_a[43]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_54 ),
	.sharein(Xd_0__inst_i17_55 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_66 ),
	.cout(Xd_0__inst_mult_7_67 ),
	.shareout(Xd_0__inst_mult_7_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_53 (
// Equation(s):
// Xd_0__inst_i17_53_sumout  = SUM(( !din_a[41] $ (!din_b[41]) ) + ( Xd_0__inst_i17_59  ) + ( Xd_0__inst_i17_58  ))
// Xd_0__inst_i17_54  = CARRY(( !din_a[41] $ (!din_b[41]) ) + ( Xd_0__inst_i17_59  ) + ( Xd_0__inst_i17_58  ))
// Xd_0__inst_i17_55  = SHARE(GND)

	.dataa(!din_a[41]),
	.datab(!din_b[41]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_58 ),
	.sharein(Xd_0__inst_i17_59 ),
	.combout(),
	.sumout(Xd_0__inst_i17_53_sumout ),
	.cout(Xd_0__inst_i17_54 ),
	.shareout(Xd_0__inst_i17_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_57 (
// Equation(s):
// Xd_0__inst_i17_57_sumout  = SUM(( !din_a[47] $ (!din_b[47]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_58  = CARRY(( !din_a[47] $ (!din_b[47]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_59  = SHARE(GND)

	.dataa(!din_a[47]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_57_sumout ),
	.cout(Xd_0__inst_i17_58 ),
	.shareout(Xd_0__inst_i17_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_27 (
// Equation(s):
// Xd_0__inst_mult_31_87  = SUM(( (!din_a[190] & (((din_a[189] & din_b[187])))) # (din_a[190] & (!din_b[186] $ (((!din_a[189]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_31_117  ) + ( Xd_0__inst_mult_31_116  ))
// Xd_0__inst_mult_31_88  = CARRY(( (!din_a[190] & (((din_a[189] & din_b[187])))) # (din_a[190] & (!din_b[186] $ (((!din_a[189]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_31_117  ) + ( Xd_0__inst_mult_31_116  ))
// Xd_0__inst_mult_31_89  = SHARE((din_a[190] & (din_b[186] & (din_a[189] & din_b[187]))))

	.dataa(!din_a[190]),
	.datab(!din_b[186]),
	.datac(!din_a[189]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_116 ),
	.sharein(Xd_0__inst_mult_31_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_87 ),
	.cout(Xd_0__inst_mult_31_88 ),
	.shareout(Xd_0__inst_mult_31_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_20 (
// Equation(s):
// Xd_0__inst_mult_4_57  = SUM(( (din_a[24] & din_b[24]) ) + ( Xd_0__inst_mult_8_76  ) + ( Xd_0__inst_mult_8_75  ))
// Xd_0__inst_mult_4_58  = CARRY(( (din_a[24] & din_b[24]) ) + ( Xd_0__inst_mult_8_76  ) + ( Xd_0__inst_mult_8_75  ))
// Xd_0__inst_mult_4_59  = SHARE((din_b[24] & din_a[25]))

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(!din_a[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_75 ),
	.sharein(Xd_0__inst_mult_8_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_57 ),
	.cout(Xd_0__inst_mult_4_58 ),
	.shareout(Xd_0__inst_mult_4_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_22 (
// Equation(s):
// Xd_0__inst_mult_5_66  = SUM(( (din_a[30] & din_b[30]) ) + ( Xd_0__inst_mult_7_84  ) + ( Xd_0__inst_mult_7_83  ))
// Xd_0__inst_mult_5_67  = CARRY(( (din_a[30] & din_b[30]) ) + ( Xd_0__inst_mult_7_84  ) + ( Xd_0__inst_mult_7_83  ))
// Xd_0__inst_mult_5_68  = SHARE((din_b[30] & din_a[31]))

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(!din_a[31]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_83 ),
	.sharein(Xd_0__inst_mult_7_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_66 ),
	.cout(Xd_0__inst_mult_5_67 ),
	.shareout(Xd_0__inst_mult_5_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_61 (
// Equation(s):
// Xd_0__inst_i17_61_sumout  = SUM(( !din_a[29] $ (!din_b[29]) ) + ( Xd_0__inst_i17_67  ) + ( Xd_0__inst_i17_66  ))
// Xd_0__inst_i17_62  = CARRY(( !din_a[29] $ (!din_b[29]) ) + ( Xd_0__inst_i17_67  ) + ( Xd_0__inst_i17_66  ))
// Xd_0__inst_i17_63  = SHARE(GND)

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_66 ),
	.sharein(Xd_0__inst_i17_67 ),
	.combout(),
	.sumout(Xd_0__inst_i17_61_sumout ),
	.cout(Xd_0__inst_i17_62 ),
	.shareout(Xd_0__inst_i17_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_65 (
// Equation(s):
// Xd_0__inst_i17_65_sumout  = SUM(( !din_a[35] $ (!din_b[35]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_66  = CARRY(( !din_a[35] $ (!din_b[35]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_67  = SHARE(GND)

	.dataa(!din_a[35]),
	.datab(!din_b[35]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_65_sumout ),
	.cout(Xd_0__inst_i17_66 ),
	.shareout(Xd_0__inst_i17_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_22 (
// Equation(s):
// Xd_0__inst_mult_2_66  = SUM(( (din_a[12] & din_b[12]) ) + ( Xd_0__inst_i17_39  ) + ( Xd_0__inst_i17_38  ))
// Xd_0__inst_mult_2_67  = CARRY(( (din_a[12] & din_b[12]) ) + ( Xd_0__inst_i17_39  ) + ( Xd_0__inst_i17_38  ))
// Xd_0__inst_mult_2_68  = SHARE((din_b[12] & din_a[13]))

	.dataa(!din_a[12]),
	.datab(!din_b[12]),
	.datac(!din_a[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_38 ),
	.sharein(Xd_0__inst_i17_39 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_66 ),
	.cout(Xd_0__inst_mult_2_67 ),
	.shareout(Xd_0__inst_mult_2_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_22 (
// Equation(s):
// Xd_0__inst_mult_3_66  = SUM(( (din_a[18] & din_b[18]) ) + ( Xd_0__inst_mult_2_84  ) + ( Xd_0__inst_mult_2_83  ))
// Xd_0__inst_mult_3_67  = CARRY(( (din_a[18] & din_b[18]) ) + ( Xd_0__inst_mult_2_84  ) + ( Xd_0__inst_mult_2_83  ))
// Xd_0__inst_mult_3_68  = SHARE((din_b[18] & din_a[19]))

	.dataa(!din_a[18]),
	.datab(!din_b[18]),
	.datac(!din_a[19]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_83 ),
	.sharein(Xd_0__inst_mult_2_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_66 ),
	.cout(Xd_0__inst_mult_3_67 ),
	.shareout(Xd_0__inst_mult_3_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_69 (
// Equation(s):
// Xd_0__inst_i17_69_sumout  = SUM(( !din_a[17] $ (!din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_70  = CARRY(( !din_a[17] $ (!din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_71  = SHARE(GND)

	.dataa(!din_a[17]),
	.datab(!din_b[17]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_69_sumout ),
	.cout(Xd_0__inst_i17_70 ),
	.shareout(Xd_0__inst_i17_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_73 (
// Equation(s):
// Xd_0__inst_i17_73_sumout  = SUM(( !din_a[23] $ (!din_b[23]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_74  = CARRY(( !din_a[23] $ (!din_b[23]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_75  = SHARE(GND)

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_73_sumout ),
	.cout(Xd_0__inst_i17_74 ),
	.shareout(Xd_0__inst_i17_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_22 (
// Equation(s):
// Xd_0__inst_mult_0_66  = SUM(( (din_a[0] & din_b[0]) ) + ( Xd_0__inst_i17_47  ) + ( Xd_0__inst_i17_46  ))
// Xd_0__inst_mult_0_67  = CARRY(( (din_a[0] & din_b[0]) ) + ( Xd_0__inst_i17_47  ) + ( Xd_0__inst_i17_46  ))
// Xd_0__inst_mult_0_68  = SHARE((din_b[0] & din_a[1]))

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_a[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_46 ),
	.sharein(Xd_0__inst_i17_47 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_66 ),
	.cout(Xd_0__inst_mult_0_67 ),
	.shareout(Xd_0__inst_mult_0_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_22 (
// Equation(s):
// Xd_0__inst_mult_1_66  = SUM(( (din_a[6] & din_b[6]) ) + ( Xd_0__inst_mult_0_84  ) + ( Xd_0__inst_mult_0_83  ))
// Xd_0__inst_mult_1_67  = CARRY(( (din_a[6] & din_b[6]) ) + ( Xd_0__inst_mult_0_84  ) + ( Xd_0__inst_mult_0_83  ))
// Xd_0__inst_mult_1_68  = SHARE((din_b[6] & din_a[7]))

	.dataa(!din_a[6]),
	.datab(!din_b[6]),
	.datac(!din_a[7]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_83 ),
	.sharein(Xd_0__inst_mult_0_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_66 ),
	.cout(Xd_0__inst_mult_1_67 ),
	.shareout(Xd_0__inst_mult_1_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_77 (
// Equation(s):
// Xd_0__inst_i17_77_sumout  = SUM(( !din_a[5] $ (!din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_78  = CARRY(( !din_a[5] $ (!din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_79  = SHARE(GND)

	.dataa(!din_a[5]),
	.datab(!din_b[5]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_77_sumout ),
	.cout(Xd_0__inst_i17_78 ),
	.shareout(Xd_0__inst_i17_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_81 (
// Equation(s):
// Xd_0__inst_i17_81_sumout  = SUM(( !din_a[11] $ (!din_b[11]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_82  = CARRY(( !din_a[11] $ (!din_b[11]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_83  = SHARE(GND)

	.dataa(!din_a[11]),
	.datab(!din_b[11]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_81_sumout ),
	.cout(Xd_0__inst_i17_82 ),
	.shareout(Xd_0__inst_i17_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_24 (
// Equation(s):
// Xd_0__inst_mult_11_75  = SUM(( (!din_a[70] & (((din_a[69] & din_b[67])))) # (din_a[70] & (!din_b[66] $ (((!din_a[69]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_11_97  ) + ( Xd_0__inst_mult_11_96  ))
// Xd_0__inst_mult_11_76  = CARRY(( (!din_a[70] & (((din_a[69] & din_b[67])))) # (din_a[70] & (!din_b[66] $ (((!din_a[69]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_11_97  ) + ( Xd_0__inst_mult_11_96  ))
// Xd_0__inst_mult_11_77  = SHARE((din_a[70] & (din_b[66] & (din_a[69] & din_b[67]))))

	.dataa(!din_a[70]),
	.datab(!din_b[66]),
	.datac(!din_a[69]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_96 ),
	.sharein(Xd_0__inst_mult_11_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_75 ),
	.cout(Xd_0__inst_mult_11_76 ),
	.shareout(Xd_0__inst_mult_11_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_25 (
// Equation(s):
// Xd_0__inst_mult_28_79  = SUM(( (din_a[168] & din_b[168]) ) + ( Xd_0__inst_mult_21_85  ) + ( Xd_0__inst_mult_21_84  ))
// Xd_0__inst_mult_28_80  = CARRY(( (din_a[168] & din_b[168]) ) + ( Xd_0__inst_mult_21_85  ) + ( Xd_0__inst_mult_21_84  ))
// Xd_0__inst_mult_28_81  = SHARE((din_b[168] & din_a[169]))

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(!din_a[169]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_84 ),
	.sharein(Xd_0__inst_mult_21_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_79 ),
	.cout(Xd_0__inst_mult_28_80 ),
	.shareout(Xd_0__inst_mult_28_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_24 (
// Equation(s):
// Xd_0__inst_mult_29_75  = SUM(( (din_a[174] & din_b[174]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_29_76  = CARRY(( (din_a[174] & din_b[174]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_29_77  = SHARE((din_b[174] & din_a[175]))

	.dataa(!din_a[174]),
	.datab(!din_b[174]),
	.datac(!din_a[175]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_29_75 ),
	.cout(Xd_0__inst_mult_29_76 ),
	.shareout(Xd_0__inst_mult_29_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_85 (
// Equation(s):
// Xd_0__inst_i17_85_sumout  = SUM(( !din_a[173] $ (!din_b[173]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_86  = CARRY(( !din_a[173] $ (!din_b[173]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_87  = SHARE(GND)

	.dataa(!din_a[173]),
	.datab(!din_b[173]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_85_sumout ),
	.cout(Xd_0__inst_i17_86 ),
	.shareout(Xd_0__inst_i17_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_89 (
// Equation(s):
// Xd_0__inst_i17_89_sumout  = SUM(( !din_a[179] $ (!din_b[179]) ) + ( Xd_0__inst_i17_87  ) + ( Xd_0__inst_i17_86  ))
// Xd_0__inst_i17_90  = CARRY(( !din_a[179] $ (!din_b[179]) ) + ( Xd_0__inst_i17_87  ) + ( Xd_0__inst_i17_86  ))
// Xd_0__inst_i17_91  = SHARE(GND)

	.dataa(!din_a[179]),
	.datab(!din_b[179]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_86 ),
	.sharein(Xd_0__inst_i17_87 ),
	.combout(),
	.sumout(Xd_0__inst_i17_89_sumout ),
	.cout(Xd_0__inst_i17_90 ),
	.shareout(Xd_0__inst_i17_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_25 (
// Equation(s):
// Xd_0__inst_mult_26_79  = SUM(( (din_a[156] & din_b[156]) ) + ( Xd_0__inst_i17_19  ) + ( Xd_0__inst_i17_18  ))
// Xd_0__inst_mult_26_80  = CARRY(( (din_a[156] & din_b[156]) ) + ( Xd_0__inst_i17_19  ) + ( Xd_0__inst_i17_18  ))
// Xd_0__inst_mult_26_81  = SHARE((din_b[156] & din_a[157]))

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(!din_a[157]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_18 ),
	.sharein(Xd_0__inst_i17_19 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_79 ),
	.cout(Xd_0__inst_mult_26_80 ),
	.shareout(Xd_0__inst_mult_26_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_23 (
// Equation(s):
// Xd_0__inst_mult_27_71  = SUM(( (din_a[162] & din_b[162]) ) + ( Xd_0__inst_mult_26_97  ) + ( Xd_0__inst_mult_26_96  ))
// Xd_0__inst_mult_27_72  = CARRY(( (din_a[162] & din_b[162]) ) + ( Xd_0__inst_mult_26_97  ) + ( Xd_0__inst_mult_26_96  ))
// Xd_0__inst_mult_27_73  = SHARE((din_b[162] & din_a[163]))

	.dataa(!din_a[162]),
	.datab(!din_b[162]),
	.datac(!din_a[163]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_96 ),
	.sharein(Xd_0__inst_mult_26_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_71 ),
	.cout(Xd_0__inst_mult_27_72 ),
	.shareout(Xd_0__inst_mult_27_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_93 (
// Equation(s):
// Xd_0__inst_i17_93_sumout  = SUM(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i17_43  ) + ( Xd_0__inst_i17_42  ))
// Xd_0__inst_i17_94  = CARRY(( !din_a[167] $ (!din_b[167]) ) + ( Xd_0__inst_i17_43  ) + ( Xd_0__inst_i17_42  ))
// Xd_0__inst_i17_95  = SHARE(GND)

	.dataa(!din_a[167]),
	.datab(!din_b[167]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_42 ),
	.sharein(Xd_0__inst_i17_43 ),
	.combout(),
	.sumout(Xd_0__inst_i17_93_sumout ),
	.cout(Xd_0__inst_i17_94 ),
	.shareout(Xd_0__inst_i17_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_25 (
// Equation(s):
// Xd_0__inst_mult_24_79  = SUM(( (din_a[144] & din_b[144]) ) + ( Xd_0__inst_i17_103  ) + ( Xd_0__inst_i17_102  ))
// Xd_0__inst_mult_24_80  = CARRY(( (din_a[144] & din_b[144]) ) + ( Xd_0__inst_i17_103  ) + ( Xd_0__inst_i17_102  ))
// Xd_0__inst_mult_24_81  = SHARE((din_b[144] & din_a[145]))

	.dataa(!din_a[144]),
	.datab(!din_b[144]),
	.datac(!din_a[145]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_102 ),
	.sharein(Xd_0__inst_i17_103 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_79 ),
	.cout(Xd_0__inst_mult_24_80 ),
	.shareout(Xd_0__inst_mult_24_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_23 (
// Equation(s):
// Xd_0__inst_mult_25_71  = SUM(( (din_a[150] & din_b[150]) ) + ( Xd_0__inst_mult_24_97  ) + ( Xd_0__inst_mult_24_96  ))
// Xd_0__inst_mult_25_72  = CARRY(( (din_a[150] & din_b[150]) ) + ( Xd_0__inst_mult_24_97  ) + ( Xd_0__inst_mult_24_96  ))
// Xd_0__inst_mult_25_73  = SHARE((din_b[150] & din_a[151]))

	.dataa(!din_a[150]),
	.datab(!din_b[150]),
	.datac(!din_a[151]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_96 ),
	.sharein(Xd_0__inst_mult_24_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_71 ),
	.cout(Xd_0__inst_mult_25_72 ),
	.shareout(Xd_0__inst_mult_25_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_97 (
// Equation(s):
// Xd_0__inst_i17_97_sumout  = SUM(( !din_a[149] $ (!din_b[149]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_98  = CARRY(( !din_a[149] $ (!din_b[149]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_99  = SHARE(GND)

	.dataa(!din_a[149]),
	.datab(!din_b[149]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_97_sumout ),
	.cout(Xd_0__inst_i17_98 ),
	.shareout(Xd_0__inst_i17_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_101 (
// Equation(s):
// Xd_0__inst_i17_101_sumout  = SUM(( !din_a[155] $ (!din_b[155]) ) + ( Xd_0__inst_i17_99  ) + ( Xd_0__inst_i17_98  ))
// Xd_0__inst_i17_102  = CARRY(( !din_a[155] $ (!din_b[155]) ) + ( Xd_0__inst_i17_99  ) + ( Xd_0__inst_i17_98  ))
// Xd_0__inst_i17_103  = SHARE(GND)

	.dataa(!din_a[155]),
	.datab(!din_b[155]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_98 ),
	.sharein(Xd_0__inst_i17_99 ),
	.combout(),
	.sumout(Xd_0__inst_i17_101_sumout ),
	.cout(Xd_0__inst_i17_102 ),
	.shareout(Xd_0__inst_i17_103 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_24 (
// Equation(s):
// Xd_0__inst_mult_25_75  = SUM(( (!din_a[154] & (((din_a[153] & din_b[151])))) # (din_a[154] & (!din_b[150] $ (((!din_a[153]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_25_93  ) + ( Xd_0__inst_mult_25_92  ))
// Xd_0__inst_mult_25_76  = CARRY(( (!din_a[154] & (((din_a[153] & din_b[151])))) # (din_a[154] & (!din_b[150] $ (((!din_a[153]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_25_93  ) + ( Xd_0__inst_mult_25_92  ))
// Xd_0__inst_mult_25_77  = SHARE((din_a[154] & (din_b[150] & (din_a[153] & din_b[151]))))

	.dataa(!din_a[154]),
	.datab(!din_b[150]),
	.datac(!din_a[153]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_92 ),
	.sharein(Xd_0__inst_mult_25_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_75 ),
	.cout(Xd_0__inst_mult_25_76 ),
	.shareout(Xd_0__inst_mult_25_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_25 (
// Equation(s):
// Xd_0__inst_mult_22_79  = SUM(( (din_a[132] & din_b[132]) ) + ( Xd_0__inst_i17_111  ) + ( Xd_0__inst_i17_110  ))
// Xd_0__inst_mult_22_80  = CARRY(( (din_a[132] & din_b[132]) ) + ( Xd_0__inst_i17_111  ) + ( Xd_0__inst_i17_110  ))
// Xd_0__inst_mult_22_81  = SHARE((din_b[132] & din_a[133]))

	.dataa(!din_a[132]),
	.datab(!din_b[132]),
	.datac(!din_a[133]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_110 ),
	.sharein(Xd_0__inst_i17_111 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_79 ),
	.cout(Xd_0__inst_mult_22_80 ),
	.shareout(Xd_0__inst_mult_22_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_25 (
// Equation(s):
// Xd_0__inst_mult_23_79  = SUM(( (din_a[138] & din_b[138]) ) + ( Xd_0__inst_mult_19_97  ) + ( Xd_0__inst_mult_19_96  ))
// Xd_0__inst_mult_23_80  = CARRY(( (din_a[138] & din_b[138]) ) + ( Xd_0__inst_mult_19_97  ) + ( Xd_0__inst_mult_19_96  ))
// Xd_0__inst_mult_23_81  = SHARE((din_b[138] & din_a[139]))

	.dataa(!din_a[138]),
	.datab(!din_b[138]),
	.datac(!din_a[139]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_96 ),
	.sharein(Xd_0__inst_mult_19_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_79 ),
	.cout(Xd_0__inst_mult_23_80 ),
	.shareout(Xd_0__inst_mult_23_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_105 (
// Equation(s):
// Xd_0__inst_i17_105_sumout  = SUM(( !din_a[137] $ (!din_b[137]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_106  = CARRY(( !din_a[137] $ (!din_b[137]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_107  = SHARE(GND)

	.dataa(!din_a[137]),
	.datab(!din_b[137]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_105_sumout ),
	.cout(Xd_0__inst_i17_106 ),
	.shareout(Xd_0__inst_i17_107 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_109 (
// Equation(s):
// Xd_0__inst_i17_109_sumout  = SUM(( !din_a[143] $ (!din_b[143]) ) + ( Xd_0__inst_i17_107  ) + ( Xd_0__inst_i17_106  ))
// Xd_0__inst_i17_110  = CARRY(( !din_a[143] $ (!din_b[143]) ) + ( Xd_0__inst_i17_107  ) + ( Xd_0__inst_i17_106  ))
// Xd_0__inst_i17_111  = SHARE(GND)

	.dataa(!din_a[143]),
	.datab(!din_b[143]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_106 ),
	.sharein(Xd_0__inst_i17_107 ),
	.combout(),
	.sumout(Xd_0__inst_i17_109_sumout ),
	.cout(Xd_0__inst_i17_110 ),
	.shareout(Xd_0__inst_i17_111 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_25 (
// Equation(s):
// Xd_0__inst_mult_20_79  = SUM(( (din_a[120] & din_b[120]) ) + ( Xd_0__inst_mult_17_85  ) + ( Xd_0__inst_mult_17_84  ))
// Xd_0__inst_mult_20_80  = CARRY(( (din_a[120] & din_b[120]) ) + ( Xd_0__inst_mult_17_85  ) + ( Xd_0__inst_mult_17_84  ))
// Xd_0__inst_mult_20_81  = SHARE((din_b[120] & din_a[121]))

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(!din_a[121]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_84 ),
	.sharein(Xd_0__inst_mult_17_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_79 ),
	.cout(Xd_0__inst_mult_20_80 ),
	.shareout(Xd_0__inst_mult_20_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_22 (
// Equation(s):
// Xd_0__inst_mult_21_67  = SUM(( (din_a[126] & din_b[126]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_21_68  = CARRY(( (din_a[126] & din_b[126]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_21_69  = SHARE((din_b[126] & din_a[127]))

	.dataa(!din_a[126]),
	.datab(!din_b[126]),
	.datac(!din_a[127]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_21_67 ),
	.cout(Xd_0__inst_mult_21_68 ),
	.shareout(Xd_0__inst_mult_21_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_113 (
// Equation(s):
// Xd_0__inst_i17_113_sumout  = SUM(( !din_a[125] $ (!din_b[125]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_114  = CARRY(( !din_a[125] $ (!din_b[125]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_115  = SHARE(GND)

	.dataa(!din_a[125]),
	.datab(!din_b[125]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_113_sumout ),
	.cout(Xd_0__inst_i17_114 ),
	.shareout(Xd_0__inst_i17_115 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_117 (
// Equation(s):
// Xd_0__inst_i17_117_sumout  = SUM(( !din_a[131] $ (!din_b[131]) ) + ( Xd_0__inst_i17_115  ) + ( Xd_0__inst_i17_114  ))
// Xd_0__inst_i17_118  = CARRY(( !din_a[131] $ (!din_b[131]) ) + ( Xd_0__inst_i17_115  ) + ( Xd_0__inst_i17_114  ))
// Xd_0__inst_i17_119  = SHARE(GND)

	.dataa(!din_a[131]),
	.datab(!din_b[131]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_114 ),
	.sharein(Xd_0__inst_i17_115 ),
	.combout(),
	.sumout(Xd_0__inst_i17_117_sumout ),
	.cout(Xd_0__inst_i17_118 ),
	.shareout(Xd_0__inst_i17_119 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_20 (
// Equation(s):
// Xd_0__inst_mult_18_58  = SUM(( (din_a[108] & din_b[108]) ) + ( Xd_0__inst_mult_12_76  ) + ( Xd_0__inst_mult_12_75  ))
// Xd_0__inst_mult_18_59  = CARRY(( (din_a[108] & din_b[108]) ) + ( Xd_0__inst_mult_12_76  ) + ( Xd_0__inst_mult_12_75  ))
// Xd_0__inst_mult_18_60  = SHARE((din_b[108] & din_a[109]))

	.dataa(!din_a[108]),
	.datab(!din_b[108]),
	.datac(!din_a[109]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_75 ),
	.sharein(Xd_0__inst_mult_12_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_58 ),
	.cout(Xd_0__inst_mult_18_59 ),
	.shareout(Xd_0__inst_mult_18_60 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_25 (
// Equation(s):
// Xd_0__inst_mult_19_79  = SUM(( (din_a[114] & din_b[114]) ) + ( Xd_0__inst_i17_91  ) + ( Xd_0__inst_i17_90  ))
// Xd_0__inst_mult_19_80  = CARRY(( (din_a[114] & din_b[114]) ) + ( Xd_0__inst_i17_91  ) + ( Xd_0__inst_i17_90  ))
// Xd_0__inst_mult_19_81  = SHARE((din_b[114] & din_a[115]))

	.dataa(!din_a[114]),
	.datab(!din_b[114]),
	.datac(!din_a[115]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_90 ),
	.sharein(Xd_0__inst_i17_91 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_79 ),
	.cout(Xd_0__inst_mult_19_80 ),
	.shareout(Xd_0__inst_mult_19_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_121 (
// Equation(s):
// Xd_0__inst_i17_121_sumout  = SUM(( !din_a[113] $ (!din_b[113]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_122  = CARRY(( !din_a[113] $ (!din_b[113]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_123  = SHARE(GND)

	.dataa(!din_a[113]),
	.datab(!din_b[113]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_121_sumout ),
	.cout(Xd_0__inst_i17_122 ),
	.shareout(Xd_0__inst_i17_123 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i17_125 (
// Equation(s):
// Xd_0__inst_i17_125_sumout  = SUM(( !din_a[119] $ (!din_b[119]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_126  = CARRY(( !din_a[119] $ (!din_b[119]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i17_127  = SHARE(GND)

	.dataa(!din_a[119]),
	.datab(!din_b[119]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i17_125_sumout ),
	.cout(Xd_0__inst_i17_126 ),
	.shareout(Xd_0__inst_i17_127 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_24 (
// Equation(s):
// Xd_0__inst_mult_27_75  = SUM(( (!din_a[166] & (((din_a[165] & din_b[163])))) # (din_a[166] & (!din_b[162] $ (((!din_a[165]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_27_93  ) + ( Xd_0__inst_mult_27_92  ))
// Xd_0__inst_mult_27_76  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[163])))) # (din_a[166] & (!din_b[162] $ (((!din_a[165]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_27_93  ) + ( Xd_0__inst_mult_27_92  ))
// Xd_0__inst_mult_27_77  = SHARE((din_a[166] & (din_b[162] & (din_a[165] & din_b[163]))))

	.dataa(!din_a[166]),
	.datab(!din_b[162]),
	.datac(!din_a[165]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_92 ),
	.sharein(Xd_0__inst_mult_27_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_75 ),
	.cout(Xd_0__inst_mult_27_76 ),
	.shareout(Xd_0__inst_mult_27_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_30_29 (
// Equation(s):
// Xd_0__inst_mult_30_95  = SUM(( GND ) + ( Xd_0__inst_mult_30_117  ) + ( Xd_0__inst_mult_30_116  ))
// Xd_0__inst_mult_30_96  = CARRY(( GND ) + ( Xd_0__inst_mult_30_117  ) + ( Xd_0__inst_mult_30_116  ))
// Xd_0__inst_mult_30_97  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_116 ),
	.sharein(Xd_0__inst_mult_30_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_95 ),
	.cout(Xd_0__inst_mult_30_96 ),
	.shareout(Xd_0__inst_mult_30_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_16_21 (
// Equation(s):
// Xd_0__inst_mult_16_62  = SUM(( (din_a[96] & din_b[97]) ) + ( Xd_0__inst_mult_16_60  ) + ( Xd_0__inst_mult_16_59  ))
// Xd_0__inst_mult_16_63  = CARRY(( (din_a[96] & din_b[97]) ) + ( Xd_0__inst_mult_16_60  ) + ( Xd_0__inst_mult_16_59  ))
// Xd_0__inst_mult_16_64  = SHARE((din_b[96] & din_a[98]))

	.dataa(!din_a[96]),
	.datab(!din_b[96]),
	.datac(!din_b[97]),
	.datad(!din_a[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_59 ),
	.sharein(Xd_0__inst_mult_16_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_62 ),
	.cout(Xd_0__inst_mult_16_63 ),
	.shareout(Xd_0__inst_mult_16_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_17_23 (
// Equation(s):
// Xd_0__inst_mult_17_71  = SUM(( (din_a[102] & din_b[103]) ) + ( Xd_0__inst_mult_17_69  ) + ( Xd_0__inst_mult_17_68  ))
// Xd_0__inst_mult_17_72  = CARRY(( (din_a[102] & din_b[103]) ) + ( Xd_0__inst_mult_17_69  ) + ( Xd_0__inst_mult_17_68  ))
// Xd_0__inst_mult_17_73  = SHARE((din_b[102] & din_a[104]))

	.dataa(!din_a[102]),
	.datab(!din_b[102]),
	.datac(!din_b[103]),
	.datad(!din_a[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_68 ),
	.sharein(Xd_0__inst_mult_17_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_71 ),
	.cout(Xd_0__inst_mult_17_72 ),
	.shareout(Xd_0__inst_mult_17_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_14_21 (
// Equation(s):
// Xd_0__inst_mult_14_62  = SUM(( (din_a[84] & din_b[85]) ) + ( Xd_0__inst_mult_14_60  ) + ( Xd_0__inst_mult_14_59  ))
// Xd_0__inst_mult_14_63  = CARRY(( (din_a[84] & din_b[85]) ) + ( Xd_0__inst_mult_14_60  ) + ( Xd_0__inst_mult_14_59  ))
// Xd_0__inst_mult_14_64  = SHARE((din_b[84] & din_a[86]))

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(!din_a[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_59 ),
	.sharein(Xd_0__inst_mult_14_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_62 ),
	.cout(Xd_0__inst_mult_14_63 ),
	.shareout(Xd_0__inst_mult_14_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_15_23 (
// Equation(s):
// Xd_0__inst_mult_15_71  = SUM(( (din_a[90] & din_b[91]) ) + ( Xd_0__inst_mult_15_69  ) + ( Xd_0__inst_mult_15_68  ))
// Xd_0__inst_mult_15_72  = CARRY(( (din_a[90] & din_b[91]) ) + ( Xd_0__inst_mult_15_69  ) + ( Xd_0__inst_mult_15_68  ))
// Xd_0__inst_mult_15_73  = SHARE((din_b[90] & din_a[92]))

	.dataa(!din_a[90]),
	.datab(!din_b[90]),
	.datac(!din_b[91]),
	.datad(!din_a[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_68 ),
	.sharein(Xd_0__inst_mult_15_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_71 ),
	.cout(Xd_0__inst_mult_15_72 ),
	.shareout(Xd_0__inst_mult_15_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_12_21 (
// Equation(s):
// Xd_0__inst_mult_12_62  = SUM(( (din_a[72] & din_b[73]) ) + ( Xd_0__inst_mult_12_60  ) + ( Xd_0__inst_mult_12_59  ))
// Xd_0__inst_mult_12_63  = CARRY(( (din_a[72] & din_b[73]) ) + ( Xd_0__inst_mult_12_60  ) + ( Xd_0__inst_mult_12_59  ))
// Xd_0__inst_mult_12_64  = SHARE((din_b[72] & din_a[74]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_b[73]),
	.datad(!din_a[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_59 ),
	.sharein(Xd_0__inst_mult_12_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_62 ),
	.cout(Xd_0__inst_mult_12_63 ),
	.shareout(Xd_0__inst_mult_12_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_13_23 (
// Equation(s):
// Xd_0__inst_mult_13_71  = SUM(( (din_a[78] & din_b[79]) ) + ( Xd_0__inst_mult_13_69  ) + ( Xd_0__inst_mult_13_68  ))
// Xd_0__inst_mult_13_72  = CARRY(( (din_a[78] & din_b[79]) ) + ( Xd_0__inst_mult_13_69  ) + ( Xd_0__inst_mult_13_68  ))
// Xd_0__inst_mult_13_73  = SHARE((din_b[78] & din_a[80]))

	.dataa(!din_a[78]),
	.datab(!din_b[78]),
	.datac(!din_b[79]),
	.datad(!din_a[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_68 ),
	.sharein(Xd_0__inst_mult_13_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_71 ),
	.cout(Xd_0__inst_mult_13_72 ),
	.shareout(Xd_0__inst_mult_13_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_10_21 (
// Equation(s):
// Xd_0__inst_mult_10_62  = SUM(( (din_a[60] & din_b[61]) ) + ( Xd_0__inst_mult_10_60  ) + ( Xd_0__inst_mult_10_59  ))
// Xd_0__inst_mult_10_63  = CARRY(( (din_a[60] & din_b[61]) ) + ( Xd_0__inst_mult_10_60  ) + ( Xd_0__inst_mult_10_59  ))
// Xd_0__inst_mult_10_64  = SHARE((din_b[60] & din_a[62]))

	.dataa(!din_a[60]),
	.datab(!din_b[60]),
	.datac(!din_b[61]),
	.datad(!din_a[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_59 ),
	.sharein(Xd_0__inst_mult_10_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_62 ),
	.cout(Xd_0__inst_mult_10_63 ),
	.shareout(Xd_0__inst_mult_10_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_11_25 (
// Equation(s):
// Xd_0__inst_mult_11_79  = SUM(( (din_a[66] & din_b[67]) ) + ( Xd_0__inst_mult_11_73  ) + ( Xd_0__inst_mult_11_72  ))
// Xd_0__inst_mult_11_80  = CARRY(( (din_a[66] & din_b[67]) ) + ( Xd_0__inst_mult_11_73  ) + ( Xd_0__inst_mult_11_72  ))
// Xd_0__inst_mult_11_81  = SHARE((din_b[66] & din_a[68]))

	.dataa(!din_a[66]),
	.datab(!din_b[66]),
	.datac(!din_b[67]),
	.datad(!din_a[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_72 ),
	.sharein(Xd_0__inst_mult_11_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_79 ),
	.cout(Xd_0__inst_mult_11_80 ),
	.shareout(Xd_0__inst_mult_11_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_8_21 (
// Equation(s):
// Xd_0__inst_mult_8_62  = SUM(( (din_a[48] & din_b[49]) ) + ( Xd_0__inst_mult_8_60  ) + ( Xd_0__inst_mult_8_59  ))
// Xd_0__inst_mult_8_63  = CARRY(( (din_a[48] & din_b[49]) ) + ( Xd_0__inst_mult_8_60  ) + ( Xd_0__inst_mult_8_59  ))
// Xd_0__inst_mult_8_64  = SHARE((din_b[48] & din_a[50]))

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(!din_b[49]),
	.datad(!din_a[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_59 ),
	.sharein(Xd_0__inst_mult_8_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_62 ),
	.cout(Xd_0__inst_mult_8_63 ),
	.shareout(Xd_0__inst_mult_8_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_9_23 (
// Equation(s):
// Xd_0__inst_mult_9_71  = SUM(( (din_a[54] & din_b[55]) ) + ( Xd_0__inst_mult_9_69  ) + ( Xd_0__inst_mult_9_68  ))
// Xd_0__inst_mult_9_72  = CARRY(( (din_a[54] & din_b[55]) ) + ( Xd_0__inst_mult_9_69  ) + ( Xd_0__inst_mult_9_68  ))
// Xd_0__inst_mult_9_73  = SHARE((din_b[54] & din_a[56]))

	.dataa(!din_a[54]),
	.datab(!din_b[54]),
	.datac(!din_b[55]),
	.datad(!din_a[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_68 ),
	.sharein(Xd_0__inst_mult_9_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_71 ),
	.cout(Xd_0__inst_mult_9_72 ),
	.shareout(Xd_0__inst_mult_9_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_6_21 (
// Equation(s):
// Xd_0__inst_mult_6_61  = SUM(( (din_a[36] & din_b[37]) ) + ( Xd_0__inst_mult_6_59  ) + ( Xd_0__inst_mult_6_58  ))
// Xd_0__inst_mult_6_62  = CARRY(( (din_a[36] & din_b[37]) ) + ( Xd_0__inst_mult_6_59  ) + ( Xd_0__inst_mult_6_58  ))
// Xd_0__inst_mult_6_63  = SHARE((din_b[36] & din_a[38]))

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(!din_a[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_58 ),
	.sharein(Xd_0__inst_mult_6_59 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_61 ),
	.cout(Xd_0__inst_mult_6_62 ),
	.shareout(Xd_0__inst_mult_6_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_7_23 (
// Equation(s):
// Xd_0__inst_mult_7_70  = SUM(( (din_a[42] & din_b[43]) ) + ( Xd_0__inst_mult_7_68  ) + ( Xd_0__inst_mult_7_67  ))
// Xd_0__inst_mult_7_71  = CARRY(( (din_a[42] & din_b[43]) ) + ( Xd_0__inst_mult_7_68  ) + ( Xd_0__inst_mult_7_67  ))
// Xd_0__inst_mult_7_72  = SHARE((din_b[42] & din_a[44]))

	.dataa(!din_a[42]),
	.datab(!din_b[42]),
	.datac(!din_b[43]),
	.datad(!din_a[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_67 ),
	.sharein(Xd_0__inst_mult_7_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_70 ),
	.cout(Xd_0__inst_mult_7_71 ),
	.shareout(Xd_0__inst_mult_7_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_4_21 (
// Equation(s):
// Xd_0__inst_mult_4_61  = SUM(( (din_a[24] & din_b[25]) ) + ( Xd_0__inst_mult_4_59  ) + ( Xd_0__inst_mult_4_58  ))
// Xd_0__inst_mult_4_62  = CARRY(( (din_a[24] & din_b[25]) ) + ( Xd_0__inst_mult_4_59  ) + ( Xd_0__inst_mult_4_58  ))
// Xd_0__inst_mult_4_63  = SHARE((din_b[24] & din_a[26]))

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(!din_b[25]),
	.datad(!din_a[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_58 ),
	.sharein(Xd_0__inst_mult_4_59 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_61 ),
	.cout(Xd_0__inst_mult_4_62 ),
	.shareout(Xd_0__inst_mult_4_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_5_23 (
// Equation(s):
// Xd_0__inst_mult_5_70  = SUM(( (din_a[30] & din_b[31]) ) + ( Xd_0__inst_mult_5_68  ) + ( Xd_0__inst_mult_5_67  ))
// Xd_0__inst_mult_5_71  = CARRY(( (din_a[30] & din_b[31]) ) + ( Xd_0__inst_mult_5_68  ) + ( Xd_0__inst_mult_5_67  ))
// Xd_0__inst_mult_5_72  = SHARE((din_b[30] & din_a[32]))

	.dataa(!din_a[30]),
	.datab(!din_b[30]),
	.datac(!din_b[31]),
	.datad(!din_a[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_67 ),
	.sharein(Xd_0__inst_mult_5_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_70 ),
	.cout(Xd_0__inst_mult_5_71 ),
	.shareout(Xd_0__inst_mult_5_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_2_23 (
// Equation(s):
// Xd_0__inst_mult_2_70  = SUM(( (din_a[12] & din_b[13]) ) + ( Xd_0__inst_mult_2_68  ) + ( Xd_0__inst_mult_2_67  ))
// Xd_0__inst_mult_2_71  = CARRY(( (din_a[12] & din_b[13]) ) + ( Xd_0__inst_mult_2_68  ) + ( Xd_0__inst_mult_2_67  ))
// Xd_0__inst_mult_2_72  = SHARE((din_b[12] & din_a[14]))

	.dataa(!din_a[12]),
	.datab(!din_b[12]),
	.datac(!din_b[13]),
	.datad(!din_a[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_67 ),
	.sharein(Xd_0__inst_mult_2_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_70 ),
	.cout(Xd_0__inst_mult_2_71 ),
	.shareout(Xd_0__inst_mult_2_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_3_23 (
// Equation(s):
// Xd_0__inst_mult_3_70  = SUM(( (din_a[18] & din_b[19]) ) + ( Xd_0__inst_mult_3_68  ) + ( Xd_0__inst_mult_3_67  ))
// Xd_0__inst_mult_3_71  = CARRY(( (din_a[18] & din_b[19]) ) + ( Xd_0__inst_mult_3_68  ) + ( Xd_0__inst_mult_3_67  ))
// Xd_0__inst_mult_3_72  = SHARE((din_b[18] & din_a[20]))

	.dataa(!din_a[18]),
	.datab(!din_b[18]),
	.datac(!din_b[19]),
	.datad(!din_a[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_67 ),
	.sharein(Xd_0__inst_mult_3_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_70 ),
	.cout(Xd_0__inst_mult_3_71 ),
	.shareout(Xd_0__inst_mult_3_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_0_23 (
// Equation(s):
// Xd_0__inst_mult_0_70  = SUM(( (din_a[0] & din_b[1]) ) + ( Xd_0__inst_mult_0_68  ) + ( Xd_0__inst_mult_0_67  ))
// Xd_0__inst_mult_0_71  = CARRY(( (din_a[0] & din_b[1]) ) + ( Xd_0__inst_mult_0_68  ) + ( Xd_0__inst_mult_0_67  ))
// Xd_0__inst_mult_0_72  = SHARE((din_b[0] & din_a[2]))

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(!din_a[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_67 ),
	.sharein(Xd_0__inst_mult_0_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_70 ),
	.cout(Xd_0__inst_mult_0_71 ),
	.shareout(Xd_0__inst_mult_0_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_1_23 (
// Equation(s):
// Xd_0__inst_mult_1_70  = SUM(( (din_a[6] & din_b[7]) ) + ( Xd_0__inst_mult_1_68  ) + ( Xd_0__inst_mult_1_67  ))
// Xd_0__inst_mult_1_71  = CARRY(( (din_a[6] & din_b[7]) ) + ( Xd_0__inst_mult_1_68  ) + ( Xd_0__inst_mult_1_67  ))
// Xd_0__inst_mult_1_72  = SHARE((din_b[6] & din_a[8]))

	.dataa(!din_a[6]),
	.datab(!din_b[6]),
	.datac(!din_b[7]),
	.datad(!din_a[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_67 ),
	.sharein(Xd_0__inst_mult_1_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_70 ),
	.cout(Xd_0__inst_mult_1_71 ),
	.shareout(Xd_0__inst_mult_1_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_28_26 (
// Equation(s):
// Xd_0__inst_mult_28_83  = SUM(( (din_a[168] & din_b[169]) ) + ( Xd_0__inst_mult_28_81  ) + ( Xd_0__inst_mult_28_80  ))
// Xd_0__inst_mult_28_84  = CARRY(( (din_a[168] & din_b[169]) ) + ( Xd_0__inst_mult_28_81  ) + ( Xd_0__inst_mult_28_80  ))
// Xd_0__inst_mult_28_85  = SHARE((din_b[168] & din_a[170]))

	.dataa(!din_a[168]),
	.datab(!din_b[168]),
	.datac(!din_b[169]),
	.datad(!din_a[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_80 ),
	.sharein(Xd_0__inst_mult_28_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_83 ),
	.cout(Xd_0__inst_mult_28_84 ),
	.shareout(Xd_0__inst_mult_28_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_29_25 (
// Equation(s):
// Xd_0__inst_mult_29_79  = SUM(( (din_a[174] & din_b[175]) ) + ( Xd_0__inst_mult_29_77  ) + ( Xd_0__inst_mult_29_76  ))
// Xd_0__inst_mult_29_80  = CARRY(( (din_a[174] & din_b[175]) ) + ( Xd_0__inst_mult_29_77  ) + ( Xd_0__inst_mult_29_76  ))
// Xd_0__inst_mult_29_81  = SHARE((din_b[174] & din_a[176]))

	.dataa(!din_a[174]),
	.datab(!din_b[174]),
	.datac(!din_b[175]),
	.datad(!din_a[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_76 ),
	.sharein(Xd_0__inst_mult_29_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_79 ),
	.cout(Xd_0__inst_mult_29_80 ),
	.shareout(Xd_0__inst_mult_29_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_26_26 (
// Equation(s):
// Xd_0__inst_mult_26_83  = SUM(( (din_a[156] & din_b[157]) ) + ( Xd_0__inst_mult_26_81  ) + ( Xd_0__inst_mult_26_80  ))
// Xd_0__inst_mult_26_84  = CARRY(( (din_a[156] & din_b[157]) ) + ( Xd_0__inst_mult_26_81  ) + ( Xd_0__inst_mult_26_80  ))
// Xd_0__inst_mult_26_85  = SHARE((din_b[156] & din_a[158]))

	.dataa(!din_a[156]),
	.datab(!din_b[156]),
	.datac(!din_b[157]),
	.datad(!din_a[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_80 ),
	.sharein(Xd_0__inst_mult_26_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_83 ),
	.cout(Xd_0__inst_mult_26_84 ),
	.shareout(Xd_0__inst_mult_26_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_27_25 (
// Equation(s):
// Xd_0__inst_mult_27_79  = SUM(( (din_a[162] & din_b[163]) ) + ( Xd_0__inst_mult_27_73  ) + ( Xd_0__inst_mult_27_72  ))
// Xd_0__inst_mult_27_80  = CARRY(( (din_a[162] & din_b[163]) ) + ( Xd_0__inst_mult_27_73  ) + ( Xd_0__inst_mult_27_72  ))
// Xd_0__inst_mult_27_81  = SHARE((din_b[162] & din_a[164]))

	.dataa(!din_a[162]),
	.datab(!din_b[162]),
	.datac(!din_b[163]),
	.datad(!din_a[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_72 ),
	.sharein(Xd_0__inst_mult_27_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_79 ),
	.cout(Xd_0__inst_mult_27_80 ),
	.shareout(Xd_0__inst_mult_27_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_24_26 (
// Equation(s):
// Xd_0__inst_mult_24_83  = SUM(( (din_a[144] & din_b[145]) ) + ( Xd_0__inst_mult_24_81  ) + ( Xd_0__inst_mult_24_80  ))
// Xd_0__inst_mult_24_84  = CARRY(( (din_a[144] & din_b[145]) ) + ( Xd_0__inst_mult_24_81  ) + ( Xd_0__inst_mult_24_80  ))
// Xd_0__inst_mult_24_85  = SHARE((din_b[144] & din_a[146]))

	.dataa(!din_a[144]),
	.datab(!din_b[144]),
	.datac(!din_b[145]),
	.datad(!din_a[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_80 ),
	.sharein(Xd_0__inst_mult_24_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_83 ),
	.cout(Xd_0__inst_mult_24_84 ),
	.shareout(Xd_0__inst_mult_24_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_25_25 (
// Equation(s):
// Xd_0__inst_mult_25_79  = SUM(( (din_a[150] & din_b[151]) ) + ( Xd_0__inst_mult_25_73  ) + ( Xd_0__inst_mult_25_72  ))
// Xd_0__inst_mult_25_80  = CARRY(( (din_a[150] & din_b[151]) ) + ( Xd_0__inst_mult_25_73  ) + ( Xd_0__inst_mult_25_72  ))
// Xd_0__inst_mult_25_81  = SHARE((din_b[150] & din_a[152]))

	.dataa(!din_a[150]),
	.datab(!din_b[150]),
	.datac(!din_b[151]),
	.datad(!din_a[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_72 ),
	.sharein(Xd_0__inst_mult_25_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_79 ),
	.cout(Xd_0__inst_mult_25_80 ),
	.shareout(Xd_0__inst_mult_25_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_22_26 (
// Equation(s):
// Xd_0__inst_mult_22_83  = SUM(( (din_a[132] & din_b[133]) ) + ( Xd_0__inst_mult_22_81  ) + ( Xd_0__inst_mult_22_80  ))
// Xd_0__inst_mult_22_84  = CARRY(( (din_a[132] & din_b[133]) ) + ( Xd_0__inst_mult_22_81  ) + ( Xd_0__inst_mult_22_80  ))
// Xd_0__inst_mult_22_85  = SHARE((din_b[132] & din_a[134]))

	.dataa(!din_a[132]),
	.datab(!din_b[132]),
	.datac(!din_b[133]),
	.datad(!din_a[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_80 ),
	.sharein(Xd_0__inst_mult_22_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_83 ),
	.cout(Xd_0__inst_mult_22_84 ),
	.shareout(Xd_0__inst_mult_22_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_23_26 (
// Equation(s):
// Xd_0__inst_mult_23_83  = SUM(( (din_a[138] & din_b[139]) ) + ( Xd_0__inst_mult_23_81  ) + ( Xd_0__inst_mult_23_80  ))
// Xd_0__inst_mult_23_84  = CARRY(( (din_a[138] & din_b[139]) ) + ( Xd_0__inst_mult_23_81  ) + ( Xd_0__inst_mult_23_80  ))
// Xd_0__inst_mult_23_85  = SHARE((din_b[138] & din_a[140]))

	.dataa(!din_a[138]),
	.datab(!din_b[138]),
	.datac(!din_b[139]),
	.datad(!din_a[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_80 ),
	.sharein(Xd_0__inst_mult_23_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_83 ),
	.cout(Xd_0__inst_mult_23_84 ),
	.shareout(Xd_0__inst_mult_23_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_20_26 (
// Equation(s):
// Xd_0__inst_mult_20_83  = SUM(( (din_a[120] & din_b[121]) ) + ( Xd_0__inst_mult_20_81  ) + ( Xd_0__inst_mult_20_80  ))
// Xd_0__inst_mult_20_84  = CARRY(( (din_a[120] & din_b[121]) ) + ( Xd_0__inst_mult_20_81  ) + ( Xd_0__inst_mult_20_80  ))
// Xd_0__inst_mult_20_85  = SHARE((din_b[120] & din_a[122]))

	.dataa(!din_a[120]),
	.datab(!din_b[120]),
	.datac(!din_b[121]),
	.datad(!din_a[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_80 ),
	.sharein(Xd_0__inst_mult_20_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_83 ),
	.cout(Xd_0__inst_mult_20_84 ),
	.shareout(Xd_0__inst_mult_20_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_21_23 (
// Equation(s):
// Xd_0__inst_mult_21_71  = SUM(( (din_a[126] & din_b[127]) ) + ( Xd_0__inst_mult_21_69  ) + ( Xd_0__inst_mult_21_68  ))
// Xd_0__inst_mult_21_72  = CARRY(( (din_a[126] & din_b[127]) ) + ( Xd_0__inst_mult_21_69  ) + ( Xd_0__inst_mult_21_68  ))
// Xd_0__inst_mult_21_73  = SHARE((din_b[126] & din_a[128]))

	.dataa(!din_a[126]),
	.datab(!din_b[126]),
	.datac(!din_b[127]),
	.datad(!din_a[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_68 ),
	.sharein(Xd_0__inst_mult_21_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_71 ),
	.cout(Xd_0__inst_mult_21_72 ),
	.shareout(Xd_0__inst_mult_21_73 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_18_21 (
// Equation(s):
// Xd_0__inst_mult_18_62  = SUM(( (din_a[108] & din_b[109]) ) + ( Xd_0__inst_mult_18_60  ) + ( Xd_0__inst_mult_18_59  ))
// Xd_0__inst_mult_18_63  = CARRY(( (din_a[108] & din_b[109]) ) + ( Xd_0__inst_mult_18_60  ) + ( Xd_0__inst_mult_18_59  ))
// Xd_0__inst_mult_18_64  = SHARE((din_b[108] & din_a[110]))

	.dataa(!din_a[108]),
	.datab(!din_b[108]),
	.datac(!din_b[109]),
	.datad(!din_a[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_59 ),
	.sharein(Xd_0__inst_mult_18_60 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_62 ),
	.cout(Xd_0__inst_mult_18_63 ),
	.shareout(Xd_0__inst_mult_18_64 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000003300000505),
	.shared_arith("on")
) Xd_0__inst_mult_19_26 (
// Equation(s):
// Xd_0__inst_mult_19_83  = SUM(( (din_a[114] & din_b[115]) ) + ( Xd_0__inst_mult_19_81  ) + ( Xd_0__inst_mult_19_80  ))
// Xd_0__inst_mult_19_84  = CARRY(( (din_a[114] & din_b[115]) ) + ( Xd_0__inst_mult_19_81  ) + ( Xd_0__inst_mult_19_80  ))
// Xd_0__inst_mult_19_85  = SHARE((din_b[114] & din_a[116]))

	.dataa(!din_a[114]),
	.datab(!din_b[114]),
	.datac(!din_b[115]),
	.datad(!din_a[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_80 ),
	.sharein(Xd_0__inst_mult_19_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_83 ),
	.cout(Xd_0__inst_mult_19_84 ),
	.shareout(Xd_0__inst_mult_19_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_22 (
// Equation(s):
// Xd_0__inst_mult_16_66  = SUM(( (!din_a[97] & (((din_a[96] & din_b[98])))) # (din_a[97] & (!din_b[97] $ (((!din_a[96]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_16_64  ) + ( Xd_0__inst_mult_16_63  ))
// Xd_0__inst_mult_16_67  = CARRY(( (!din_a[97] & (((din_a[96] & din_b[98])))) # (din_a[97] & (!din_b[97] $ (((!din_a[96]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_16_64  ) + ( Xd_0__inst_mult_16_63  ))
// Xd_0__inst_mult_16_68  = SHARE((din_a[97] & (din_b[97] & (din_a[96] & din_b[98]))))

	.dataa(!din_a[97]),
	.datab(!din_b[97]),
	.datac(!din_a[96]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_63 ),
	.sharein(Xd_0__inst_mult_16_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_66 ),
	.cout(Xd_0__inst_mult_16_67 ),
	.shareout(Xd_0__inst_mult_16_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_24 (
// Equation(s):
// Xd_0__inst_mult_17_75  = SUM(( (!din_a[103] & (((din_a[102] & din_b[104])))) # (din_a[103] & (!din_b[103] $ (((!din_a[102]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_17_73  ) + ( Xd_0__inst_mult_17_72  ))
// Xd_0__inst_mult_17_76  = CARRY(( (!din_a[103] & (((din_a[102] & din_b[104])))) # (din_a[103] & (!din_b[103] $ (((!din_a[102]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_17_73  ) + ( Xd_0__inst_mult_17_72  ))
// Xd_0__inst_mult_17_77  = SHARE((din_a[103] & (din_b[103] & (din_a[102] & din_b[104]))))

	.dataa(!din_a[103]),
	.datab(!din_b[103]),
	.datac(!din_a[102]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_72 ),
	.sharein(Xd_0__inst_mult_17_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_75 ),
	.cout(Xd_0__inst_mult_17_76 ),
	.shareout(Xd_0__inst_mult_17_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_22 (
// Equation(s):
// Xd_0__inst_mult_14_66  = SUM(( (!din_a[85] & (((din_a[84] & din_b[86])))) # (din_a[85] & (!din_b[85] $ (((!din_a[84]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_14_64  ) + ( Xd_0__inst_mult_14_63  ))
// Xd_0__inst_mult_14_67  = CARRY(( (!din_a[85] & (((din_a[84] & din_b[86])))) # (din_a[85] & (!din_b[85] $ (((!din_a[84]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_14_64  ) + ( Xd_0__inst_mult_14_63  ))
// Xd_0__inst_mult_14_68  = SHARE((din_a[85] & (din_b[85] & (din_a[84] & din_b[86]))))

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[84]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_63 ),
	.sharein(Xd_0__inst_mult_14_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_66 ),
	.cout(Xd_0__inst_mult_14_67 ),
	.shareout(Xd_0__inst_mult_14_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_24 (
// Equation(s):
// Xd_0__inst_mult_15_75  = SUM(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_15_73  ) + ( Xd_0__inst_mult_15_72  ))
// Xd_0__inst_mult_15_76  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_15_73  ) + ( Xd_0__inst_mult_15_72  ))
// Xd_0__inst_mult_15_77  = SHARE((din_a[91] & (din_b[91] & (din_a[90] & din_b[92]))))

	.dataa(!din_a[91]),
	.datab(!din_b[91]),
	.datac(!din_a[90]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_72 ),
	.sharein(Xd_0__inst_mult_15_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_75 ),
	.cout(Xd_0__inst_mult_15_76 ),
	.shareout(Xd_0__inst_mult_15_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_22 (
// Equation(s):
// Xd_0__inst_mult_12_66  = SUM(( (!din_a[73] & (((din_a[72] & din_b[74])))) # (din_a[73] & (!din_b[73] $ (((!din_a[72]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_12_64  ) + ( Xd_0__inst_mult_12_63  ))
// Xd_0__inst_mult_12_67  = CARRY(( (!din_a[73] & (((din_a[72] & din_b[74])))) # (din_a[73] & (!din_b[73] $ (((!din_a[72]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_12_64  ) + ( Xd_0__inst_mult_12_63  ))
// Xd_0__inst_mult_12_68  = SHARE((din_a[73] & (din_b[73] & (din_a[72] & din_b[74]))))

	.dataa(!din_a[73]),
	.datab(!din_b[73]),
	.datac(!din_a[72]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_63 ),
	.sharein(Xd_0__inst_mult_12_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_66 ),
	.cout(Xd_0__inst_mult_12_67 ),
	.shareout(Xd_0__inst_mult_12_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_24 (
// Equation(s):
// Xd_0__inst_mult_13_75  = SUM(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_13_73  ) + ( Xd_0__inst_mult_13_72  ))
// Xd_0__inst_mult_13_76  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_13_73  ) + ( Xd_0__inst_mult_13_72  ))
// Xd_0__inst_mult_13_77  = SHARE((din_a[79] & (din_b[79] & (din_a[78] & din_b[80]))))

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(!din_a[78]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_72 ),
	.sharein(Xd_0__inst_mult_13_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_75 ),
	.cout(Xd_0__inst_mult_13_76 ),
	.shareout(Xd_0__inst_mult_13_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_22 (
// Equation(s):
// Xd_0__inst_mult_10_66  = SUM(( (!din_a[61] & (((din_a[60] & din_b[62])))) # (din_a[61] & (!din_b[61] $ (((!din_a[60]) # (!din_b[62]))))) ) + ( Xd_0__inst_mult_10_64  ) + ( Xd_0__inst_mult_10_63  ))
// Xd_0__inst_mult_10_67  = CARRY(( (!din_a[61] & (((din_a[60] & din_b[62])))) # (din_a[61] & (!din_b[61] $ (((!din_a[60]) # (!din_b[62]))))) ) + ( Xd_0__inst_mult_10_64  ) + ( Xd_0__inst_mult_10_63  ))
// Xd_0__inst_mult_10_68  = SHARE((din_a[61] & (din_b[61] & (din_a[60] & din_b[62]))))

	.dataa(!din_a[61]),
	.datab(!din_b[61]),
	.datac(!din_a[60]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_63 ),
	.sharein(Xd_0__inst_mult_10_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_66 ),
	.cout(Xd_0__inst_mult_10_67 ),
	.shareout(Xd_0__inst_mult_10_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_26 (
// Equation(s):
// Xd_0__inst_mult_11_83  = SUM(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_11_81  ) + ( Xd_0__inst_mult_11_80  ))
// Xd_0__inst_mult_11_84  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_11_81  ) + ( Xd_0__inst_mult_11_80  ))
// Xd_0__inst_mult_11_85  = SHARE((din_a[67] & (din_b[67] & (din_a[66] & din_b[68]))))

	.dataa(!din_a[67]),
	.datab(!din_b[67]),
	.datac(!din_a[66]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_80 ),
	.sharein(Xd_0__inst_mult_11_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_83 ),
	.cout(Xd_0__inst_mult_11_84 ),
	.shareout(Xd_0__inst_mult_11_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_22 (
// Equation(s):
// Xd_0__inst_mult_8_66  = SUM(( (!din_a[49] & (((din_a[48] & din_b[50])))) # (din_a[49] & (!din_b[49] $ (((!din_a[48]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_8_64  ) + ( Xd_0__inst_mult_8_63  ))
// Xd_0__inst_mult_8_67  = CARRY(( (!din_a[49] & (((din_a[48] & din_b[50])))) # (din_a[49] & (!din_b[49] $ (((!din_a[48]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_8_64  ) + ( Xd_0__inst_mult_8_63  ))
// Xd_0__inst_mult_8_68  = SHARE((din_a[49] & (din_b[49] & (din_a[48] & din_b[50]))))

	.dataa(!din_a[49]),
	.datab(!din_b[49]),
	.datac(!din_a[48]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_63 ),
	.sharein(Xd_0__inst_mult_8_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_66 ),
	.cout(Xd_0__inst_mult_8_67 ),
	.shareout(Xd_0__inst_mult_8_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_24 (
// Equation(s):
// Xd_0__inst_mult_9_75  = SUM(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_9_73  ) + ( Xd_0__inst_mult_9_72  ))
// Xd_0__inst_mult_9_76  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_9_73  ) + ( Xd_0__inst_mult_9_72  ))
// Xd_0__inst_mult_9_77  = SHARE((din_a[55] & (din_b[55] & (din_a[54] & din_b[56]))))

	.dataa(!din_a[55]),
	.datab(!din_b[55]),
	.datac(!din_a[54]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_72 ),
	.sharein(Xd_0__inst_mult_9_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_75 ),
	.cout(Xd_0__inst_mult_9_76 ),
	.shareout(Xd_0__inst_mult_9_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_22 (
// Equation(s):
// Xd_0__inst_mult_6_65  = SUM(( (!din_a[37] & (((din_a[36] & din_b[38])))) # (din_a[37] & (!din_b[37] $ (((!din_a[36]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_6_63  ) + ( Xd_0__inst_mult_6_62  ))
// Xd_0__inst_mult_6_66  = CARRY(( (!din_a[37] & (((din_a[36] & din_b[38])))) # (din_a[37] & (!din_b[37] $ (((!din_a[36]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_6_63  ) + ( Xd_0__inst_mult_6_62  ))
// Xd_0__inst_mult_6_67  = SHARE((din_a[37] & (din_b[37] & (din_a[36] & din_b[38]))))

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[36]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_62 ),
	.sharein(Xd_0__inst_mult_6_63 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_65 ),
	.cout(Xd_0__inst_mult_6_66 ),
	.shareout(Xd_0__inst_mult_6_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_24 (
// Equation(s):
// Xd_0__inst_mult_7_74  = SUM(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_7_72  ) + ( Xd_0__inst_mult_7_71  ))
// Xd_0__inst_mult_7_75  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_7_72  ) + ( Xd_0__inst_mult_7_71  ))
// Xd_0__inst_mult_7_76  = SHARE((din_a[43] & (din_b[43] & (din_a[42] & din_b[44]))))

	.dataa(!din_a[43]),
	.datab(!din_b[43]),
	.datac(!din_a[42]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_71 ),
	.sharein(Xd_0__inst_mult_7_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_74 ),
	.cout(Xd_0__inst_mult_7_75 ),
	.shareout(Xd_0__inst_mult_7_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_22 (
// Equation(s):
// Xd_0__inst_mult_4_65  = SUM(( (!din_a[25] & (((din_a[24] & din_b[26])))) # (din_a[25] & (!din_b[25] $ (((!din_a[24]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_4_63  ) + ( Xd_0__inst_mult_4_62  ))
// Xd_0__inst_mult_4_66  = CARRY(( (!din_a[25] & (((din_a[24] & din_b[26])))) # (din_a[25] & (!din_b[25] $ (((!din_a[24]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_4_63  ) + ( Xd_0__inst_mult_4_62  ))
// Xd_0__inst_mult_4_67  = SHARE((din_a[25] & (din_b[25] & (din_a[24] & din_b[26]))))

	.dataa(!din_a[25]),
	.datab(!din_b[25]),
	.datac(!din_a[24]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_62 ),
	.sharein(Xd_0__inst_mult_4_63 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_65 ),
	.cout(Xd_0__inst_mult_4_66 ),
	.shareout(Xd_0__inst_mult_4_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_24 (
// Equation(s):
// Xd_0__inst_mult_5_74  = SUM(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_5_72  ) + ( Xd_0__inst_mult_5_71  ))
// Xd_0__inst_mult_5_75  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_5_72  ) + ( Xd_0__inst_mult_5_71  ))
// Xd_0__inst_mult_5_76  = SHARE((din_a[31] & (din_b[31] & (din_a[30] & din_b[32]))))

	.dataa(!din_a[31]),
	.datab(!din_b[31]),
	.datac(!din_a[30]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_71 ),
	.sharein(Xd_0__inst_mult_5_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_74 ),
	.cout(Xd_0__inst_mult_5_75 ),
	.shareout(Xd_0__inst_mult_5_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_24 (
// Equation(s):
// Xd_0__inst_mult_2_74  = SUM(( (!din_a[13] & (((din_a[12] & din_b[14])))) # (din_a[13] & (!din_b[13] $ (((!din_a[12]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_72  ) + ( Xd_0__inst_mult_2_71  ))
// Xd_0__inst_mult_2_75  = CARRY(( (!din_a[13] & (((din_a[12] & din_b[14])))) # (din_a[13] & (!din_b[13] $ (((!din_a[12]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_72  ) + ( Xd_0__inst_mult_2_71  ))
// Xd_0__inst_mult_2_76  = SHARE((din_a[13] & (din_b[13] & (din_a[12] & din_b[14]))))

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(!din_a[12]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_71 ),
	.sharein(Xd_0__inst_mult_2_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_74 ),
	.cout(Xd_0__inst_mult_2_75 ),
	.shareout(Xd_0__inst_mult_2_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_24 (
// Equation(s):
// Xd_0__inst_mult_3_74  = SUM(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_3_72  ) + ( Xd_0__inst_mult_3_71  ))
// Xd_0__inst_mult_3_75  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_3_72  ) + ( Xd_0__inst_mult_3_71  ))
// Xd_0__inst_mult_3_76  = SHARE((din_a[19] & (din_b[19] & (din_a[18] & din_b[20]))))

	.dataa(!din_a[19]),
	.datab(!din_b[19]),
	.datac(!din_a[18]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_71 ),
	.sharein(Xd_0__inst_mult_3_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_74 ),
	.cout(Xd_0__inst_mult_3_75 ),
	.shareout(Xd_0__inst_mult_3_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_24 (
// Equation(s):
// Xd_0__inst_mult_0_74  = SUM(( (!din_a[1] & (((din_a[0] & din_b[2])))) # (din_a[1] & (!din_b[1] $ (((!din_a[0]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_72  ) + ( Xd_0__inst_mult_0_71  ))
// Xd_0__inst_mult_0_75  = CARRY(( (!din_a[1] & (((din_a[0] & din_b[2])))) # (din_a[1] & (!din_b[1] $ (((!din_a[0]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_72  ) + ( Xd_0__inst_mult_0_71  ))
// Xd_0__inst_mult_0_76  = SHARE((din_a[1] & (din_b[1] & (din_a[0] & din_b[2]))))

	.dataa(!din_a[1]),
	.datab(!din_b[1]),
	.datac(!din_a[0]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_71 ),
	.sharein(Xd_0__inst_mult_0_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_74 ),
	.cout(Xd_0__inst_mult_0_75 ),
	.shareout(Xd_0__inst_mult_0_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_24 (
// Equation(s):
// Xd_0__inst_mult_1_74  = SUM(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_72  ) + ( Xd_0__inst_mult_1_71  ))
// Xd_0__inst_mult_1_75  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_72  ) + ( Xd_0__inst_mult_1_71  ))
// Xd_0__inst_mult_1_76  = SHARE((din_a[7] & (din_b[7] & (din_a[6] & din_b[8]))))

	.dataa(!din_a[7]),
	.datab(!din_b[7]),
	.datac(!din_a[6]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_71 ),
	.sharein(Xd_0__inst_mult_1_72 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_74 ),
	.cout(Xd_0__inst_mult_1_75 ),
	.shareout(Xd_0__inst_mult_1_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_27 (
// Equation(s):
// Xd_0__inst_mult_28_87  = SUM(( (!din_a[169] & (((din_a[168] & din_b[170])))) # (din_a[169] & (!din_b[169] $ (((!din_a[168]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_28_85  ) + ( Xd_0__inst_mult_28_84  ))
// Xd_0__inst_mult_28_88  = CARRY(( (!din_a[169] & (((din_a[168] & din_b[170])))) # (din_a[169] & (!din_b[169] $ (((!din_a[168]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_28_85  ) + ( Xd_0__inst_mult_28_84  ))
// Xd_0__inst_mult_28_89  = SHARE((din_a[169] & (din_b[169] & (din_a[168] & din_b[170]))))

	.dataa(!din_a[169]),
	.datab(!din_b[169]),
	.datac(!din_a[168]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_84 ),
	.sharein(Xd_0__inst_mult_28_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_87 ),
	.cout(Xd_0__inst_mult_28_88 ),
	.shareout(Xd_0__inst_mult_28_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_26 (
// Equation(s):
// Xd_0__inst_mult_29_83  = SUM(( (!din_a[175] & (((din_a[174] & din_b[176])))) # (din_a[175] & (!din_b[175] $ (((!din_a[174]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_29_81  ) + ( Xd_0__inst_mult_29_80  ))
// Xd_0__inst_mult_29_84  = CARRY(( (!din_a[175] & (((din_a[174] & din_b[176])))) # (din_a[175] & (!din_b[175] $ (((!din_a[174]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_29_81  ) + ( Xd_0__inst_mult_29_80  ))
// Xd_0__inst_mult_29_85  = SHARE((din_a[175] & (din_b[175] & (din_a[174] & din_b[176]))))

	.dataa(!din_a[175]),
	.datab(!din_b[175]),
	.datac(!din_a[174]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_80 ),
	.sharein(Xd_0__inst_mult_29_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_83 ),
	.cout(Xd_0__inst_mult_29_84 ),
	.shareout(Xd_0__inst_mult_29_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_27 (
// Equation(s):
// Xd_0__inst_mult_26_87  = SUM(( (!din_a[157] & (((din_a[156] & din_b[158])))) # (din_a[157] & (!din_b[157] $ (((!din_a[156]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_26_85  ) + ( Xd_0__inst_mult_26_84  ))
// Xd_0__inst_mult_26_88  = CARRY(( (!din_a[157] & (((din_a[156] & din_b[158])))) # (din_a[157] & (!din_b[157] $ (((!din_a[156]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_26_85  ) + ( Xd_0__inst_mult_26_84  ))
// Xd_0__inst_mult_26_89  = SHARE((din_a[157] & (din_b[157] & (din_a[156] & din_b[158]))))

	.dataa(!din_a[157]),
	.datab(!din_b[157]),
	.datac(!din_a[156]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_84 ),
	.sharein(Xd_0__inst_mult_26_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_87 ),
	.cout(Xd_0__inst_mult_26_88 ),
	.shareout(Xd_0__inst_mult_26_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_26 (
// Equation(s):
// Xd_0__inst_mult_27_83  = SUM(( (!din_a[163] & (((din_a[162] & din_b[164])))) # (din_a[163] & (!din_b[163] $ (((!din_a[162]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_27_81  ) + ( Xd_0__inst_mult_27_80  ))
// Xd_0__inst_mult_27_84  = CARRY(( (!din_a[163] & (((din_a[162] & din_b[164])))) # (din_a[163] & (!din_b[163] $ (((!din_a[162]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_27_81  ) + ( Xd_0__inst_mult_27_80  ))
// Xd_0__inst_mult_27_85  = SHARE((din_a[163] & (din_b[163] & (din_a[162] & din_b[164]))))

	.dataa(!din_a[163]),
	.datab(!din_b[163]),
	.datac(!din_a[162]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_80 ),
	.sharein(Xd_0__inst_mult_27_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_83 ),
	.cout(Xd_0__inst_mult_27_84 ),
	.shareout(Xd_0__inst_mult_27_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_27 (
// Equation(s):
// Xd_0__inst_mult_24_87  = SUM(( (!din_a[145] & (((din_a[144] & din_b[146])))) # (din_a[145] & (!din_b[145] $ (((!din_a[144]) # (!din_b[146]))))) ) + ( Xd_0__inst_mult_24_85  ) + ( Xd_0__inst_mult_24_84  ))
// Xd_0__inst_mult_24_88  = CARRY(( (!din_a[145] & (((din_a[144] & din_b[146])))) # (din_a[145] & (!din_b[145] $ (((!din_a[144]) # (!din_b[146]))))) ) + ( Xd_0__inst_mult_24_85  ) + ( Xd_0__inst_mult_24_84  ))
// Xd_0__inst_mult_24_89  = SHARE((din_a[145] & (din_b[145] & (din_a[144] & din_b[146]))))

	.dataa(!din_a[145]),
	.datab(!din_b[145]),
	.datac(!din_a[144]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_84 ),
	.sharein(Xd_0__inst_mult_24_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_87 ),
	.cout(Xd_0__inst_mult_24_88 ),
	.shareout(Xd_0__inst_mult_24_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_26 (
// Equation(s):
// Xd_0__inst_mult_25_83  = SUM(( (!din_a[151] & (((din_a[150] & din_b[152])))) # (din_a[151] & (!din_b[151] $ (((!din_a[150]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_25_81  ) + ( Xd_0__inst_mult_25_80  ))
// Xd_0__inst_mult_25_84  = CARRY(( (!din_a[151] & (((din_a[150] & din_b[152])))) # (din_a[151] & (!din_b[151] $ (((!din_a[150]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_25_81  ) + ( Xd_0__inst_mult_25_80  ))
// Xd_0__inst_mult_25_85  = SHARE((din_a[151] & (din_b[151] & (din_a[150] & din_b[152]))))

	.dataa(!din_a[151]),
	.datab(!din_b[151]),
	.datac(!din_a[150]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_80 ),
	.sharein(Xd_0__inst_mult_25_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_83 ),
	.cout(Xd_0__inst_mult_25_84 ),
	.shareout(Xd_0__inst_mult_25_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_27 (
// Equation(s):
// Xd_0__inst_mult_22_87  = SUM(( (!din_a[133] & (((din_a[132] & din_b[134])))) # (din_a[133] & (!din_b[133] $ (((!din_a[132]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_22_85  ) + ( Xd_0__inst_mult_22_84  ))
// Xd_0__inst_mult_22_88  = CARRY(( (!din_a[133] & (((din_a[132] & din_b[134])))) # (din_a[133] & (!din_b[133] $ (((!din_a[132]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_22_85  ) + ( Xd_0__inst_mult_22_84  ))
// Xd_0__inst_mult_22_89  = SHARE((din_a[133] & (din_b[133] & (din_a[132] & din_b[134]))))

	.dataa(!din_a[133]),
	.datab(!din_b[133]),
	.datac(!din_a[132]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_84 ),
	.sharein(Xd_0__inst_mult_22_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_87 ),
	.cout(Xd_0__inst_mult_22_88 ),
	.shareout(Xd_0__inst_mult_22_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_27 (
// Equation(s):
// Xd_0__inst_mult_23_87  = SUM(( (!din_a[139] & (((din_a[138] & din_b[140])))) # (din_a[139] & (!din_b[139] $ (((!din_a[138]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_23_85  ) + ( Xd_0__inst_mult_23_84  ))
// Xd_0__inst_mult_23_88  = CARRY(( (!din_a[139] & (((din_a[138] & din_b[140])))) # (din_a[139] & (!din_b[139] $ (((!din_a[138]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_23_85  ) + ( Xd_0__inst_mult_23_84  ))
// Xd_0__inst_mult_23_89  = SHARE((din_a[139] & (din_b[139] & (din_a[138] & din_b[140]))))

	.dataa(!din_a[139]),
	.datab(!din_b[139]),
	.datac(!din_a[138]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_84 ),
	.sharein(Xd_0__inst_mult_23_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_87 ),
	.cout(Xd_0__inst_mult_23_88 ),
	.shareout(Xd_0__inst_mult_23_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_27 (
// Equation(s):
// Xd_0__inst_mult_20_87  = SUM(( (!din_a[121] & (((din_a[120] & din_b[122])))) # (din_a[121] & (!din_b[121] $ (((!din_a[120]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_20_85  ) + ( Xd_0__inst_mult_20_84  ))
// Xd_0__inst_mult_20_88  = CARRY(( (!din_a[121] & (((din_a[120] & din_b[122])))) # (din_a[121] & (!din_b[121] $ (((!din_a[120]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_20_85  ) + ( Xd_0__inst_mult_20_84  ))
// Xd_0__inst_mult_20_89  = SHARE((din_a[121] & (din_b[121] & (din_a[120] & din_b[122]))))

	.dataa(!din_a[121]),
	.datab(!din_b[121]),
	.datac(!din_a[120]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_84 ),
	.sharein(Xd_0__inst_mult_20_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_87 ),
	.cout(Xd_0__inst_mult_20_88 ),
	.shareout(Xd_0__inst_mult_20_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_24 (
// Equation(s):
// Xd_0__inst_mult_21_75  = SUM(( (!din_a[127] & (((din_a[126] & din_b[128])))) # (din_a[127] & (!din_b[127] $ (((!din_a[126]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_21_73  ) + ( Xd_0__inst_mult_21_72  ))
// Xd_0__inst_mult_21_76  = CARRY(( (!din_a[127] & (((din_a[126] & din_b[128])))) # (din_a[127] & (!din_b[127] $ (((!din_a[126]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_21_73  ) + ( Xd_0__inst_mult_21_72  ))
// Xd_0__inst_mult_21_77  = SHARE((din_a[127] & (din_b[127] & (din_a[126] & din_b[128]))))

	.dataa(!din_a[127]),
	.datab(!din_b[127]),
	.datac(!din_a[126]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_72 ),
	.sharein(Xd_0__inst_mult_21_73 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_75 ),
	.cout(Xd_0__inst_mult_21_76 ),
	.shareout(Xd_0__inst_mult_21_77 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_22 (
// Equation(s):
// Xd_0__inst_mult_18_66  = SUM(( (!din_a[109] & (((din_a[108] & din_b[110])))) # (din_a[109] & (!din_b[109] $ (((!din_a[108]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_18_64  ) + ( Xd_0__inst_mult_18_63  ))
// Xd_0__inst_mult_18_67  = CARRY(( (!din_a[109] & (((din_a[108] & din_b[110])))) # (din_a[109] & (!din_b[109] $ (((!din_a[108]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_18_64  ) + ( Xd_0__inst_mult_18_63  ))
// Xd_0__inst_mult_18_68  = SHARE((din_a[109] & (din_b[109] & (din_a[108] & din_b[110]))))

	.dataa(!din_a[109]),
	.datab(!din_b[109]),
	.datac(!din_a[108]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_63 ),
	.sharein(Xd_0__inst_mult_18_64 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_66 ),
	.cout(Xd_0__inst_mult_18_67 ),
	.shareout(Xd_0__inst_mult_18_68 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_27 (
// Equation(s):
// Xd_0__inst_mult_19_87  = SUM(( (!din_a[115] & (((din_a[114] & din_b[116])))) # (din_a[115] & (!din_b[115] $ (((!din_a[114]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_19_85  ) + ( Xd_0__inst_mult_19_84  ))
// Xd_0__inst_mult_19_88  = CARRY(( (!din_a[115] & (((din_a[114] & din_b[116])))) # (din_a[115] & (!din_b[115] $ (((!din_a[114]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_19_85  ) + ( Xd_0__inst_mult_19_84  ))
// Xd_0__inst_mult_19_89  = SHARE((din_a[115] & (din_b[115] & (din_a[114] & din_b[116]))))

	.dataa(!din_a[115]),
	.datab(!din_b[115]),
	.datac(!din_a[114]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_84 ),
	.sharein(Xd_0__inst_mult_19_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_87 ),
	.cout(Xd_0__inst_mult_19_88 ),
	.shareout(Xd_0__inst_mult_19_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_23 (
// Equation(s):
// Xd_0__inst_mult_16_71  = CARRY(( (Xd_0__inst_mult_16_0_q  & Xd_0__inst_mult_16_1_q ) ) + ( Xd_0__inst_mult_16_80  ) + ( Xd_0__inst_mult_16_79  ))
// Xd_0__inst_mult_16_72  = SHARE((Xd_0__inst_mult_16_2_q  & Xd_0__inst_mult_16_3_q ))

	.dataa(!Xd_0__inst_mult_16_0_q ),
	.datab(!Xd_0__inst_mult_16_1_q ),
	.datac(!Xd_0__inst_mult_16_2_q ),
	.datad(!Xd_0__inst_mult_16_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_79 ),
	.sharein(Xd_0__inst_mult_16_80 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_71 ),
	.shareout(Xd_0__inst_mult_16_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_25 (
// Equation(s):
// Xd_0__inst_mult_17_80  = CARRY(( (Xd_0__inst_mult_17_0_q  & Xd_0__inst_mult_17_1_q ) ) + ( Xd_0__inst_mult_17_61  ) + ( Xd_0__inst_mult_17_60  ))
// Xd_0__inst_mult_17_81  = SHARE((Xd_0__inst_mult_17_2_q  & Xd_0__inst_mult_17_3_q ))

	.dataa(!Xd_0__inst_mult_17_0_q ),
	.datab(!Xd_0__inst_mult_17_1_q ),
	.datac(!Xd_0__inst_mult_17_2_q ),
	.datad(!Xd_0__inst_mult_17_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_60 ),
	.sharein(Xd_0__inst_mult_17_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_80 ),
	.shareout(Xd_0__inst_mult_17_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_23 (
// Equation(s):
// Xd_0__inst_mult_14_71  = CARRY(( (Xd_0__inst_mult_14_0_q  & Xd_0__inst_mult_14_1_q ) ) + ( Xd_0__inst_mult_14_80  ) + ( Xd_0__inst_mult_14_79  ))
// Xd_0__inst_mult_14_72  = SHARE((Xd_0__inst_mult_14_2_q  & Xd_0__inst_mult_14_3_q ))

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(!Xd_0__inst_mult_14_2_q ),
	.datad(!Xd_0__inst_mult_14_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_79 ),
	.sharein(Xd_0__inst_mult_14_80 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_71 ),
	.shareout(Xd_0__inst_mult_14_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_25 (
// Equation(s):
// Xd_0__inst_mult_15_80  = CARRY(( (Xd_0__inst_mult_15_0_q  & Xd_0__inst_mult_15_1_q ) ) + ( Xd_0__inst_mult_15_61  ) + ( Xd_0__inst_mult_15_60  ))
// Xd_0__inst_mult_15_81  = SHARE((Xd_0__inst_mult_15_2_q  & Xd_0__inst_mult_15_3_q ))

	.dataa(!Xd_0__inst_mult_15_0_q ),
	.datab(!Xd_0__inst_mult_15_1_q ),
	.datac(!Xd_0__inst_mult_15_2_q ),
	.datad(!Xd_0__inst_mult_15_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_60 ),
	.sharein(Xd_0__inst_mult_15_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_80 ),
	.shareout(Xd_0__inst_mult_15_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_23 (
// Equation(s):
// Xd_0__inst_mult_12_71  = CARRY(( (Xd_0__inst_mult_12_0_q  & Xd_0__inst_mult_12_1_q ) ) + ( Xd_0__inst_mult_12_84  ) + ( Xd_0__inst_mult_12_83  ))
// Xd_0__inst_mult_12_72  = SHARE((Xd_0__inst_mult_12_2_q  & Xd_0__inst_mult_12_3_q ))

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(!Xd_0__inst_mult_12_2_q ),
	.datad(!Xd_0__inst_mult_12_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_83 ),
	.sharein(Xd_0__inst_mult_12_84 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_71 ),
	.shareout(Xd_0__inst_mult_12_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_25 (
// Equation(s):
// Xd_0__inst_mult_13_80  = CARRY(( (Xd_0__inst_mult_13_0_q  & Xd_0__inst_mult_13_1_q ) ) + ( Xd_0__inst_mult_13_61  ) + ( Xd_0__inst_mult_13_60  ))
// Xd_0__inst_mult_13_81  = SHARE((Xd_0__inst_mult_13_2_q  & Xd_0__inst_mult_13_3_q ))

	.dataa(!Xd_0__inst_mult_13_0_q ),
	.datab(!Xd_0__inst_mult_13_1_q ),
	.datac(!Xd_0__inst_mult_13_2_q ),
	.datad(!Xd_0__inst_mult_13_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_60 ),
	.sharein(Xd_0__inst_mult_13_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_80 ),
	.shareout(Xd_0__inst_mult_13_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_23 (
// Equation(s):
// Xd_0__inst_mult_10_71  = CARRY(( (Xd_0__inst_mult_10_0_q  & Xd_0__inst_mult_10_1_q ) ) + ( Xd_0__inst_mult_10_80  ) + ( Xd_0__inst_mult_10_79  ))
// Xd_0__inst_mult_10_72  = SHARE((Xd_0__inst_mult_10_2_q  & Xd_0__inst_mult_10_3_q ))

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(!Xd_0__inst_mult_10_2_q ),
	.datad(!Xd_0__inst_mult_10_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_79 ),
	.sharein(Xd_0__inst_mult_10_80 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_71 ),
	.shareout(Xd_0__inst_mult_10_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_27 (
// Equation(s):
// Xd_0__inst_mult_11_88  = CARRY(( (Xd_0__inst_mult_11_0_q  & Xd_0__inst_mult_11_1_q ) ) + ( Xd_0__inst_mult_11_38  ) + ( Xd_0__inst_mult_11_37  ))
// Xd_0__inst_mult_11_89  = SHARE((Xd_0__inst_mult_11_2_q  & Xd_0__inst_mult_11_3_q ))

	.dataa(!Xd_0__inst_mult_11_0_q ),
	.datab(!Xd_0__inst_mult_11_1_q ),
	.datac(!Xd_0__inst_mult_11_2_q ),
	.datad(!Xd_0__inst_mult_11_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_37 ),
	.sharein(Xd_0__inst_mult_11_38 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_88 ),
	.shareout(Xd_0__inst_mult_11_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_23 (
// Equation(s):
// Xd_0__inst_mult_8_71  = CARRY(( (Xd_0__inst_mult_8_0_q  & Xd_0__inst_mult_8_1_q ) ) + ( Xd_0__inst_mult_8_84  ) + ( Xd_0__inst_mult_8_83  ))
// Xd_0__inst_mult_8_72  = SHARE((Xd_0__inst_mult_8_2_q  & Xd_0__inst_mult_8_3_q ))

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(!Xd_0__inst_mult_8_2_q ),
	.datad(!Xd_0__inst_mult_8_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_83 ),
	.sharein(Xd_0__inst_mult_8_84 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_71 ),
	.shareout(Xd_0__inst_mult_8_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_25 (
// Equation(s):
// Xd_0__inst_mult_9_80  = CARRY(( (Xd_0__inst_mult_9_0_q  & Xd_0__inst_mult_9_1_q ) ) + ( Xd_0__inst_mult_9_61  ) + ( Xd_0__inst_mult_9_60  ))
// Xd_0__inst_mult_9_81  = SHARE((Xd_0__inst_mult_9_2_q  & Xd_0__inst_mult_9_3_q ))

	.dataa(!Xd_0__inst_mult_9_0_q ),
	.datab(!Xd_0__inst_mult_9_1_q ),
	.datac(!Xd_0__inst_mult_9_2_q ),
	.datad(!Xd_0__inst_mult_9_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_60 ),
	.sharein(Xd_0__inst_mult_9_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_80 ),
	.shareout(Xd_0__inst_mult_9_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_23 (
// Equation(s):
// Xd_0__inst_mult_6_70  = CARRY(( (Xd_0__inst_mult_6_0_q  & Xd_0__inst_mult_6_1_q ) ) + ( Xd_0__inst_mult_6_79  ) + ( Xd_0__inst_mult_6_78  ))
// Xd_0__inst_mult_6_71  = SHARE((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_3_q ))

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(!Xd_0__inst_mult_6_2_q ),
	.datad(!Xd_0__inst_mult_6_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_78 ),
	.sharein(Xd_0__inst_mult_6_79 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_70 ),
	.shareout(Xd_0__inst_mult_6_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_25 (
// Equation(s):
// Xd_0__inst_mult_7_79  = CARRY(( (Xd_0__inst_mult_7_0_q  & Xd_0__inst_mult_7_1_q ) ) + ( Xd_0__inst_mult_7_60  ) + ( Xd_0__inst_mult_7_59  ))
// Xd_0__inst_mult_7_80  = SHARE((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_3_q ))

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(!Xd_0__inst_mult_7_2_q ),
	.datad(!Xd_0__inst_mult_7_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_59 ),
	.sharein(Xd_0__inst_mult_7_60 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_79 ),
	.shareout(Xd_0__inst_mult_7_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_23 (
// Equation(s):
// Xd_0__inst_mult_4_70  = CARRY(( (Xd_0__inst_mult_4_0_q  & Xd_0__inst_mult_4_1_q ) ) + ( Xd_0__inst_mult_4_79  ) + ( Xd_0__inst_mult_4_78  ))
// Xd_0__inst_mult_4_71  = SHARE((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_3_q ))

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(!Xd_0__inst_mult_4_2_q ),
	.datad(!Xd_0__inst_mult_4_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_78 ),
	.sharein(Xd_0__inst_mult_4_79 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_70 ),
	.shareout(Xd_0__inst_mult_4_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_25 (
// Equation(s):
// Xd_0__inst_mult_5_79  = CARRY(( (Xd_0__inst_mult_5_0_q  & Xd_0__inst_mult_5_1_q ) ) + ( Xd_0__inst_mult_5_60  ) + ( Xd_0__inst_mult_5_59  ))
// Xd_0__inst_mult_5_80  = SHARE((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_3_q ))

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(!Xd_0__inst_mult_5_2_q ),
	.datad(!Xd_0__inst_mult_5_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_59 ),
	.sharein(Xd_0__inst_mult_5_60 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_79 ),
	.shareout(Xd_0__inst_mult_5_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_25 (
// Equation(s):
// Xd_0__inst_mult_2_79  = CARRY(( (Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_1_q ) ) + ( Xd_0__inst_mult_2_37  ) + ( Xd_0__inst_mult_2_36  ))
// Xd_0__inst_mult_2_80  = SHARE((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_3_q ))

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(!Xd_0__inst_mult_2_2_q ),
	.datad(!Xd_0__inst_mult_2_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_36 ),
	.sharein(Xd_0__inst_mult_2_37 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_79 ),
	.shareout(Xd_0__inst_mult_2_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_25 (
// Equation(s):
// Xd_0__inst_mult_3_79  = CARRY(( (Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_1_q ) ) + ( Xd_0__inst_mult_3_37  ) + ( Xd_0__inst_mult_3_36  ))
// Xd_0__inst_mult_3_80  = SHARE((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_3_q ))

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(!Xd_0__inst_mult_3_2_q ),
	.datad(!Xd_0__inst_mult_3_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_36 ),
	.sharein(Xd_0__inst_mult_3_37 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_79 ),
	.shareout(Xd_0__inst_mult_3_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_25 (
// Equation(s):
// Xd_0__inst_mult_0_79  = CARRY(( (Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_1_q ) ) + ( Xd_0__inst_mult_0_37  ) + ( Xd_0__inst_mult_0_36  ))
// Xd_0__inst_mult_0_80  = SHARE((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_3_q ))

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(!Xd_0__inst_mult_0_2_q ),
	.datad(!Xd_0__inst_mult_0_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_36 ),
	.sharein(Xd_0__inst_mult_0_37 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_79 ),
	.shareout(Xd_0__inst_mult_0_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_25 (
// Equation(s):
// Xd_0__inst_mult_1_79  = CARRY(( (Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_1_q ) ) + ( Xd_0__inst_mult_1_37  ) + ( Xd_0__inst_mult_1_36  ))
// Xd_0__inst_mult_1_80  = SHARE((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_3_q ))

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(!Xd_0__inst_mult_1_2_q ),
	.datad(!Xd_0__inst_mult_1_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_36 ),
	.sharein(Xd_0__inst_mult_1_37 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_79 ),
	.shareout(Xd_0__inst_mult_1_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_28 (
// Equation(s):
// Xd_0__inst_mult_28_92  = CARRY(( (Xd_0__inst_mult_28_0_q  & Xd_0__inst_mult_28_1_q ) ) + ( Xd_0__inst_mult_28_45  ) + ( Xd_0__inst_mult_28_44  ))
// Xd_0__inst_mult_28_93  = SHARE((Xd_0__inst_mult_28_2_q  & Xd_0__inst_mult_28_3_q ))

	.dataa(!Xd_0__inst_mult_28_0_q ),
	.datab(!Xd_0__inst_mult_28_1_q ),
	.datac(!Xd_0__inst_mult_28_2_q ),
	.datad(!Xd_0__inst_mult_28_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_44 ),
	.sharein(Xd_0__inst_mult_28_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_28_92 ),
	.shareout(Xd_0__inst_mult_28_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_27 (
// Equation(s):
// Xd_0__inst_mult_29_88  = CARRY(( (Xd_0__inst_mult_29_0_q  & Xd_0__inst_mult_29_1_q ) ) + ( Xd_0__inst_mult_29_38  ) + ( Xd_0__inst_mult_29_37  ))
// Xd_0__inst_mult_29_89  = SHARE((Xd_0__inst_mult_29_2_q  & Xd_0__inst_mult_29_3_q ))

	.dataa(!Xd_0__inst_mult_29_0_q ),
	.datab(!Xd_0__inst_mult_29_1_q ),
	.datac(!Xd_0__inst_mult_29_2_q ),
	.datad(!Xd_0__inst_mult_29_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_37 ),
	.sharein(Xd_0__inst_mult_29_38 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_88 ),
	.shareout(Xd_0__inst_mult_29_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_28 (
// Equation(s):
// Xd_0__inst_mult_26_92  = CARRY(( (Xd_0__inst_mult_26_0_q  & Xd_0__inst_mult_26_1_q ) ) + ( Xd_0__inst_mult_26_45  ) + ( Xd_0__inst_mult_26_44  ))
// Xd_0__inst_mult_26_93  = SHARE((Xd_0__inst_mult_26_2_q  & Xd_0__inst_mult_26_3_q ))

	.dataa(!Xd_0__inst_mult_26_0_q ),
	.datab(!Xd_0__inst_mult_26_1_q ),
	.datac(!Xd_0__inst_mult_26_2_q ),
	.datad(!Xd_0__inst_mult_26_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_44 ),
	.sharein(Xd_0__inst_mult_26_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_26_92 ),
	.shareout(Xd_0__inst_mult_26_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_27 (
// Equation(s):
// Xd_0__inst_mult_27_88  = CARRY(( (Xd_0__inst_mult_27_0_q  & Xd_0__inst_mult_27_1_q ) ) + ( Xd_0__inst_mult_27_38  ) + ( Xd_0__inst_mult_27_37  ))
// Xd_0__inst_mult_27_89  = SHARE((Xd_0__inst_mult_27_2_q  & Xd_0__inst_mult_27_3_q ))

	.dataa(!Xd_0__inst_mult_27_0_q ),
	.datab(!Xd_0__inst_mult_27_1_q ),
	.datac(!Xd_0__inst_mult_27_2_q ),
	.datad(!Xd_0__inst_mult_27_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_37 ),
	.sharein(Xd_0__inst_mult_27_38 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_88 ),
	.shareout(Xd_0__inst_mult_27_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_28 (
// Equation(s):
// Xd_0__inst_mult_24_92  = CARRY(( (Xd_0__inst_mult_24_0_q  & Xd_0__inst_mult_24_1_q ) ) + ( Xd_0__inst_mult_24_49  ) + ( Xd_0__inst_mult_24_48  ))
// Xd_0__inst_mult_24_93  = SHARE((Xd_0__inst_mult_24_2_q  & Xd_0__inst_mult_24_3_q ))

	.dataa(!Xd_0__inst_mult_24_0_q ),
	.datab(!Xd_0__inst_mult_24_1_q ),
	.datac(!Xd_0__inst_mult_24_2_q ),
	.datad(!Xd_0__inst_mult_24_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_48 ),
	.sharein(Xd_0__inst_mult_24_49 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_24_92 ),
	.shareout(Xd_0__inst_mult_24_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_27 (
// Equation(s):
// Xd_0__inst_mult_25_88  = CARRY(( (Xd_0__inst_mult_25_0_q  & Xd_0__inst_mult_25_1_q ) ) + ( Xd_0__inst_mult_25_38  ) + ( Xd_0__inst_mult_25_37  ))
// Xd_0__inst_mult_25_89  = SHARE((Xd_0__inst_mult_25_2_q  & Xd_0__inst_mult_25_3_q ))

	.dataa(!Xd_0__inst_mult_25_0_q ),
	.datab(!Xd_0__inst_mult_25_1_q ),
	.datac(!Xd_0__inst_mult_25_2_q ),
	.datad(!Xd_0__inst_mult_25_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_37 ),
	.sharein(Xd_0__inst_mult_25_38 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_88 ),
	.shareout(Xd_0__inst_mult_25_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_28 (
// Equation(s):
// Xd_0__inst_mult_22_92  = CARRY(( (Xd_0__inst_mult_22_0_q  & Xd_0__inst_mult_22_1_q ) ) + ( Xd_0__inst_mult_22_45  ) + ( Xd_0__inst_mult_22_44  ))
// Xd_0__inst_mult_22_93  = SHARE((Xd_0__inst_mult_22_2_q  & Xd_0__inst_mult_22_3_q ))

	.dataa(!Xd_0__inst_mult_22_0_q ),
	.datab(!Xd_0__inst_mult_22_1_q ),
	.datac(!Xd_0__inst_mult_22_2_q ),
	.datad(!Xd_0__inst_mult_22_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_44 ),
	.sharein(Xd_0__inst_mult_22_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_22_92 ),
	.shareout(Xd_0__inst_mult_22_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_28 (
// Equation(s):
// Xd_0__inst_mult_23_92  = CARRY(( (Xd_0__inst_mult_23_0_q  & Xd_0__inst_mult_23_1_q ) ) + ( Xd_0__inst_mult_23_49  ) + ( Xd_0__inst_mult_23_48  ))
// Xd_0__inst_mult_23_93  = SHARE((Xd_0__inst_mult_23_2_q  & Xd_0__inst_mult_23_3_q ))

	.dataa(!Xd_0__inst_mult_23_0_q ),
	.datab(!Xd_0__inst_mult_23_1_q ),
	.datac(!Xd_0__inst_mult_23_2_q ),
	.datad(!Xd_0__inst_mult_23_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_48 ),
	.sharein(Xd_0__inst_mult_23_49 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_23_92 ),
	.shareout(Xd_0__inst_mult_23_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_28 (
// Equation(s):
// Xd_0__inst_mult_20_92  = CARRY(( (Xd_0__inst_mult_20_0_q  & Xd_0__inst_mult_20_1_q ) ) + ( Xd_0__inst_mult_20_49  ) + ( Xd_0__inst_mult_20_48  ))
// Xd_0__inst_mult_20_93  = SHARE((Xd_0__inst_mult_20_2_q  & Xd_0__inst_mult_20_3_q ))

	.dataa(!Xd_0__inst_mult_20_0_q ),
	.datab(!Xd_0__inst_mult_20_1_q ),
	.datac(!Xd_0__inst_mult_20_2_q ),
	.datad(!Xd_0__inst_mult_20_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_48 ),
	.sharein(Xd_0__inst_mult_20_49 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_20_92 ),
	.shareout(Xd_0__inst_mult_20_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_25 (
// Equation(s):
// Xd_0__inst_mult_21_80  = CARRY(( (Xd_0__inst_mult_21_0_q  & Xd_0__inst_mult_21_1_q ) ) + ( Xd_0__inst_mult_21_61  ) + ( Xd_0__inst_mult_21_60  ))
// Xd_0__inst_mult_21_81  = SHARE((Xd_0__inst_mult_21_2_q  & Xd_0__inst_mult_21_3_q ))

	.dataa(!Xd_0__inst_mult_21_0_q ),
	.datab(!Xd_0__inst_mult_21_1_q ),
	.datac(!Xd_0__inst_mult_21_2_q ),
	.datad(!Xd_0__inst_mult_21_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_60 ),
	.sharein(Xd_0__inst_mult_21_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_80 ),
	.shareout(Xd_0__inst_mult_21_81 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_23 (
// Equation(s):
// Xd_0__inst_mult_18_71  = CARRY(( (Xd_0__inst_mult_18_0_q  & Xd_0__inst_mult_18_1_q ) ) + ( Xd_0__inst_mult_18_80  ) + ( Xd_0__inst_mult_18_79  ))
// Xd_0__inst_mult_18_72  = SHARE((Xd_0__inst_mult_18_2_q  & Xd_0__inst_mult_18_3_q ))

	.dataa(!Xd_0__inst_mult_18_0_q ),
	.datab(!Xd_0__inst_mult_18_1_q ),
	.datac(!Xd_0__inst_mult_18_2_q ),
	.datad(!Xd_0__inst_mult_18_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_79 ),
	.sharein(Xd_0__inst_mult_18_80 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_71 ),
	.shareout(Xd_0__inst_mult_18_72 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_28 (
// Equation(s):
// Xd_0__inst_mult_19_92  = CARRY(( (Xd_0__inst_mult_19_0_q  & Xd_0__inst_mult_19_1_q ) ) + ( Xd_0__inst_mult_19_73  ) + ( Xd_0__inst_mult_19_72  ))
// Xd_0__inst_mult_19_93  = SHARE((Xd_0__inst_mult_19_2_q  & Xd_0__inst_mult_19_3_q ))

	.dataa(!Xd_0__inst_mult_19_0_q ),
	.datab(!Xd_0__inst_mult_19_1_q ),
	.datac(!Xd_0__inst_mult_19_2_q ),
	.datad(!Xd_0__inst_mult_19_3_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_72 ),
	.sharein(Xd_0__inst_mult_19_73 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_19_92 ),
	.shareout(Xd_0__inst_mult_19_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_30 (
// Equation(s):
// Xd_0__inst_mult_30_99  = SUM(( (!din_a[181] & (((din_a[182] & din_b[181])))) # (din_a[181] & (!din_b[182] $ (((!din_a[182]) # (!din_b[181]))))) ) + ( Xd_0__inst_mult_30_89  ) + ( Xd_0__inst_mult_30_88  ))
// Xd_0__inst_mult_30_100  = CARRY(( (!din_a[181] & (((din_a[182] & din_b[181])))) # (din_a[181] & (!din_b[182] $ (((!din_a[182]) # (!din_b[181]))))) ) + ( Xd_0__inst_mult_30_89  ) + ( Xd_0__inst_mult_30_88  ))
// Xd_0__inst_mult_30_101  = SHARE((din_a[181] & (din_b[182] & (din_a[182] & din_b[181]))))

	.dataa(!din_a[181]),
	.datab(!din_b[182]),
	.datac(!din_a[182]),
	.datad(!din_b[181]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_88 ),
	.sharein(Xd_0__inst_mult_30_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_99 ),
	.cout(Xd_0__inst_mult_30_100 ),
	.shareout(Xd_0__inst_mult_30_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_28 (
// Equation(s):
// Xd_0__inst_mult_31_91  = SUM(( (!din_a[187] & (((din_a[188] & din_b[187])))) # (din_a[187] & (!din_b[188] $ (((!din_a[188]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_31_81  ) + ( Xd_0__inst_mult_31_80  ))
// Xd_0__inst_mult_31_92  = CARRY(( (!din_a[187] & (((din_a[188] & din_b[187])))) # (din_a[187] & (!din_b[188] $ (((!din_a[188]) # (!din_b[187]))))) ) + ( Xd_0__inst_mult_31_81  ) + ( Xd_0__inst_mult_31_80  ))
// Xd_0__inst_mult_31_93  = SHARE((din_a[187] & (din_b[188] & (din_a[188] & din_b[187]))))

	.dataa(!din_a[187]),
	.datab(!din_b[188]),
	.datac(!din_a[188]),
	.datad(!din_b[187]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_80 ),
	.sharein(Xd_0__inst_mult_31_81 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_91 ),
	.cout(Xd_0__inst_mult_31_92 ),
	.shareout(Xd_0__inst_mult_31_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_31 (
// Equation(s):
// Xd_0__inst_mult_30_103  = SUM(( (din_a[182] & din_b[182]) ) + ( Xd_0__inst_mult_30_101  ) + ( Xd_0__inst_mult_30_100  ))
// Xd_0__inst_mult_30_104  = CARRY(( (din_a[182] & din_b[182]) ) + ( Xd_0__inst_mult_30_101  ) + ( Xd_0__inst_mult_30_100  ))
// Xd_0__inst_mult_30_105  = SHARE((din_a[182] & din_b[183]))

	.dataa(!din_a[182]),
	.datab(!din_b[182]),
	.datac(!din_b[183]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_100 ),
	.sharein(Xd_0__inst_mult_30_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_103 ),
	.cout(Xd_0__inst_mult_30_104 ),
	.shareout(Xd_0__inst_mult_30_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_29 (
// Equation(s):
// Xd_0__inst_mult_31_95  = SUM(( (din_a[188] & din_b[188]) ) + ( Xd_0__inst_mult_31_93  ) + ( Xd_0__inst_mult_31_92  ))
// Xd_0__inst_mult_31_96  = CARRY(( (din_a[188] & din_b[188]) ) + ( Xd_0__inst_mult_31_93  ) + ( Xd_0__inst_mult_31_92  ))
// Xd_0__inst_mult_31_97  = SHARE((din_a[188] & din_b[189]))

	.dataa(!din_a[188]),
	.datab(!din_b[188]),
	.datac(!din_b[189]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_92 ),
	.sharein(Xd_0__inst_mult_31_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_95 ),
	.cout(Xd_0__inst_mult_31_96 ),
	.shareout(Xd_0__inst_mult_31_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_32 (
// Equation(s):
// Xd_0__inst_mult_30_107  = SUM(( (!din_a[184] & (((din_a[183] & din_b[182])))) # (din_a[184] & (!din_b[181] $ (((!din_a[183]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_30_105  ) + ( Xd_0__inst_mult_30_104  ))
// Xd_0__inst_mult_30_108  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[182])))) # (din_a[184] & (!din_b[181] $ (((!din_a[183]) # (!din_b[182]))))) ) + ( Xd_0__inst_mult_30_105  ) + ( Xd_0__inst_mult_30_104  ))
// Xd_0__inst_mult_30_109  = SHARE((din_a[184] & (din_b[181] & (din_a[183] & din_b[182]))))

	.dataa(!din_a[184]),
	.datab(!din_b[181]),
	.datac(!din_a[183]),
	.datad(!din_b[182]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_104 ),
	.sharein(Xd_0__inst_mult_30_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_107 ),
	.cout(Xd_0__inst_mult_30_108 ),
	.shareout(Xd_0__inst_mult_30_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_30 (
// Equation(s):
// Xd_0__inst_mult_31_99  = SUM(( (!din_a[190] & (((din_a[189] & din_b[188])))) # (din_a[190] & (!din_b[187] $ (((!din_a[189]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_31_97  ) + ( Xd_0__inst_mult_31_96  ))
// Xd_0__inst_mult_31_100  = CARRY(( (!din_a[190] & (((din_a[189] & din_b[188])))) # (din_a[190] & (!din_b[187] $ (((!din_a[189]) # (!din_b[188]))))) ) + ( Xd_0__inst_mult_31_97  ) + ( Xd_0__inst_mult_31_96  ))
// Xd_0__inst_mult_31_101  = SHARE((din_a[190] & (din_b[187] & (din_a[189] & din_b[188]))))

	.dataa(!din_a[190]),
	.datab(!din_b[187]),
	.datac(!din_a[189]),
	.datad(!din_b[188]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_96 ),
	.sharein(Xd_0__inst_mult_31_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_99 ),
	.cout(Xd_0__inst_mult_31_100 ),
	.shareout(Xd_0__inst_mult_31_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_30_33 (
// Equation(s):
// Xd_0__inst_mult_30_111  = SUM(( (!din_a[184] & (((din_a[183] & din_b[183])))) # (din_a[184] & (!din_b[182] $ (((!din_a[183]) # (!din_b[183]))))) ) + ( Xd_0__inst_mult_30_109  ) + ( Xd_0__inst_mult_30_108  ))
// Xd_0__inst_mult_30_112  = CARRY(( (!din_a[184] & (((din_a[183] & din_b[183])))) # (din_a[184] & (!din_b[182] $ (((!din_a[183]) # (!din_b[183]))))) ) + ( Xd_0__inst_mult_30_109  ) + ( Xd_0__inst_mult_30_108  ))
// Xd_0__inst_mult_30_113  = SHARE((din_a[184] & (din_b[182] & (din_a[183] & din_b[183]))))

	.dataa(!din_a[184]),
	.datab(!din_b[182]),
	.datac(!din_a[183]),
	.datad(!din_b[183]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_108 ),
	.sharein(Xd_0__inst_mult_30_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_111 ),
	.cout(Xd_0__inst_mult_30_112 ),
	.shareout(Xd_0__inst_mult_30_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_31_31 (
// Equation(s):
// Xd_0__inst_mult_31_103  = SUM(( (!din_a[190] & (((din_a[189] & din_b[189])))) # (din_a[190] & (!din_b[188] $ (((!din_a[189]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_31_101  ) + ( Xd_0__inst_mult_31_100  ))
// Xd_0__inst_mult_31_104  = CARRY(( (!din_a[190] & (((din_a[189] & din_b[189])))) # (din_a[190] & (!din_b[188] $ (((!din_a[189]) # (!din_b[189]))))) ) + ( Xd_0__inst_mult_31_101  ) + ( Xd_0__inst_mult_31_100  ))
// Xd_0__inst_mult_31_105  = SHARE((din_a[190] & (din_b[188] & (din_a[189] & din_b[189]))))

	.dataa(!din_a[190]),
	.datab(!din_b[188]),
	.datac(!din_a[189]),
	.datad(!din_b[189]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_100 ),
	.sharein(Xd_0__inst_mult_31_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_103 ),
	.cout(Xd_0__inst_mult_31_104 ),
	.shareout(Xd_0__inst_mult_31_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_30_34 (
// Equation(s):
// Xd_0__inst_mult_30_115  = SUM(( (din_a[184] & din_b[183]) ) + ( Xd_0__inst_mult_30_113  ) + ( Xd_0__inst_mult_30_112  ))
// Xd_0__inst_mult_30_116  = CARRY(( (din_a[184] & din_b[183]) ) + ( Xd_0__inst_mult_30_113  ) + ( Xd_0__inst_mult_30_112  ))
// Xd_0__inst_mult_30_117  = SHARE(GND)

	.dataa(!din_a[184]),
	.datab(!din_b[183]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_30_112 ),
	.sharein(Xd_0__inst_mult_30_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_30_115 ),
	.cout(Xd_0__inst_mult_30_116 ),
	.shareout(Xd_0__inst_mult_30_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_31_32 (
// Equation(s):
// Xd_0__inst_mult_31_107  = SUM(( (din_a[190] & din_b[189]) ) + ( Xd_0__inst_mult_31_105  ) + ( Xd_0__inst_mult_31_104  ))
// Xd_0__inst_mult_31_108  = CARRY(( (din_a[190] & din_b[189]) ) + ( Xd_0__inst_mult_31_105  ) + ( Xd_0__inst_mult_31_104  ))
// Xd_0__inst_mult_31_109  = SHARE(GND)

	.dataa(!din_a[190]),
	.datab(!din_b[189]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_104 ),
	.sharein(Xd_0__inst_mult_31_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_107 ),
	.cout(Xd_0__inst_mult_31_108 ),
	.shareout(Xd_0__inst_mult_31_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_33 (
// Equation(s):
// Xd_0__inst_mult_31_111  = SUM(( GND ) + ( Xd_0__inst_mult_31_109  ) + ( Xd_0__inst_mult_31_108  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_31_108 ),
	.sharein(Xd_0__inst_mult_31_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_31_111 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_22_29 (
// Equation(s):
// Xd_0__inst_mult_22_95  = SUM(( GND ) + ( Xd_0__inst_mult_22_117  ) + ( Xd_0__inst_mult_22_116  ))
// Xd_0__inst_mult_22_96  = CARRY(( GND ) + ( Xd_0__inst_mult_22_117  ) + ( Xd_0__inst_mult_22_116  ))
// Xd_0__inst_mult_22_97  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_116 ),
	.sharein(Xd_0__inst_mult_22_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_95 ),
	.cout(Xd_0__inst_mult_22_96 ),
	.shareout(Xd_0__inst_mult_22_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_26 (
// Equation(s):
// Xd_0__inst_mult_15_83  = SUM(( GND ) + ( Xd_0__inst_mult_15_113  ) + ( Xd_0__inst_mult_15_112  ))
// Xd_0__inst_mult_15_84  = CARRY(( GND ) + ( Xd_0__inst_mult_15_113  ) + ( Xd_0__inst_mult_15_112  ))
// Xd_0__inst_mult_15_85  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_112 ),
	.sharein(Xd_0__inst_mult_15_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_83 ),
	.cout(Xd_0__inst_mult_15_84 ),
	.shareout(Xd_0__inst_mult_15_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_28 (
// Equation(s):
// Xd_0__inst_mult_29_91  = SUM(( GND ) + ( Xd_0__inst_mult_29_117  ) + ( Xd_0__inst_mult_29_116  ))
// Xd_0__inst_mult_29_92  = CARRY(( GND ) + ( Xd_0__inst_mult_29_117  ) + ( Xd_0__inst_mult_29_116  ))
// Xd_0__inst_mult_29_93  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_116 ),
	.sharein(Xd_0__inst_mult_29_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_91 ),
	.cout(Xd_0__inst_mult_29_92 ),
	.shareout(Xd_0__inst_mult_29_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_29_29 (
// Equation(s):
// Xd_0__inst_mult_29_96  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_29_97  = SHARE((din_b[177] & din_a[175]))

	.dataa(!din_b[177]),
	.datab(!din_a[175]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_29_96 ),
	.shareout(Xd_0__inst_mult_29_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_28 (
// Equation(s):
// Xd_0__inst_mult_11_91  = SUM(( GND ) + ( Xd_0__inst_mult_11_117  ) + ( Xd_0__inst_mult_11_116  ))
// Xd_0__inst_mult_11_92  = CARRY(( GND ) + ( Xd_0__inst_mult_11_117  ) + ( Xd_0__inst_mult_11_116  ))
// Xd_0__inst_mult_11_93  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_116 ),
	.sharein(Xd_0__inst_mult_11_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_91 ),
	.cout(Xd_0__inst_mult_11_92 ),
	.shareout(Xd_0__inst_mult_11_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_26 (
// Equation(s):
// Xd_0__inst_mult_9_83  = SUM(( GND ) + ( Xd_0__inst_mult_9_113  ) + ( Xd_0__inst_mult_9_112  ))
// Xd_0__inst_mult_9_84  = CARRY(( GND ) + ( Xd_0__inst_mult_9_113  ) + ( Xd_0__inst_mult_9_112  ))
// Xd_0__inst_mult_9_85  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_112 ),
	.sharein(Xd_0__inst_mult_9_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_83 ),
	.cout(Xd_0__inst_mult_9_84 ),
	.shareout(Xd_0__inst_mult_9_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_31_34 (
// Equation(s):
// Xd_0__inst_mult_31_116  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_31_117  = SHARE((din_b[189] & din_a[187]))

	.dataa(!din_b[189]),
	.datab(!din_a[187]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_31_116 ),
	.shareout(Xd_0__inst_mult_31_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_24 (
// Equation(s):
// Xd_0__inst_mult_8_74  = SUM(( GND ) + ( Xd_0__inst_mult_8_108  ) + ( Xd_0__inst_mult_8_107  ))
// Xd_0__inst_mult_8_75  = CARRY(( GND ) + ( Xd_0__inst_mult_8_108  ) + ( Xd_0__inst_mult_8_107  ))
// Xd_0__inst_mult_8_76  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_107 ),
	.sharein(Xd_0__inst_mult_8_108 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_74 ),
	.cout(Xd_0__inst_mult_8_75 ),
	.shareout(Xd_0__inst_mult_8_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_26 (
// Equation(s):
// Xd_0__inst_mult_7_82  = SUM(( GND ) + ( Xd_0__inst_mult_7_108  ) + ( Xd_0__inst_mult_7_107  ))
// Xd_0__inst_mult_7_83  = CARRY(( GND ) + ( Xd_0__inst_mult_7_108  ) + ( Xd_0__inst_mult_7_107  ))
// Xd_0__inst_mult_7_84  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_107 ),
	.sharein(Xd_0__inst_mult_7_108 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_82 ),
	.cout(Xd_0__inst_mult_7_83 ),
	.shareout(Xd_0__inst_mult_7_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_26 (
// Equation(s):
// Xd_0__inst_mult_2_82  = SUM(( GND ) + ( Xd_0__inst_mult_2_108  ) + ( Xd_0__inst_mult_2_107  ))
// Xd_0__inst_mult_2_83  = CARRY(( GND ) + ( Xd_0__inst_mult_2_108  ) + ( Xd_0__inst_mult_2_107  ))
// Xd_0__inst_mult_2_84  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_107 ),
	.sharein(Xd_0__inst_mult_2_108 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_82 ),
	.cout(Xd_0__inst_mult_2_83 ),
	.shareout(Xd_0__inst_mult_2_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_26 (
// Equation(s):
// Xd_0__inst_mult_0_82  = SUM(( GND ) + ( Xd_0__inst_mult_0_108  ) + ( Xd_0__inst_mult_0_107  ))
// Xd_0__inst_mult_0_83  = CARRY(( GND ) + ( Xd_0__inst_mult_0_108  ) + ( Xd_0__inst_mult_0_107  ))
// Xd_0__inst_mult_0_84  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_107 ),
	.sharein(Xd_0__inst_mult_0_108 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_82 ),
	.cout(Xd_0__inst_mult_0_83 ),
	.shareout(Xd_0__inst_mult_0_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_11_29 (
// Equation(s):
// Xd_0__inst_mult_11_96  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_11_97  = SHARE((din_b[69] & din_a[67]))

	.dataa(!din_b[69]),
	.datab(!din_a[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_11_96 ),
	.shareout(Xd_0__inst_mult_11_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_26 (
// Equation(s):
// Xd_0__inst_mult_21_83  = SUM(( GND ) + ( Xd_0__inst_mult_21_113  ) + ( Xd_0__inst_mult_21_112  ))
// Xd_0__inst_mult_21_84  = CARRY(( GND ) + ( Xd_0__inst_mult_21_113  ) + ( Xd_0__inst_mult_21_112  ))
// Xd_0__inst_mult_21_85  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_112 ),
	.sharein(Xd_0__inst_mult_21_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_83 ),
	.cout(Xd_0__inst_mult_21_84 ),
	.shareout(Xd_0__inst_mult_21_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_26_29 (
// Equation(s):
// Xd_0__inst_mult_26_95  = SUM(( GND ) + ( Xd_0__inst_mult_26_117  ) + ( Xd_0__inst_mult_26_116  ))
// Xd_0__inst_mult_26_96  = CARRY(( GND ) + ( Xd_0__inst_mult_26_117  ) + ( Xd_0__inst_mult_26_116  ))
// Xd_0__inst_mult_26_97  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_116 ),
	.sharein(Xd_0__inst_mult_26_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_95 ),
	.cout(Xd_0__inst_mult_26_96 ),
	.shareout(Xd_0__inst_mult_26_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_24_29 (
// Equation(s):
// Xd_0__inst_mult_24_95  = SUM(( GND ) + ( Xd_0__inst_mult_24_117  ) + ( Xd_0__inst_mult_24_116  ))
// Xd_0__inst_mult_24_96  = CARRY(( GND ) + ( Xd_0__inst_mult_24_117  ) + ( Xd_0__inst_mult_24_116  ))
// Xd_0__inst_mult_24_97  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_116 ),
	.sharein(Xd_0__inst_mult_24_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_95 ),
	.cout(Xd_0__inst_mult_24_96 ),
	.shareout(Xd_0__inst_mult_24_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_28 (
// Equation(s):
// Xd_0__inst_mult_25_92  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_25_93  = SHARE((din_b[153] & din_a[151]))

	.dataa(!din_b[153]),
	.datab(!din_a[151]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_25_92 ),
	.shareout(Xd_0__inst_mult_25_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_19_29 (
// Equation(s):
// Xd_0__inst_mult_19_95  = SUM(( GND ) + ( Xd_0__inst_mult_19_117  ) + ( Xd_0__inst_mult_19_116  ))
// Xd_0__inst_mult_19_96  = CARRY(( GND ) + ( Xd_0__inst_mult_19_117  ) + ( Xd_0__inst_mult_19_116  ))
// Xd_0__inst_mult_19_97  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_116 ),
	.sharein(Xd_0__inst_mult_19_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_95 ),
	.cout(Xd_0__inst_mult_19_96 ),
	.shareout(Xd_0__inst_mult_19_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_26 (
// Equation(s):
// Xd_0__inst_mult_17_83  = SUM(( GND ) + ( Xd_0__inst_mult_17_113  ) + ( Xd_0__inst_mult_17_112  ))
// Xd_0__inst_mult_17_84  = CARRY(( GND ) + ( Xd_0__inst_mult_17_113  ) + ( Xd_0__inst_mult_17_112  ))
// Xd_0__inst_mult_17_85  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_112 ),
	.sharein(Xd_0__inst_mult_17_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_83 ),
	.cout(Xd_0__inst_mult_17_84 ),
	.shareout(Xd_0__inst_mult_17_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_24 (
// Equation(s):
// Xd_0__inst_mult_12_74  = SUM(( GND ) + ( Xd_0__inst_mult_12_108  ) + ( Xd_0__inst_mult_12_107  ))
// Xd_0__inst_mult_12_75  = CARRY(( GND ) + ( Xd_0__inst_mult_12_108  ) + ( Xd_0__inst_mult_12_107  ))
// Xd_0__inst_mult_12_76  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_107 ),
	.sharein(Xd_0__inst_mult_12_108 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_74 ),
	.cout(Xd_0__inst_mult_12_75 ),
	.shareout(Xd_0__inst_mult_12_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_28 (
// Equation(s):
// Xd_0__inst_mult_27_92  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_27_93  = SHARE((din_b[165] & din_a[163]))

	.dataa(!din_b[165]),
	.datab(!din_a[163]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_27_92 ),
	.shareout(Xd_0__inst_mult_27_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_24 (
// Equation(s):
// Xd_0__inst_mult_16_74  = SUM(( (!din_a[97] & (((din_a[98] & din_b[97])))) # (din_a[97] & (!din_b[98] $ (((!din_a[98]) # (!din_b[97]))))) ) + ( Xd_0__inst_mult_16_68  ) + ( Xd_0__inst_mult_16_67  ))
// Xd_0__inst_mult_16_75  = CARRY(( (!din_a[97] & (((din_a[98] & din_b[97])))) # (din_a[97] & (!din_b[98] $ (((!din_a[98]) # (!din_b[97]))))) ) + ( Xd_0__inst_mult_16_68  ) + ( Xd_0__inst_mult_16_67  ))
// Xd_0__inst_mult_16_76  = SHARE((din_a[97] & (din_b[98] & (din_a[98] & din_b[97]))))

	.dataa(!din_a[97]),
	.datab(!din_b[98]),
	.datac(!din_a[98]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_67 ),
	.sharein(Xd_0__inst_mult_16_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_74 ),
	.cout(Xd_0__inst_mult_16_75 ),
	.shareout(Xd_0__inst_mult_16_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_25 (
// Equation(s):
// Xd_0__inst_mult_16_78  = SUM(( GND ) + ( Xd_0__inst_mult_7_96  ) + ( Xd_0__inst_mult_7_95  ))
// Xd_0__inst_mult_16_79  = CARRY(( GND ) + ( Xd_0__inst_mult_7_96  ) + ( Xd_0__inst_mult_7_95  ))
// Xd_0__inst_mult_16_80  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_16_0_q ),
	.datab(!Xd_0__inst_mult_16_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_95 ),
	.sharein(Xd_0__inst_mult_7_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_78 ),
	.cout(Xd_0__inst_mult_16_79 ),
	.shareout(Xd_0__inst_mult_16_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_27 (
// Equation(s):
// Xd_0__inst_mult_17_87  = SUM(( (!din_a[103] & (((din_a[104] & din_b[103])))) # (din_a[103] & (!din_b[104] $ (((!din_a[104]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_17_77  ) + ( Xd_0__inst_mult_17_76  ))
// Xd_0__inst_mult_17_88  = CARRY(( (!din_a[103] & (((din_a[104] & din_b[103])))) # (din_a[103] & (!din_b[104] $ (((!din_a[104]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_17_77  ) + ( Xd_0__inst_mult_17_76  ))
// Xd_0__inst_mult_17_89  = SHARE((din_a[103] & (din_b[104] & (din_a[104] & din_b[103]))))

	.dataa(!din_a[103]),
	.datab(!din_b[104]),
	.datac(!din_a[104]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_76 ),
	.sharein(Xd_0__inst_mult_17_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_87 ),
	.cout(Xd_0__inst_mult_17_88 ),
	.shareout(Xd_0__inst_mult_17_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_24 (
// Equation(s):
// Xd_0__inst_mult_14_74  = SUM(( (!din_a[85] & (((din_a[86] & din_b[85])))) # (din_a[85] & (!din_b[86] $ (((!din_a[86]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_14_68  ) + ( Xd_0__inst_mult_14_67  ))
// Xd_0__inst_mult_14_75  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[85])))) # (din_a[85] & (!din_b[86] $ (((!din_a[86]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_14_68  ) + ( Xd_0__inst_mult_14_67  ))
// Xd_0__inst_mult_14_76  = SHARE((din_a[85] & (din_b[86] & (din_a[86] & din_b[85]))))

	.dataa(!din_a[85]),
	.datab(!din_b[86]),
	.datac(!din_a[86]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_67 ),
	.sharein(Xd_0__inst_mult_14_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_74 ),
	.cout(Xd_0__inst_mult_14_75 ),
	.shareout(Xd_0__inst_mult_14_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_25 (
// Equation(s):
// Xd_0__inst_mult_14_78  = SUM(( GND ) + ( Xd_0__inst_mult_4_87  ) + ( Xd_0__inst_mult_4_86  ))
// Xd_0__inst_mult_14_79  = CARRY(( GND ) + ( Xd_0__inst_mult_4_87  ) + ( Xd_0__inst_mult_4_86  ))
// Xd_0__inst_mult_14_80  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_14_0_q ),
	.datab(!Xd_0__inst_mult_14_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_86 ),
	.sharein(Xd_0__inst_mult_4_87 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_78 ),
	.cout(Xd_0__inst_mult_14_79 ),
	.shareout(Xd_0__inst_mult_14_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_27 (
// Equation(s):
// Xd_0__inst_mult_15_87  = SUM(( (!din_a[91] & (((din_a[92] & din_b[91])))) # (din_a[91] & (!din_b[92] $ (((!din_a[92]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_15_77  ) + ( Xd_0__inst_mult_15_76  ))
// Xd_0__inst_mult_15_88  = CARRY(( (!din_a[91] & (((din_a[92] & din_b[91])))) # (din_a[91] & (!din_b[92] $ (((!din_a[92]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_15_77  ) + ( Xd_0__inst_mult_15_76  ))
// Xd_0__inst_mult_15_89  = SHARE((din_a[91] & (din_b[92] & (din_a[92] & din_b[91]))))

	.dataa(!din_a[91]),
	.datab(!din_b[92]),
	.datac(!din_a[92]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_76 ),
	.sharein(Xd_0__inst_mult_15_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_87 ),
	.cout(Xd_0__inst_mult_15_88 ),
	.shareout(Xd_0__inst_mult_15_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_25 (
// Equation(s):
// Xd_0__inst_mult_12_78  = SUM(( (!din_a[73] & (((din_a[74] & din_b[73])))) # (din_a[73] & (!din_b[74] $ (((!din_a[74]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_12_68  ) + ( Xd_0__inst_mult_12_67  ))
// Xd_0__inst_mult_12_79  = CARRY(( (!din_a[73] & (((din_a[74] & din_b[73])))) # (din_a[73] & (!din_b[74] $ (((!din_a[74]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_12_68  ) + ( Xd_0__inst_mult_12_67  ))
// Xd_0__inst_mult_12_80  = SHARE((din_a[73] & (din_b[74] & (din_a[74] & din_b[73]))))

	.dataa(!din_a[73]),
	.datab(!din_b[74]),
	.datac(!din_a[74]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_67 ),
	.sharein(Xd_0__inst_mult_12_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_78 ),
	.cout(Xd_0__inst_mult_12_79 ),
	.shareout(Xd_0__inst_mult_12_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_26 (
// Equation(s):
// Xd_0__inst_mult_12_82  = SUM(( GND ) + ( Xd_0__inst_mult_5_92  ) + ( Xd_0__inst_mult_5_91  ))
// Xd_0__inst_mult_12_83  = CARRY(( GND ) + ( Xd_0__inst_mult_5_92  ) + ( Xd_0__inst_mult_5_91  ))
// Xd_0__inst_mult_12_84  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_12_0_q ),
	.datab(!Xd_0__inst_mult_12_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_91 ),
	.sharein(Xd_0__inst_mult_5_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_82 ),
	.cout(Xd_0__inst_mult_12_83 ),
	.shareout(Xd_0__inst_mult_12_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_26 (
// Equation(s):
// Xd_0__inst_mult_13_83  = SUM(( (!din_a[79] & (((din_a[80] & din_b[79])))) # (din_a[79] & (!din_b[80] $ (((!din_a[80]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_13_77  ) + ( Xd_0__inst_mult_13_76  ))
// Xd_0__inst_mult_13_84  = CARRY(( (!din_a[79] & (((din_a[80] & din_b[79])))) # (din_a[79] & (!din_b[80] $ (((!din_a[80]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_13_77  ) + ( Xd_0__inst_mult_13_76  ))
// Xd_0__inst_mult_13_85  = SHARE((din_a[79] & (din_b[80] & (din_a[80] & din_b[79]))))

	.dataa(!din_a[79]),
	.datab(!din_b[80]),
	.datac(!din_a[80]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_76 ),
	.sharein(Xd_0__inst_mult_13_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_83 ),
	.cout(Xd_0__inst_mult_13_84 ),
	.shareout(Xd_0__inst_mult_13_85 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_24 (
// Equation(s):
// Xd_0__inst_mult_10_74  = SUM(( (!din_a[61] & (((din_a[62] & din_b[61])))) # (din_a[61] & (!din_b[62] $ (((!din_a[62]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_10_68  ) + ( Xd_0__inst_mult_10_67  ))
// Xd_0__inst_mult_10_75  = CARRY(( (!din_a[61] & (((din_a[62] & din_b[61])))) # (din_a[61] & (!din_b[62] $ (((!din_a[62]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_10_68  ) + ( Xd_0__inst_mult_10_67  ))
// Xd_0__inst_mult_10_76  = SHARE((din_a[61] & (din_b[62] & (din_a[62] & din_b[61]))))

	.dataa(!din_a[61]),
	.datab(!din_b[62]),
	.datac(!din_a[62]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_67 ),
	.sharein(Xd_0__inst_mult_10_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_74 ),
	.cout(Xd_0__inst_mult_10_75 ),
	.shareout(Xd_0__inst_mult_10_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_25 (
// Equation(s):
// Xd_0__inst_mult_10_78  = SUM(( GND ) + ( Xd_0__inst_mult_2_96  ) + ( Xd_0__inst_mult_2_95  ))
// Xd_0__inst_mult_10_79  = CARRY(( GND ) + ( Xd_0__inst_mult_2_96  ) + ( Xd_0__inst_mult_2_95  ))
// Xd_0__inst_mult_10_80  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_10_0_q ),
	.datab(!Xd_0__inst_mult_10_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_95 ),
	.sharein(Xd_0__inst_mult_2_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_78 ),
	.cout(Xd_0__inst_mult_10_79 ),
	.shareout(Xd_0__inst_mult_10_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_30 (
// Equation(s):
// Xd_0__inst_mult_11_99  = SUM(( (!din_a[67] & (((din_a[68] & din_b[67])))) # (din_a[67] & (!din_b[68] $ (((!din_a[68]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_11_85  ) + ( Xd_0__inst_mult_11_84  ))
// Xd_0__inst_mult_11_100  = CARRY(( (!din_a[67] & (((din_a[68] & din_b[67])))) # (din_a[67] & (!din_b[68] $ (((!din_a[68]) # (!din_b[67]))))) ) + ( Xd_0__inst_mult_11_85  ) + ( Xd_0__inst_mult_11_84  ))
// Xd_0__inst_mult_11_101  = SHARE((din_a[67] & (din_b[68] & (din_a[68] & din_b[67]))))

	.dataa(!din_a[67]),
	.datab(!din_b[68]),
	.datac(!din_a[68]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_84 ),
	.sharein(Xd_0__inst_mult_11_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_99 ),
	.cout(Xd_0__inst_mult_11_100 ),
	.shareout(Xd_0__inst_mult_11_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_25 (
// Equation(s):
// Xd_0__inst_mult_8_78  = SUM(( (!din_a[49] & (((din_a[50] & din_b[49])))) # (din_a[49] & (!din_b[50] $ (((!din_a[50]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_8_68  ) + ( Xd_0__inst_mult_8_67  ))
// Xd_0__inst_mult_8_79  = CARRY(( (!din_a[49] & (((din_a[50] & din_b[49])))) # (din_a[49] & (!din_b[50] $ (((!din_a[50]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_8_68  ) + ( Xd_0__inst_mult_8_67  ))
// Xd_0__inst_mult_8_80  = SHARE((din_a[49] & (din_b[50] & (din_a[50] & din_b[49]))))

	.dataa(!din_a[49]),
	.datab(!din_b[50]),
	.datac(!din_a[50]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_67 ),
	.sharein(Xd_0__inst_mult_8_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_78 ),
	.cout(Xd_0__inst_mult_8_79 ),
	.shareout(Xd_0__inst_mult_8_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_26 (
// Equation(s):
// Xd_0__inst_mult_8_82  = SUM(( GND ) + ( Xd_0__inst_mult_3_92  ) + ( Xd_0__inst_mult_3_91  ))
// Xd_0__inst_mult_8_83  = CARRY(( GND ) + ( Xd_0__inst_mult_3_92  ) + ( Xd_0__inst_mult_3_91  ))
// Xd_0__inst_mult_8_84  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_8_0_q ),
	.datab(!Xd_0__inst_mult_8_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_91 ),
	.sharein(Xd_0__inst_mult_3_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_82 ),
	.cout(Xd_0__inst_mult_8_83 ),
	.shareout(Xd_0__inst_mult_8_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_27 (
// Equation(s):
// Xd_0__inst_mult_9_87  = SUM(( (!din_a[55] & (((din_a[56] & din_b[55])))) # (din_a[55] & (!din_b[56] $ (((!din_a[56]) # (!din_b[55]))))) ) + ( Xd_0__inst_mult_9_77  ) + ( Xd_0__inst_mult_9_76  ))
// Xd_0__inst_mult_9_88  = CARRY(( (!din_a[55] & (((din_a[56] & din_b[55])))) # (din_a[55] & (!din_b[56] $ (((!din_a[56]) # (!din_b[55]))))) ) + ( Xd_0__inst_mult_9_77  ) + ( Xd_0__inst_mult_9_76  ))
// Xd_0__inst_mult_9_89  = SHARE((din_a[55] & (din_b[56] & (din_a[56] & din_b[55]))))

	.dataa(!din_a[55]),
	.datab(!din_b[56]),
	.datac(!din_a[56]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_76 ),
	.sharein(Xd_0__inst_mult_9_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_87 ),
	.cout(Xd_0__inst_mult_9_88 ),
	.shareout(Xd_0__inst_mult_9_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_24 (
// Equation(s):
// Xd_0__inst_mult_6_73  = SUM(( (!din_a[37] & (((din_a[38] & din_b[37])))) # (din_a[37] & (!din_b[38] $ (((!din_a[38]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_6_67  ) + ( Xd_0__inst_mult_6_66  ))
// Xd_0__inst_mult_6_74  = CARRY(( (!din_a[37] & (((din_a[38] & din_b[37])))) # (din_a[37] & (!din_b[38] $ (((!din_a[38]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_6_67  ) + ( Xd_0__inst_mult_6_66  ))
// Xd_0__inst_mult_6_75  = SHARE((din_a[37] & (din_b[38] & (din_a[38] & din_b[37]))))

	.dataa(!din_a[37]),
	.datab(!din_b[38]),
	.datac(!din_a[38]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_66 ),
	.sharein(Xd_0__inst_mult_6_67 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_73 ),
	.cout(Xd_0__inst_mult_6_74 ),
	.shareout(Xd_0__inst_mult_6_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_25 (
// Equation(s):
// Xd_0__inst_mult_6_77  = SUM(( GND ) + ( Xd_0__inst_mult_0_96  ) + ( Xd_0__inst_mult_0_95  ))
// Xd_0__inst_mult_6_78  = CARRY(( GND ) + ( Xd_0__inst_mult_0_96  ) + ( Xd_0__inst_mult_0_95  ))
// Xd_0__inst_mult_6_79  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_95 ),
	.sharein(Xd_0__inst_mult_0_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_77 ),
	.cout(Xd_0__inst_mult_6_78 ),
	.shareout(Xd_0__inst_mult_6_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_27 (
// Equation(s):
// Xd_0__inst_mult_7_86  = SUM(( (!din_a[43] & (((din_a[44] & din_b[43])))) # (din_a[43] & (!din_b[44] $ (((!din_a[44]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_7_76  ) + ( Xd_0__inst_mult_7_75  ))
// Xd_0__inst_mult_7_87  = CARRY(( (!din_a[43] & (((din_a[44] & din_b[43])))) # (din_a[43] & (!din_b[44] $ (((!din_a[44]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_7_76  ) + ( Xd_0__inst_mult_7_75  ))
// Xd_0__inst_mult_7_88  = SHARE((din_a[43] & (din_b[44] & (din_a[44] & din_b[43]))))

	.dataa(!din_a[43]),
	.datab(!din_b[44]),
	.datac(!din_a[44]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_75 ),
	.sharein(Xd_0__inst_mult_7_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_86 ),
	.cout(Xd_0__inst_mult_7_87 ),
	.shareout(Xd_0__inst_mult_7_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_24 (
// Equation(s):
// Xd_0__inst_mult_4_73  = SUM(( (!din_a[25] & (((din_a[26] & din_b[25])))) # (din_a[25] & (!din_b[26] $ (((!din_a[26]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_4_67  ) + ( Xd_0__inst_mult_4_66  ))
// Xd_0__inst_mult_4_74  = CARRY(( (!din_a[25] & (((din_a[26] & din_b[25])))) # (din_a[25] & (!din_b[26] $ (((!din_a[26]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_4_67  ) + ( Xd_0__inst_mult_4_66  ))
// Xd_0__inst_mult_4_75  = SHARE((din_a[25] & (din_b[26] & (din_a[26] & din_b[25]))))

	.dataa(!din_a[25]),
	.datab(!din_b[26]),
	.datac(!din_a[26]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_66 ),
	.sharein(Xd_0__inst_mult_4_67 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_73 ),
	.cout(Xd_0__inst_mult_4_74 ),
	.shareout(Xd_0__inst_mult_4_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_25 (
// Equation(s):
// Xd_0__inst_mult_4_77  = SUM(( GND ) + ( Xd_0__inst_mult_1_92  ) + ( Xd_0__inst_mult_1_91  ))
// Xd_0__inst_mult_4_78  = CARRY(( GND ) + ( Xd_0__inst_mult_1_92  ) + ( Xd_0__inst_mult_1_91  ))
// Xd_0__inst_mult_4_79  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_91 ),
	.sharein(Xd_0__inst_mult_1_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_77 ),
	.cout(Xd_0__inst_mult_4_78 ),
	.shareout(Xd_0__inst_mult_4_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_26 (
// Equation(s):
// Xd_0__inst_mult_5_82  = SUM(( (!din_a[31] & (((din_a[32] & din_b[31])))) # (din_a[31] & (!din_b[32] $ (((!din_a[32]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_5_76  ) + ( Xd_0__inst_mult_5_75  ))
// Xd_0__inst_mult_5_83  = CARRY(( (!din_a[31] & (((din_a[32] & din_b[31])))) # (din_a[31] & (!din_b[32] $ (((!din_a[32]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_5_76  ) + ( Xd_0__inst_mult_5_75  ))
// Xd_0__inst_mult_5_84  = SHARE((din_a[31] & (din_b[32] & (din_a[32] & din_b[31]))))

	.dataa(!din_a[31]),
	.datab(!din_b[32]),
	.datac(!din_a[32]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_75 ),
	.sharein(Xd_0__inst_mult_5_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_82 ),
	.cout(Xd_0__inst_mult_5_83 ),
	.shareout(Xd_0__inst_mult_5_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_27 (
// Equation(s):
// Xd_0__inst_mult_2_86  = SUM(( (!din_a[13] & (((din_a[14] & din_b[13])))) # (din_a[13] & (!din_b[14] $ (((!din_a[14]) # (!din_b[13]))))) ) + ( Xd_0__inst_mult_2_76  ) + ( Xd_0__inst_mult_2_75  ))
// Xd_0__inst_mult_2_87  = CARRY(( (!din_a[13] & (((din_a[14] & din_b[13])))) # (din_a[13] & (!din_b[14] $ (((!din_a[14]) # (!din_b[13]))))) ) + ( Xd_0__inst_mult_2_76  ) + ( Xd_0__inst_mult_2_75  ))
// Xd_0__inst_mult_2_88  = SHARE((din_a[13] & (din_b[14] & (din_a[14] & din_b[13]))))

	.dataa(!din_a[13]),
	.datab(!din_b[14]),
	.datac(!din_a[14]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_75 ),
	.sharein(Xd_0__inst_mult_2_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_86 ),
	.cout(Xd_0__inst_mult_2_87 ),
	.shareout(Xd_0__inst_mult_2_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_26 (
// Equation(s):
// Xd_0__inst_mult_3_82  = SUM(( (!din_a[19] & (((din_a[20] & din_b[19])))) # (din_a[19] & (!din_b[20] $ (((!din_a[20]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_3_76  ) + ( Xd_0__inst_mult_3_75  ))
// Xd_0__inst_mult_3_83  = CARRY(( (!din_a[19] & (((din_a[20] & din_b[19])))) # (din_a[19] & (!din_b[20] $ (((!din_a[20]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_3_76  ) + ( Xd_0__inst_mult_3_75  ))
// Xd_0__inst_mult_3_84  = SHARE((din_a[19] & (din_b[20] & (din_a[20] & din_b[19]))))

	.dataa(!din_a[19]),
	.datab(!din_b[20]),
	.datac(!din_a[20]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_75 ),
	.sharein(Xd_0__inst_mult_3_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_82 ),
	.cout(Xd_0__inst_mult_3_83 ),
	.shareout(Xd_0__inst_mult_3_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_27 (
// Equation(s):
// Xd_0__inst_mult_0_86  = SUM(( (!din_a[1] & (((din_a[2] & din_b[1])))) # (din_a[1] & (!din_b[2] $ (((!din_a[2]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_76  ) + ( Xd_0__inst_mult_0_75  ))
// Xd_0__inst_mult_0_87  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[1])))) # (din_a[1] & (!din_b[2] $ (((!din_a[2]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_76  ) + ( Xd_0__inst_mult_0_75  ))
// Xd_0__inst_mult_0_88  = SHARE((din_a[1] & (din_b[2] & (din_a[2] & din_b[1]))))

	.dataa(!din_a[1]),
	.datab(!din_b[2]),
	.datac(!din_a[2]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_75 ),
	.sharein(Xd_0__inst_mult_0_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_86 ),
	.cout(Xd_0__inst_mult_0_87 ),
	.shareout(Xd_0__inst_mult_0_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_26 (
// Equation(s):
// Xd_0__inst_mult_1_82  = SUM(( (!din_a[7] & (((din_a[8] & din_b[7])))) # (din_a[7] & (!din_b[8] $ (((!din_a[8]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_76  ) + ( Xd_0__inst_mult_1_75  ))
// Xd_0__inst_mult_1_83  = CARRY(( (!din_a[7] & (((din_a[8] & din_b[7])))) # (din_a[7] & (!din_b[8] $ (((!din_a[8]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_76  ) + ( Xd_0__inst_mult_1_75  ))
// Xd_0__inst_mult_1_84  = SHARE((din_a[7] & (din_b[8] & (din_a[8] & din_b[7]))))

	.dataa(!din_a[7]),
	.datab(!din_b[8]),
	.datac(!din_a[8]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_75 ),
	.sharein(Xd_0__inst_mult_1_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_82 ),
	.cout(Xd_0__inst_mult_1_83 ),
	.shareout(Xd_0__inst_mult_1_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_29 (
// Equation(s):
// Xd_0__inst_mult_28_95  = SUM(( (!din_a[169] & (((din_a[170] & din_b[169])))) # (din_a[169] & (!din_b[170] $ (((!din_a[170]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_28_89  ) + ( Xd_0__inst_mult_28_88  ))
// Xd_0__inst_mult_28_96  = CARRY(( (!din_a[169] & (((din_a[170] & din_b[169])))) # (din_a[169] & (!din_b[170] $ (((!din_a[170]) # (!din_b[169]))))) ) + ( Xd_0__inst_mult_28_89  ) + ( Xd_0__inst_mult_28_88  ))
// Xd_0__inst_mult_28_97  = SHARE((din_a[169] & (din_b[170] & (din_a[170] & din_b[169]))))

	.dataa(!din_a[169]),
	.datab(!din_b[170]),
	.datac(!din_a[170]),
	.datad(!din_b[169]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_88 ),
	.sharein(Xd_0__inst_mult_28_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_95 ),
	.cout(Xd_0__inst_mult_28_96 ),
	.shareout(Xd_0__inst_mult_28_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_30 (
// Equation(s):
// Xd_0__inst_mult_29_99  = SUM(( (!din_a[175] & (((din_a[176] & din_b[175])))) # (din_a[175] & (!din_b[176] $ (((!din_a[176]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_29_85  ) + ( Xd_0__inst_mult_29_84  ))
// Xd_0__inst_mult_29_100  = CARRY(( (!din_a[175] & (((din_a[176] & din_b[175])))) # (din_a[175] & (!din_b[176] $ (((!din_a[176]) # (!din_b[175]))))) ) + ( Xd_0__inst_mult_29_85  ) + ( Xd_0__inst_mult_29_84  ))
// Xd_0__inst_mult_29_101  = SHARE((din_a[175] & (din_b[176] & (din_a[176] & din_b[175]))))

	.dataa(!din_a[175]),
	.datab(!din_b[176]),
	.datac(!din_a[176]),
	.datad(!din_b[175]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_84 ),
	.sharein(Xd_0__inst_mult_29_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_99 ),
	.cout(Xd_0__inst_mult_29_100 ),
	.shareout(Xd_0__inst_mult_29_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_30 (
// Equation(s):
// Xd_0__inst_mult_26_99  = SUM(( (!din_a[157] & (((din_a[158] & din_b[157])))) # (din_a[157] & (!din_b[158] $ (((!din_a[158]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_26_89  ) + ( Xd_0__inst_mult_26_88  ))
// Xd_0__inst_mult_26_100  = CARRY(( (!din_a[157] & (((din_a[158] & din_b[157])))) # (din_a[157] & (!din_b[158] $ (((!din_a[158]) # (!din_b[157]))))) ) + ( Xd_0__inst_mult_26_89  ) + ( Xd_0__inst_mult_26_88  ))
// Xd_0__inst_mult_26_101  = SHARE((din_a[157] & (din_b[158] & (din_a[158] & din_b[157]))))

	.dataa(!din_a[157]),
	.datab(!din_b[158]),
	.datac(!din_a[158]),
	.datad(!din_b[157]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_88 ),
	.sharein(Xd_0__inst_mult_26_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_99 ),
	.cout(Xd_0__inst_mult_26_100 ),
	.shareout(Xd_0__inst_mult_26_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_29 (
// Equation(s):
// Xd_0__inst_mult_27_95  = SUM(( (!din_a[163] & (((din_a[164] & din_b[163])))) # (din_a[163] & (!din_b[164] $ (((!din_a[164]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_27_85  ) + ( Xd_0__inst_mult_27_84  ))
// Xd_0__inst_mult_27_96  = CARRY(( (!din_a[163] & (((din_a[164] & din_b[163])))) # (din_a[163] & (!din_b[164] $ (((!din_a[164]) # (!din_b[163]))))) ) + ( Xd_0__inst_mult_27_85  ) + ( Xd_0__inst_mult_27_84  ))
// Xd_0__inst_mult_27_97  = SHARE((din_a[163] & (din_b[164] & (din_a[164] & din_b[163]))))

	.dataa(!din_a[163]),
	.datab(!din_b[164]),
	.datac(!din_a[164]),
	.datad(!din_b[163]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_84 ),
	.sharein(Xd_0__inst_mult_27_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_95 ),
	.cout(Xd_0__inst_mult_27_96 ),
	.shareout(Xd_0__inst_mult_27_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_30 (
// Equation(s):
// Xd_0__inst_mult_24_99  = SUM(( (!din_a[145] & (((din_a[146] & din_b[145])))) # (din_a[145] & (!din_b[146] $ (((!din_a[146]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_24_89  ) + ( Xd_0__inst_mult_24_88  ))
// Xd_0__inst_mult_24_100  = CARRY(( (!din_a[145] & (((din_a[146] & din_b[145])))) # (din_a[145] & (!din_b[146] $ (((!din_a[146]) # (!din_b[145]))))) ) + ( Xd_0__inst_mult_24_89  ) + ( Xd_0__inst_mult_24_88  ))
// Xd_0__inst_mult_24_101  = SHARE((din_a[145] & (din_b[146] & (din_a[146] & din_b[145]))))

	.dataa(!din_a[145]),
	.datab(!din_b[146]),
	.datac(!din_a[146]),
	.datad(!din_b[145]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_88 ),
	.sharein(Xd_0__inst_mult_24_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_99 ),
	.cout(Xd_0__inst_mult_24_100 ),
	.shareout(Xd_0__inst_mult_24_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_29 (
// Equation(s):
// Xd_0__inst_mult_25_95  = SUM(( (!din_a[151] & (((din_a[152] & din_b[151])))) # (din_a[151] & (!din_b[152] $ (((!din_a[152]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_25_85  ) + ( Xd_0__inst_mult_25_84  ))
// Xd_0__inst_mult_25_96  = CARRY(( (!din_a[151] & (((din_a[152] & din_b[151])))) # (din_a[151] & (!din_b[152] $ (((!din_a[152]) # (!din_b[151]))))) ) + ( Xd_0__inst_mult_25_85  ) + ( Xd_0__inst_mult_25_84  ))
// Xd_0__inst_mult_25_97  = SHARE((din_a[151] & (din_b[152] & (din_a[152] & din_b[151]))))

	.dataa(!din_a[151]),
	.datab(!din_b[152]),
	.datac(!din_a[152]),
	.datad(!din_b[151]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_84 ),
	.sharein(Xd_0__inst_mult_25_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_95 ),
	.cout(Xd_0__inst_mult_25_96 ),
	.shareout(Xd_0__inst_mult_25_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_30 (
// Equation(s):
// Xd_0__inst_mult_22_99  = SUM(( (!din_a[133] & (((din_a[134] & din_b[133])))) # (din_a[133] & (!din_b[134] $ (((!din_a[134]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_22_89  ) + ( Xd_0__inst_mult_22_88  ))
// Xd_0__inst_mult_22_100  = CARRY(( (!din_a[133] & (((din_a[134] & din_b[133])))) # (din_a[133] & (!din_b[134] $ (((!din_a[134]) # (!din_b[133]))))) ) + ( Xd_0__inst_mult_22_89  ) + ( Xd_0__inst_mult_22_88  ))
// Xd_0__inst_mult_22_101  = SHARE((din_a[133] & (din_b[134] & (din_a[134] & din_b[133]))))

	.dataa(!din_a[133]),
	.datab(!din_b[134]),
	.datac(!din_a[134]),
	.datad(!din_b[133]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_88 ),
	.sharein(Xd_0__inst_mult_22_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_99 ),
	.cout(Xd_0__inst_mult_22_100 ),
	.shareout(Xd_0__inst_mult_22_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_29 (
// Equation(s):
// Xd_0__inst_mult_23_95  = SUM(( (!din_a[139] & (((din_a[140] & din_b[139])))) # (din_a[139] & (!din_b[140] $ (((!din_a[140]) # (!din_b[139]))))) ) + ( Xd_0__inst_mult_23_89  ) + ( Xd_0__inst_mult_23_88  ))
// Xd_0__inst_mult_23_96  = CARRY(( (!din_a[139] & (((din_a[140] & din_b[139])))) # (din_a[139] & (!din_b[140] $ (((!din_a[140]) # (!din_b[139]))))) ) + ( Xd_0__inst_mult_23_89  ) + ( Xd_0__inst_mult_23_88  ))
// Xd_0__inst_mult_23_97  = SHARE((din_a[139] & (din_b[140] & (din_a[140] & din_b[139]))))

	.dataa(!din_a[139]),
	.datab(!din_b[140]),
	.datac(!din_a[140]),
	.datad(!din_b[139]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_88 ),
	.sharein(Xd_0__inst_mult_23_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_95 ),
	.cout(Xd_0__inst_mult_23_96 ),
	.shareout(Xd_0__inst_mult_23_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_29 (
// Equation(s):
// Xd_0__inst_mult_20_95  = SUM(( (!din_a[121] & (((din_a[122] & din_b[121])))) # (din_a[121] & (!din_b[122] $ (((!din_a[122]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_20_89  ) + ( Xd_0__inst_mult_20_88  ))
// Xd_0__inst_mult_20_96  = CARRY(( (!din_a[121] & (((din_a[122] & din_b[121])))) # (din_a[121] & (!din_b[122] $ (((!din_a[122]) # (!din_b[121]))))) ) + ( Xd_0__inst_mult_20_89  ) + ( Xd_0__inst_mult_20_88  ))
// Xd_0__inst_mult_20_97  = SHARE((din_a[121] & (din_b[122] & (din_a[122] & din_b[121]))))

	.dataa(!din_a[121]),
	.datab(!din_b[122]),
	.datac(!din_a[122]),
	.datad(!din_b[121]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_88 ),
	.sharein(Xd_0__inst_mult_20_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_95 ),
	.cout(Xd_0__inst_mult_20_96 ),
	.shareout(Xd_0__inst_mult_20_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_27 (
// Equation(s):
// Xd_0__inst_mult_21_87  = SUM(( (!din_a[127] & (((din_a[128] & din_b[127])))) # (din_a[127] & (!din_b[128] $ (((!din_a[128]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_21_77  ) + ( Xd_0__inst_mult_21_76  ))
// Xd_0__inst_mult_21_88  = CARRY(( (!din_a[127] & (((din_a[128] & din_b[127])))) # (din_a[127] & (!din_b[128] $ (((!din_a[128]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_21_77  ) + ( Xd_0__inst_mult_21_76  ))
// Xd_0__inst_mult_21_89  = SHARE((din_a[127] & (din_b[128] & (din_a[128] & din_b[127]))))

	.dataa(!din_a[127]),
	.datab(!din_b[128]),
	.datac(!din_a[128]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_76 ),
	.sharein(Xd_0__inst_mult_21_77 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_87 ),
	.cout(Xd_0__inst_mult_21_88 ),
	.shareout(Xd_0__inst_mult_21_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_24 (
// Equation(s):
// Xd_0__inst_mult_18_74  = SUM(( (!din_a[109] & (((din_a[110] & din_b[109])))) # (din_a[109] & (!din_b[110] $ (((!din_a[110]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_18_68  ) + ( Xd_0__inst_mult_18_67  ))
// Xd_0__inst_mult_18_75  = CARRY(( (!din_a[109] & (((din_a[110] & din_b[109])))) # (din_a[109] & (!din_b[110] $ (((!din_a[110]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_18_68  ) + ( Xd_0__inst_mult_18_67  ))
// Xd_0__inst_mult_18_76  = SHARE((din_a[109] & (din_b[110] & (din_a[110] & din_b[109]))))

	.dataa(!din_a[109]),
	.datab(!din_b[110]),
	.datac(!din_a[110]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_67 ),
	.sharein(Xd_0__inst_mult_18_68 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_74 ),
	.cout(Xd_0__inst_mult_18_75 ),
	.shareout(Xd_0__inst_mult_18_76 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_25 (
// Equation(s):
// Xd_0__inst_mult_18_78  = SUM(( GND ) + ( Xd_0__inst_mult_6_87  ) + ( Xd_0__inst_mult_6_86  ))
// Xd_0__inst_mult_18_79  = CARRY(( GND ) + ( Xd_0__inst_mult_6_87  ) + ( Xd_0__inst_mult_6_86  ))
// Xd_0__inst_mult_18_80  = SHARE(VCC)

	.dataa(!Xd_0__inst_mult_18_0_q ),
	.datab(!Xd_0__inst_mult_18_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_86 ),
	.sharein(Xd_0__inst_mult_6_87 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_78 ),
	.cout(Xd_0__inst_mult_18_79 ),
	.shareout(Xd_0__inst_mult_18_80 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_30 (
// Equation(s):
// Xd_0__inst_mult_19_99  = SUM(( (!din_a[115] & (((din_a[116] & din_b[115])))) # (din_a[115] & (!din_b[116] $ (((!din_a[116]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_19_89  ) + ( Xd_0__inst_mult_19_88  ))
// Xd_0__inst_mult_19_100  = CARRY(( (!din_a[115] & (((din_a[116] & din_b[115])))) # (din_a[115] & (!din_b[116] $ (((!din_a[116]) # (!din_b[115]))))) ) + ( Xd_0__inst_mult_19_89  ) + ( Xd_0__inst_mult_19_88  ))
// Xd_0__inst_mult_19_101  = SHARE((din_a[115] & (din_b[116] & (din_a[116] & din_b[115]))))

	.dataa(!din_a[115]),
	.datab(!din_b[116]),
	.datac(!din_a[116]),
	.datad(!din_b[115]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_88 ),
	.sharein(Xd_0__inst_mult_19_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_99 ),
	.cout(Xd_0__inst_mult_19_100 ),
	.shareout(Xd_0__inst_mult_19_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_26 (
// Equation(s):
// Xd_0__inst_mult_16_82  = SUM(( (din_a[98] & din_b[98]) ) + ( Xd_0__inst_mult_16_76  ) + ( Xd_0__inst_mult_16_75  ))
// Xd_0__inst_mult_16_83  = CARRY(( (din_a[98] & din_b[98]) ) + ( Xd_0__inst_mult_16_76  ) + ( Xd_0__inst_mult_16_75  ))
// Xd_0__inst_mult_16_84  = SHARE((din_a[98] & din_b[99]))

	.dataa(!din_a[98]),
	.datab(!din_b[98]),
	.datac(!din_b[99]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_75 ),
	.sharein(Xd_0__inst_mult_16_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_82 ),
	.cout(Xd_0__inst_mult_16_83 ),
	.shareout(Xd_0__inst_mult_16_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_27 (
// Equation(s):
// Xd_0__inst_mult_16_86  = SUM(( (!din_a[100] & (((din_a[99] & din_b[97])))) # (din_a[100] & (!din_b[96] $ (((!din_a[99]) # (!din_b[97]))))) ) + ( Xd_0__inst_mult_16_112  ) + ( Xd_0__inst_mult_16_111  ))
// Xd_0__inst_mult_16_87  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[97])))) # (din_a[100] & (!din_b[96] $ (((!din_a[99]) # (!din_b[97]))))) ) + ( Xd_0__inst_mult_16_112  ) + ( Xd_0__inst_mult_16_111  ))
// Xd_0__inst_mult_16_88  = SHARE((din_a[100] & (din_b[96] & (din_a[99] & din_b[97]))))

	.dataa(!din_a[100]),
	.datab(!din_b[96]),
	.datac(!din_a[99]),
	.datad(!din_b[97]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_111 ),
	.sharein(Xd_0__inst_mult_16_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_86 ),
	.cout(Xd_0__inst_mult_16_87 ),
	.shareout(Xd_0__inst_mult_16_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_28 (
// Equation(s):
// Xd_0__inst_mult_17_91  = SUM(( (din_a[104] & din_b[104]) ) + ( Xd_0__inst_mult_17_89  ) + ( Xd_0__inst_mult_17_88  ))
// Xd_0__inst_mult_17_92  = CARRY(( (din_a[104] & din_b[104]) ) + ( Xd_0__inst_mult_17_89  ) + ( Xd_0__inst_mult_17_88  ))
// Xd_0__inst_mult_17_93  = SHARE((din_a[104] & din_b[105]))

	.dataa(!din_a[104]),
	.datab(!din_b[104]),
	.datac(!din_b[105]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_88 ),
	.sharein(Xd_0__inst_mult_17_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_91 ),
	.cout(Xd_0__inst_mult_17_92 ),
	.shareout(Xd_0__inst_mult_17_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_29 (
// Equation(s):
// Xd_0__inst_mult_17_95  = SUM(( (!din_a[106] & (((din_a[105] & din_b[103])))) # (din_a[106] & (!din_b[102] $ (((!din_a[105]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_17_117  ) + ( Xd_0__inst_mult_17_116  ))
// Xd_0__inst_mult_17_96  = CARRY(( (!din_a[106] & (((din_a[105] & din_b[103])))) # (din_a[106] & (!din_b[102] $ (((!din_a[105]) # (!din_b[103]))))) ) + ( Xd_0__inst_mult_17_117  ) + ( Xd_0__inst_mult_17_116  ))
// Xd_0__inst_mult_17_97  = SHARE((din_a[106] & (din_b[102] & (din_a[105] & din_b[103]))))

	.dataa(!din_a[106]),
	.datab(!din_b[102]),
	.datac(!din_a[105]),
	.datad(!din_b[103]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_116 ),
	.sharein(Xd_0__inst_mult_17_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_95 ),
	.cout(Xd_0__inst_mult_17_96 ),
	.shareout(Xd_0__inst_mult_17_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_26 (
// Equation(s):
// Xd_0__inst_mult_14_82  = SUM(( (din_a[86] & din_b[86]) ) + ( Xd_0__inst_mult_14_76  ) + ( Xd_0__inst_mult_14_75  ))
// Xd_0__inst_mult_14_83  = CARRY(( (din_a[86] & din_b[86]) ) + ( Xd_0__inst_mult_14_76  ) + ( Xd_0__inst_mult_14_75  ))
// Xd_0__inst_mult_14_84  = SHARE((din_a[86] & din_b[87]))

	.dataa(!din_a[86]),
	.datab(!din_b[86]),
	.datac(!din_b[87]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_75 ),
	.sharein(Xd_0__inst_mult_14_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_82 ),
	.cout(Xd_0__inst_mult_14_83 ),
	.shareout(Xd_0__inst_mult_14_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_27 (
// Equation(s):
// Xd_0__inst_mult_14_86  = SUM(( (!din_a[88] & (((din_a[87] & din_b[85])))) # (din_a[88] & (!din_b[84] $ (((!din_a[87]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_14_112  ) + ( Xd_0__inst_mult_14_111  ))
// Xd_0__inst_mult_14_87  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[85])))) # (din_a[88] & (!din_b[84] $ (((!din_a[87]) # (!din_b[85]))))) ) + ( Xd_0__inst_mult_14_112  ) + ( Xd_0__inst_mult_14_111  ))
// Xd_0__inst_mult_14_88  = SHARE((din_a[88] & (din_b[84] & (din_a[87] & din_b[85]))))

	.dataa(!din_a[88]),
	.datab(!din_b[84]),
	.datac(!din_a[87]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_111 ),
	.sharein(Xd_0__inst_mult_14_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_86 ),
	.cout(Xd_0__inst_mult_14_87 ),
	.shareout(Xd_0__inst_mult_14_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_28 (
// Equation(s):
// Xd_0__inst_mult_15_91  = SUM(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_15_89  ) + ( Xd_0__inst_mult_15_88  ))
// Xd_0__inst_mult_15_92  = CARRY(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_15_89  ) + ( Xd_0__inst_mult_15_88  ))
// Xd_0__inst_mult_15_93  = SHARE((din_a[92] & din_b[93]))

	.dataa(!din_a[92]),
	.datab(!din_b[92]),
	.datac(!din_b[93]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_88 ),
	.sharein(Xd_0__inst_mult_15_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_91 ),
	.cout(Xd_0__inst_mult_15_92 ),
	.shareout(Xd_0__inst_mult_15_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_29 (
// Equation(s):
// Xd_0__inst_mult_15_95  = SUM(( (!din_a[94] & (((din_a[93] & din_b[91])))) # (din_a[94] & (!din_b[90] $ (((!din_a[93]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_15_117  ) + ( Xd_0__inst_mult_15_116  ))
// Xd_0__inst_mult_15_96  = CARRY(( (!din_a[94] & (((din_a[93] & din_b[91])))) # (din_a[94] & (!din_b[90] $ (((!din_a[93]) # (!din_b[91]))))) ) + ( Xd_0__inst_mult_15_117  ) + ( Xd_0__inst_mult_15_116  ))
// Xd_0__inst_mult_15_97  = SHARE((din_a[94] & (din_b[90] & (din_a[93] & din_b[91]))))

	.dataa(!din_a[94]),
	.datab(!din_b[90]),
	.datac(!din_a[93]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_116 ),
	.sharein(Xd_0__inst_mult_15_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_95 ),
	.cout(Xd_0__inst_mult_15_96 ),
	.shareout(Xd_0__inst_mult_15_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_27 (
// Equation(s):
// Xd_0__inst_mult_12_86  = SUM(( (din_a[74] & din_b[74]) ) + ( Xd_0__inst_mult_12_80  ) + ( Xd_0__inst_mult_12_79  ))
// Xd_0__inst_mult_12_87  = CARRY(( (din_a[74] & din_b[74]) ) + ( Xd_0__inst_mult_12_80  ) + ( Xd_0__inst_mult_12_79  ))
// Xd_0__inst_mult_12_88  = SHARE((din_a[74] & din_b[75]))

	.dataa(!din_a[74]),
	.datab(!din_b[74]),
	.datac(!din_b[75]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_79 ),
	.sharein(Xd_0__inst_mult_12_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_86 ),
	.cout(Xd_0__inst_mult_12_87 ),
	.shareout(Xd_0__inst_mult_12_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_28 (
// Equation(s):
// Xd_0__inst_mult_12_90  = SUM(( (!din_a[76] & (((din_a[75] & din_b[73])))) # (din_a[76] & (!din_b[72] $ (((!din_a[75]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_12_112  ) + ( Xd_0__inst_mult_12_111  ))
// Xd_0__inst_mult_12_91  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[73])))) # (din_a[76] & (!din_b[72] $ (((!din_a[75]) # (!din_b[73]))))) ) + ( Xd_0__inst_mult_12_112  ) + ( Xd_0__inst_mult_12_111  ))
// Xd_0__inst_mult_12_92  = SHARE((din_a[76] & (din_b[72] & (din_a[75] & din_b[73]))))

	.dataa(!din_a[76]),
	.datab(!din_b[72]),
	.datac(!din_a[75]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_111 ),
	.sharein(Xd_0__inst_mult_12_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_90 ),
	.cout(Xd_0__inst_mult_12_91 ),
	.shareout(Xd_0__inst_mult_12_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_27 (
// Equation(s):
// Xd_0__inst_mult_13_87  = SUM(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_13_85  ) + ( Xd_0__inst_mult_13_84  ))
// Xd_0__inst_mult_13_88  = CARRY(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_13_85  ) + ( Xd_0__inst_mult_13_84  ))
// Xd_0__inst_mult_13_89  = SHARE((din_a[80] & din_b[81]))

	.dataa(!din_a[80]),
	.datab(!din_b[80]),
	.datac(!din_b[81]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_84 ),
	.sharein(Xd_0__inst_mult_13_85 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_87 ),
	.cout(Xd_0__inst_mult_13_88 ),
	.shareout(Xd_0__inst_mult_13_89 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_28 (
// Equation(s):
// Xd_0__inst_mult_13_91  = SUM(( (!din_a[82] & (((din_a[81] & din_b[79])))) # (din_a[82] & (!din_b[78] $ (((!din_a[81]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_13_117  ) + ( Xd_0__inst_mult_13_116  ))
// Xd_0__inst_mult_13_92  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[79])))) # (din_a[82] & (!din_b[78] $ (((!din_a[81]) # (!din_b[79]))))) ) + ( Xd_0__inst_mult_13_117  ) + ( Xd_0__inst_mult_13_116  ))
// Xd_0__inst_mult_13_93  = SHARE((din_a[82] & (din_b[78] & (din_a[81] & din_b[79]))))

	.dataa(!din_a[82]),
	.datab(!din_b[78]),
	.datac(!din_a[81]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_116 ),
	.sharein(Xd_0__inst_mult_13_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_91 ),
	.cout(Xd_0__inst_mult_13_92 ),
	.shareout(Xd_0__inst_mult_13_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_26 (
// Equation(s):
// Xd_0__inst_mult_10_82  = SUM(( (din_a[62] & din_b[62]) ) + ( Xd_0__inst_mult_10_76  ) + ( Xd_0__inst_mult_10_75  ))
// Xd_0__inst_mult_10_83  = CARRY(( (din_a[62] & din_b[62]) ) + ( Xd_0__inst_mult_10_76  ) + ( Xd_0__inst_mult_10_75  ))
// Xd_0__inst_mult_10_84  = SHARE((din_a[62] & din_b[63]))

	.dataa(!din_a[62]),
	.datab(!din_b[62]),
	.datac(!din_b[63]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_75 ),
	.sharein(Xd_0__inst_mult_10_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_82 ),
	.cout(Xd_0__inst_mult_10_83 ),
	.shareout(Xd_0__inst_mult_10_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_27 (
// Equation(s):
// Xd_0__inst_mult_10_86  = SUM(( (!din_a[64] & (((din_a[63] & din_b[61])))) # (din_a[64] & (!din_b[60] $ (((!din_a[63]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_10_112  ) + ( Xd_0__inst_mult_10_111  ))
// Xd_0__inst_mult_10_87  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[61])))) # (din_a[64] & (!din_b[60] $ (((!din_a[63]) # (!din_b[61]))))) ) + ( Xd_0__inst_mult_10_112  ) + ( Xd_0__inst_mult_10_111  ))
// Xd_0__inst_mult_10_88  = SHARE((din_a[64] & (din_b[60] & (din_a[63] & din_b[61]))))

	.dataa(!din_a[64]),
	.datab(!din_b[60]),
	.datac(!din_a[63]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_111 ),
	.sharein(Xd_0__inst_mult_10_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_86 ),
	.cout(Xd_0__inst_mult_10_87 ),
	.shareout(Xd_0__inst_mult_10_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_31 (
// Equation(s):
// Xd_0__inst_mult_11_103  = SUM(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_11_101  ) + ( Xd_0__inst_mult_11_100  ))
// Xd_0__inst_mult_11_104  = CARRY(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_11_101  ) + ( Xd_0__inst_mult_11_100  ))
// Xd_0__inst_mult_11_105  = SHARE((din_a[68] & din_b[69]))

	.dataa(!din_a[68]),
	.datab(!din_b[68]),
	.datac(!din_b[69]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_100 ),
	.sharein(Xd_0__inst_mult_11_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_103 ),
	.cout(Xd_0__inst_mult_11_104 ),
	.shareout(Xd_0__inst_mult_11_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_27 (
// Equation(s):
// Xd_0__inst_mult_8_86  = SUM(( (din_a[50] & din_b[50]) ) + ( Xd_0__inst_mult_8_80  ) + ( Xd_0__inst_mult_8_79  ))
// Xd_0__inst_mult_8_87  = CARRY(( (din_a[50] & din_b[50]) ) + ( Xd_0__inst_mult_8_80  ) + ( Xd_0__inst_mult_8_79  ))
// Xd_0__inst_mult_8_88  = SHARE((din_a[50] & din_b[51]))

	.dataa(!din_a[50]),
	.datab(!din_b[50]),
	.datac(!din_b[51]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_79 ),
	.sharein(Xd_0__inst_mult_8_80 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_86 ),
	.cout(Xd_0__inst_mult_8_87 ),
	.shareout(Xd_0__inst_mult_8_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_28 (
// Equation(s):
// Xd_0__inst_mult_8_90  = SUM(( (!din_a[52] & (((din_a[51] & din_b[49])))) # (din_a[52] & (!din_b[48] $ (((!din_a[51]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_8_112  ) + ( Xd_0__inst_mult_8_111  ))
// Xd_0__inst_mult_8_91  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[49])))) # (din_a[52] & (!din_b[48] $ (((!din_a[51]) # (!din_b[49]))))) ) + ( Xd_0__inst_mult_8_112  ) + ( Xd_0__inst_mult_8_111  ))
// Xd_0__inst_mult_8_92  = SHARE((din_a[52] & (din_b[48] & (din_a[51] & din_b[49]))))

	.dataa(!din_a[52]),
	.datab(!din_b[48]),
	.datac(!din_a[51]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_111 ),
	.sharein(Xd_0__inst_mult_8_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_90 ),
	.cout(Xd_0__inst_mult_8_91 ),
	.shareout(Xd_0__inst_mult_8_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_28 (
// Equation(s):
// Xd_0__inst_mult_9_91  = SUM(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_9_89  ) + ( Xd_0__inst_mult_9_88  ))
// Xd_0__inst_mult_9_92  = CARRY(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_9_89  ) + ( Xd_0__inst_mult_9_88  ))
// Xd_0__inst_mult_9_93  = SHARE((din_a[56] & din_b[57]))

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(!din_b[57]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_88 ),
	.sharein(Xd_0__inst_mult_9_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_91 ),
	.cout(Xd_0__inst_mult_9_92 ),
	.shareout(Xd_0__inst_mult_9_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_29 (
// Equation(s):
// Xd_0__inst_mult_9_95  = SUM(( (!din_a[58] & (((din_a[57] & din_b[55])))) # (din_a[58] & (!din_b[54] $ (((!din_a[57]) # (!din_b[55]))))) ) + ( Xd_0__inst_mult_9_117  ) + ( Xd_0__inst_mult_9_116  ))
// Xd_0__inst_mult_9_96  = CARRY(( (!din_a[58] & (((din_a[57] & din_b[55])))) # (din_a[58] & (!din_b[54] $ (((!din_a[57]) # (!din_b[55]))))) ) + ( Xd_0__inst_mult_9_117  ) + ( Xd_0__inst_mult_9_116  ))
// Xd_0__inst_mult_9_97  = SHARE((din_a[58] & (din_b[54] & (din_a[57] & din_b[55]))))

	.dataa(!din_a[58]),
	.datab(!din_b[54]),
	.datac(!din_a[57]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_116 ),
	.sharein(Xd_0__inst_mult_9_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_95 ),
	.cout(Xd_0__inst_mult_9_96 ),
	.shareout(Xd_0__inst_mult_9_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_26 (
// Equation(s):
// Xd_0__inst_mult_6_81  = SUM(( (din_a[38] & din_b[38]) ) + ( Xd_0__inst_mult_6_75  ) + ( Xd_0__inst_mult_6_74  ))
// Xd_0__inst_mult_6_82  = CARRY(( (din_a[38] & din_b[38]) ) + ( Xd_0__inst_mult_6_75  ) + ( Xd_0__inst_mult_6_74  ))
// Xd_0__inst_mult_6_83  = SHARE((din_a[38] & din_b[39]))

	.dataa(!din_a[38]),
	.datab(!din_b[38]),
	.datac(!din_b[39]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_74 ),
	.sharein(Xd_0__inst_mult_6_75 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_81 ),
	.cout(Xd_0__inst_mult_6_82 ),
	.shareout(Xd_0__inst_mult_6_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_27 (
// Equation(s):
// Xd_0__inst_mult_6_85  = SUM(( (!din_a[40] & (((din_a[39] & din_b[37])))) # (din_a[40] & (!din_b[36] $ (((!din_a[39]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_6_107  ) + ( Xd_0__inst_mult_6_106  ))
// Xd_0__inst_mult_6_86  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[37])))) # (din_a[40] & (!din_b[36] $ (((!din_a[39]) # (!din_b[37]))))) ) + ( Xd_0__inst_mult_6_107  ) + ( Xd_0__inst_mult_6_106  ))
// Xd_0__inst_mult_6_87  = SHARE((din_a[40] & (din_b[36] & (din_a[39] & din_b[37]))))

	.dataa(!din_a[40]),
	.datab(!din_b[36]),
	.datac(!din_a[39]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_106 ),
	.sharein(Xd_0__inst_mult_6_107 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_85 ),
	.cout(Xd_0__inst_mult_6_86 ),
	.shareout(Xd_0__inst_mult_6_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_28 (
// Equation(s):
// Xd_0__inst_mult_7_90  = SUM(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_7_88  ) + ( Xd_0__inst_mult_7_87  ))
// Xd_0__inst_mult_7_91  = CARRY(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_7_88  ) + ( Xd_0__inst_mult_7_87  ))
// Xd_0__inst_mult_7_92  = SHARE((din_a[44] & din_b[45]))

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(!din_b[45]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_87 ),
	.sharein(Xd_0__inst_mult_7_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_90 ),
	.cout(Xd_0__inst_mult_7_91 ),
	.shareout(Xd_0__inst_mult_7_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_29 (
// Equation(s):
// Xd_0__inst_mult_7_94  = SUM(( (!din_a[46] & (((din_a[45] & din_b[43])))) # (din_a[46] & (!din_b[42] $ (((!din_a[45]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_7_112  ) + ( Xd_0__inst_mult_7_111  ))
// Xd_0__inst_mult_7_95  = CARRY(( (!din_a[46] & (((din_a[45] & din_b[43])))) # (din_a[46] & (!din_b[42] $ (((!din_a[45]) # (!din_b[43]))))) ) + ( Xd_0__inst_mult_7_112  ) + ( Xd_0__inst_mult_7_111  ))
// Xd_0__inst_mult_7_96  = SHARE((din_a[46] & (din_b[42] & (din_a[45] & din_b[43]))))

	.dataa(!din_a[46]),
	.datab(!din_b[42]),
	.datac(!din_a[45]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_111 ),
	.sharein(Xd_0__inst_mult_7_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_94 ),
	.cout(Xd_0__inst_mult_7_95 ),
	.shareout(Xd_0__inst_mult_7_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_26 (
// Equation(s):
// Xd_0__inst_mult_4_81  = SUM(( (din_a[26] & din_b[26]) ) + ( Xd_0__inst_mult_4_75  ) + ( Xd_0__inst_mult_4_74  ))
// Xd_0__inst_mult_4_82  = CARRY(( (din_a[26] & din_b[26]) ) + ( Xd_0__inst_mult_4_75  ) + ( Xd_0__inst_mult_4_74  ))
// Xd_0__inst_mult_4_83  = SHARE((din_a[26] & din_b[27]))

	.dataa(!din_a[26]),
	.datab(!din_b[26]),
	.datac(!din_b[27]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_74 ),
	.sharein(Xd_0__inst_mult_4_75 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_81 ),
	.cout(Xd_0__inst_mult_4_82 ),
	.shareout(Xd_0__inst_mult_4_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_27 (
// Equation(s):
// Xd_0__inst_mult_4_85  = SUM(( (!din_a[28] & (((din_a[27] & din_b[25])))) # (din_a[28] & (!din_b[24] $ (((!din_a[27]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_4_107  ) + ( Xd_0__inst_mult_4_106  ))
// Xd_0__inst_mult_4_86  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[25])))) # (din_a[28] & (!din_b[24] $ (((!din_a[27]) # (!din_b[25]))))) ) + ( Xd_0__inst_mult_4_107  ) + ( Xd_0__inst_mult_4_106  ))
// Xd_0__inst_mult_4_87  = SHARE((din_a[28] & (din_b[24] & (din_a[27] & din_b[25]))))

	.dataa(!din_a[28]),
	.datab(!din_b[24]),
	.datac(!din_a[27]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_106 ),
	.sharein(Xd_0__inst_mult_4_107 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_85 ),
	.cout(Xd_0__inst_mult_4_86 ),
	.shareout(Xd_0__inst_mult_4_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_27 (
// Equation(s):
// Xd_0__inst_mult_5_86  = SUM(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_5_84  ) + ( Xd_0__inst_mult_5_83  ))
// Xd_0__inst_mult_5_87  = CARRY(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_5_84  ) + ( Xd_0__inst_mult_5_83  ))
// Xd_0__inst_mult_5_88  = SHARE((din_a[32] & din_b[33]))

	.dataa(!din_a[32]),
	.datab(!din_b[32]),
	.datac(!din_b[33]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_83 ),
	.sharein(Xd_0__inst_mult_5_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_86 ),
	.cout(Xd_0__inst_mult_5_87 ),
	.shareout(Xd_0__inst_mult_5_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_28 (
// Equation(s):
// Xd_0__inst_mult_5_90  = SUM(( (!din_a[34] & (((din_a[33] & din_b[31])))) # (din_a[34] & (!din_b[30] $ (((!din_a[33]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_5_112  ) + ( Xd_0__inst_mult_5_111  ))
// Xd_0__inst_mult_5_91  = CARRY(( (!din_a[34] & (((din_a[33] & din_b[31])))) # (din_a[34] & (!din_b[30] $ (((!din_a[33]) # (!din_b[31]))))) ) + ( Xd_0__inst_mult_5_112  ) + ( Xd_0__inst_mult_5_111  ))
// Xd_0__inst_mult_5_92  = SHARE((din_a[34] & (din_b[30] & (din_a[33] & din_b[31]))))

	.dataa(!din_a[34]),
	.datab(!din_b[30]),
	.datac(!din_a[33]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_111 ),
	.sharein(Xd_0__inst_mult_5_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_90 ),
	.cout(Xd_0__inst_mult_5_91 ),
	.shareout(Xd_0__inst_mult_5_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_28 (
// Equation(s):
// Xd_0__inst_mult_2_90  = SUM(( (din_a[14] & din_b[14]) ) + ( Xd_0__inst_mult_2_88  ) + ( Xd_0__inst_mult_2_87  ))
// Xd_0__inst_mult_2_91  = CARRY(( (din_a[14] & din_b[14]) ) + ( Xd_0__inst_mult_2_88  ) + ( Xd_0__inst_mult_2_87  ))
// Xd_0__inst_mult_2_92  = SHARE((din_a[14] & din_b[15]))

	.dataa(!din_a[14]),
	.datab(!din_b[14]),
	.datac(!din_b[15]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_87 ),
	.sharein(Xd_0__inst_mult_2_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_90 ),
	.cout(Xd_0__inst_mult_2_91 ),
	.shareout(Xd_0__inst_mult_2_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_29 (
// Equation(s):
// Xd_0__inst_mult_2_94  = SUM(( (!din_a[16] & (((din_a[15] & din_b[13])))) # (din_a[16] & (!din_b[12] $ (((!din_a[15]) # (!din_b[13]))))) ) + ( Xd_0__inst_mult_2_112  ) + ( Xd_0__inst_mult_2_111  ))
// Xd_0__inst_mult_2_95  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[13])))) # (din_a[16] & (!din_b[12] $ (((!din_a[15]) # (!din_b[13]))))) ) + ( Xd_0__inst_mult_2_112  ) + ( Xd_0__inst_mult_2_111  ))
// Xd_0__inst_mult_2_96  = SHARE((din_a[16] & (din_b[12] & (din_a[15] & din_b[13]))))

	.dataa(!din_a[16]),
	.datab(!din_b[12]),
	.datac(!din_a[15]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_111 ),
	.sharein(Xd_0__inst_mult_2_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_94 ),
	.cout(Xd_0__inst_mult_2_95 ),
	.shareout(Xd_0__inst_mult_2_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_27 (
// Equation(s):
// Xd_0__inst_mult_3_86  = SUM(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_3_84  ) + ( Xd_0__inst_mult_3_83  ))
// Xd_0__inst_mult_3_87  = CARRY(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_3_84  ) + ( Xd_0__inst_mult_3_83  ))
// Xd_0__inst_mult_3_88  = SHARE((din_a[20] & din_b[21]))

	.dataa(!din_a[20]),
	.datab(!din_b[20]),
	.datac(!din_b[21]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_83 ),
	.sharein(Xd_0__inst_mult_3_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_86 ),
	.cout(Xd_0__inst_mult_3_87 ),
	.shareout(Xd_0__inst_mult_3_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_28 (
// Equation(s):
// Xd_0__inst_mult_3_90  = SUM(( (!din_a[22] & (((din_a[21] & din_b[19])))) # (din_a[22] & (!din_b[18] $ (((!din_a[21]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_3_112  ) + ( Xd_0__inst_mult_3_111  ))
// Xd_0__inst_mult_3_91  = CARRY(( (!din_a[22] & (((din_a[21] & din_b[19])))) # (din_a[22] & (!din_b[18] $ (((!din_a[21]) # (!din_b[19]))))) ) + ( Xd_0__inst_mult_3_112  ) + ( Xd_0__inst_mult_3_111  ))
// Xd_0__inst_mult_3_92  = SHARE((din_a[22] & (din_b[18] & (din_a[21] & din_b[19]))))

	.dataa(!din_a[22]),
	.datab(!din_b[18]),
	.datac(!din_a[21]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_111 ),
	.sharein(Xd_0__inst_mult_3_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_90 ),
	.cout(Xd_0__inst_mult_3_91 ),
	.shareout(Xd_0__inst_mult_3_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_28 (
// Equation(s):
// Xd_0__inst_mult_0_90  = SUM(( (din_a[2] & din_b[2]) ) + ( Xd_0__inst_mult_0_88  ) + ( Xd_0__inst_mult_0_87  ))
// Xd_0__inst_mult_0_91  = CARRY(( (din_a[2] & din_b[2]) ) + ( Xd_0__inst_mult_0_88  ) + ( Xd_0__inst_mult_0_87  ))
// Xd_0__inst_mult_0_92  = SHARE((din_a[2] & din_b[3]))

	.dataa(!din_a[2]),
	.datab(!din_b[2]),
	.datac(!din_b[3]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_87 ),
	.sharein(Xd_0__inst_mult_0_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_90 ),
	.cout(Xd_0__inst_mult_0_91 ),
	.shareout(Xd_0__inst_mult_0_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_29 (
// Equation(s):
// Xd_0__inst_mult_0_94  = SUM(( (!din_a[4] & (((din_a[3] & din_b[1])))) # (din_a[4] & (!din_b[0] $ (((!din_a[3]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_112  ) + ( Xd_0__inst_mult_0_111  ))
// Xd_0__inst_mult_0_95  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[1])))) # (din_a[4] & (!din_b[0] $ (((!din_a[3]) # (!din_b[1]))))) ) + ( Xd_0__inst_mult_0_112  ) + ( Xd_0__inst_mult_0_111  ))
// Xd_0__inst_mult_0_96  = SHARE((din_a[4] & (din_b[0] & (din_a[3] & din_b[1]))))

	.dataa(!din_a[4]),
	.datab(!din_b[0]),
	.datac(!din_a[3]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_111 ),
	.sharein(Xd_0__inst_mult_0_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_94 ),
	.cout(Xd_0__inst_mult_0_95 ),
	.shareout(Xd_0__inst_mult_0_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_27 (
// Equation(s):
// Xd_0__inst_mult_1_86  = SUM(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_1_84  ) + ( Xd_0__inst_mult_1_83  ))
// Xd_0__inst_mult_1_87  = CARRY(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_1_84  ) + ( Xd_0__inst_mult_1_83  ))
// Xd_0__inst_mult_1_88  = SHARE((din_a[8] & din_b[9]))

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(!din_b[9]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_83 ),
	.sharein(Xd_0__inst_mult_1_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_86 ),
	.cout(Xd_0__inst_mult_1_87 ),
	.shareout(Xd_0__inst_mult_1_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_28 (
// Equation(s):
// Xd_0__inst_mult_1_90  = SUM(( (!din_a[10] & (((din_a[9] & din_b[7])))) # (din_a[10] & (!din_b[6] $ (((!din_a[9]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_112  ) + ( Xd_0__inst_mult_1_111  ))
// Xd_0__inst_mult_1_91  = CARRY(( (!din_a[10] & (((din_a[9] & din_b[7])))) # (din_a[10] & (!din_b[6] $ (((!din_a[9]) # (!din_b[7]))))) ) + ( Xd_0__inst_mult_1_112  ) + ( Xd_0__inst_mult_1_111  ))
// Xd_0__inst_mult_1_92  = SHARE((din_a[10] & (din_b[6] & (din_a[9] & din_b[7]))))

	.dataa(!din_a[10]),
	.datab(!din_b[6]),
	.datac(!din_a[9]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_111 ),
	.sharein(Xd_0__inst_mult_1_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_90 ),
	.cout(Xd_0__inst_mult_1_91 ),
	.shareout(Xd_0__inst_mult_1_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_30 (
// Equation(s):
// Xd_0__inst_mult_28_99  = SUM(( (din_a[170] & din_b[170]) ) + ( Xd_0__inst_mult_28_97  ) + ( Xd_0__inst_mult_28_96  ))
// Xd_0__inst_mult_28_100  = CARRY(( (din_a[170] & din_b[170]) ) + ( Xd_0__inst_mult_28_97  ) + ( Xd_0__inst_mult_28_96  ))
// Xd_0__inst_mult_28_101  = SHARE((din_a[170] & din_b[171]))

	.dataa(!din_a[170]),
	.datab(!din_b[170]),
	.datac(!din_b[171]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_96 ),
	.sharein(Xd_0__inst_mult_28_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_99 ),
	.cout(Xd_0__inst_mult_28_100 ),
	.shareout(Xd_0__inst_mult_28_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_31 (
// Equation(s):
// Xd_0__inst_mult_29_103  = SUM(( (din_a[176] & din_b[176]) ) + ( Xd_0__inst_mult_29_101  ) + ( Xd_0__inst_mult_29_100  ))
// Xd_0__inst_mult_29_104  = CARRY(( (din_a[176] & din_b[176]) ) + ( Xd_0__inst_mult_29_101  ) + ( Xd_0__inst_mult_29_100  ))
// Xd_0__inst_mult_29_105  = SHARE((din_a[176] & din_b[177]))

	.dataa(!din_a[176]),
	.datab(!din_b[176]),
	.datac(!din_b[177]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_100 ),
	.sharein(Xd_0__inst_mult_29_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_103 ),
	.cout(Xd_0__inst_mult_29_104 ),
	.shareout(Xd_0__inst_mult_29_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_31 (
// Equation(s):
// Xd_0__inst_mult_26_103  = SUM(( (din_a[158] & din_b[158]) ) + ( Xd_0__inst_mult_26_101  ) + ( Xd_0__inst_mult_26_100  ))
// Xd_0__inst_mult_26_104  = CARRY(( (din_a[158] & din_b[158]) ) + ( Xd_0__inst_mult_26_101  ) + ( Xd_0__inst_mult_26_100  ))
// Xd_0__inst_mult_26_105  = SHARE((din_a[158] & din_b[159]))

	.dataa(!din_a[158]),
	.datab(!din_b[158]),
	.datac(!din_b[159]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_100 ),
	.sharein(Xd_0__inst_mult_26_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_103 ),
	.cout(Xd_0__inst_mult_26_104 ),
	.shareout(Xd_0__inst_mult_26_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_30 (
// Equation(s):
// Xd_0__inst_mult_27_99  = SUM(( (din_a[164] & din_b[164]) ) + ( Xd_0__inst_mult_27_97  ) + ( Xd_0__inst_mult_27_96  ))
// Xd_0__inst_mult_27_100  = CARRY(( (din_a[164] & din_b[164]) ) + ( Xd_0__inst_mult_27_97  ) + ( Xd_0__inst_mult_27_96  ))
// Xd_0__inst_mult_27_101  = SHARE((din_a[164] & din_b[165]))

	.dataa(!din_a[164]),
	.datab(!din_b[164]),
	.datac(!din_b[165]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_96 ),
	.sharein(Xd_0__inst_mult_27_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_99 ),
	.cout(Xd_0__inst_mult_27_100 ),
	.shareout(Xd_0__inst_mult_27_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_31 (
// Equation(s):
// Xd_0__inst_mult_24_103  = SUM(( (din_a[146] & din_b[146]) ) + ( Xd_0__inst_mult_24_101  ) + ( Xd_0__inst_mult_24_100  ))
// Xd_0__inst_mult_24_104  = CARRY(( (din_a[146] & din_b[146]) ) + ( Xd_0__inst_mult_24_101  ) + ( Xd_0__inst_mult_24_100  ))
// Xd_0__inst_mult_24_105  = SHARE((din_a[146] & din_b[147]))

	.dataa(!din_a[146]),
	.datab(!din_b[146]),
	.datac(!din_b[147]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_100 ),
	.sharein(Xd_0__inst_mult_24_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_103 ),
	.cout(Xd_0__inst_mult_24_104 ),
	.shareout(Xd_0__inst_mult_24_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_30 (
// Equation(s):
// Xd_0__inst_mult_25_99  = SUM(( (din_a[152] & din_b[152]) ) + ( Xd_0__inst_mult_25_97  ) + ( Xd_0__inst_mult_25_96  ))
// Xd_0__inst_mult_25_100  = CARRY(( (din_a[152] & din_b[152]) ) + ( Xd_0__inst_mult_25_97  ) + ( Xd_0__inst_mult_25_96  ))
// Xd_0__inst_mult_25_101  = SHARE((din_a[152] & din_b[153]))

	.dataa(!din_a[152]),
	.datab(!din_b[152]),
	.datac(!din_b[153]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_96 ),
	.sharein(Xd_0__inst_mult_25_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_99 ),
	.cout(Xd_0__inst_mult_25_100 ),
	.shareout(Xd_0__inst_mult_25_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_31 (
// Equation(s):
// Xd_0__inst_mult_22_103  = SUM(( (din_a[134] & din_b[134]) ) + ( Xd_0__inst_mult_22_101  ) + ( Xd_0__inst_mult_22_100  ))
// Xd_0__inst_mult_22_104  = CARRY(( (din_a[134] & din_b[134]) ) + ( Xd_0__inst_mult_22_101  ) + ( Xd_0__inst_mult_22_100  ))
// Xd_0__inst_mult_22_105  = SHARE((din_a[134] & din_b[135]))

	.dataa(!din_a[134]),
	.datab(!din_b[134]),
	.datac(!din_b[135]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_100 ),
	.sharein(Xd_0__inst_mult_22_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_103 ),
	.cout(Xd_0__inst_mult_22_104 ),
	.shareout(Xd_0__inst_mult_22_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_30 (
// Equation(s):
// Xd_0__inst_mult_23_99  = SUM(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_23_97  ) + ( Xd_0__inst_mult_23_96  ))
// Xd_0__inst_mult_23_100  = CARRY(( (din_a[140] & din_b[140]) ) + ( Xd_0__inst_mult_23_97  ) + ( Xd_0__inst_mult_23_96  ))
// Xd_0__inst_mult_23_101  = SHARE((din_a[140] & din_b[141]))

	.dataa(!din_a[140]),
	.datab(!din_b[140]),
	.datac(!din_b[141]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_96 ),
	.sharein(Xd_0__inst_mult_23_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_99 ),
	.cout(Xd_0__inst_mult_23_100 ),
	.shareout(Xd_0__inst_mult_23_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_30 (
// Equation(s):
// Xd_0__inst_mult_20_99  = SUM(( (din_a[122] & din_b[122]) ) + ( Xd_0__inst_mult_20_97  ) + ( Xd_0__inst_mult_20_96  ))
// Xd_0__inst_mult_20_100  = CARRY(( (din_a[122] & din_b[122]) ) + ( Xd_0__inst_mult_20_97  ) + ( Xd_0__inst_mult_20_96  ))
// Xd_0__inst_mult_20_101  = SHARE((din_a[122] & din_b[123]))

	.dataa(!din_a[122]),
	.datab(!din_b[122]),
	.datac(!din_b[123]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_96 ),
	.sharein(Xd_0__inst_mult_20_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_99 ),
	.cout(Xd_0__inst_mult_20_100 ),
	.shareout(Xd_0__inst_mult_20_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_28 (
// Equation(s):
// Xd_0__inst_mult_21_91  = SUM(( (din_a[128] & din_b[128]) ) + ( Xd_0__inst_mult_21_89  ) + ( Xd_0__inst_mult_21_88  ))
// Xd_0__inst_mult_21_92  = CARRY(( (din_a[128] & din_b[128]) ) + ( Xd_0__inst_mult_21_89  ) + ( Xd_0__inst_mult_21_88  ))
// Xd_0__inst_mult_21_93  = SHARE((din_a[128] & din_b[129]))

	.dataa(!din_a[128]),
	.datab(!din_b[128]),
	.datac(!din_b[129]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_88 ),
	.sharein(Xd_0__inst_mult_21_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_91 ),
	.cout(Xd_0__inst_mult_21_92 ),
	.shareout(Xd_0__inst_mult_21_93 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_29 (
// Equation(s):
// Xd_0__inst_mult_21_95  = SUM(( (!din_a[130] & (((din_a[129] & din_b[127])))) # (din_a[130] & (!din_b[126] $ (((!din_a[129]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_21_117  ) + ( Xd_0__inst_mult_21_116  ))
// Xd_0__inst_mult_21_96  = CARRY(( (!din_a[130] & (((din_a[129] & din_b[127])))) # (din_a[130] & (!din_b[126] $ (((!din_a[129]) # (!din_b[127]))))) ) + ( Xd_0__inst_mult_21_117  ) + ( Xd_0__inst_mult_21_116  ))
// Xd_0__inst_mult_21_97  = SHARE((din_a[130] & (din_b[126] & (din_a[129] & din_b[127]))))

	.dataa(!din_a[130]),
	.datab(!din_b[126]),
	.datac(!din_a[129]),
	.datad(!din_b[127]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_116 ),
	.sharein(Xd_0__inst_mult_21_117 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_95 ),
	.cout(Xd_0__inst_mult_21_96 ),
	.shareout(Xd_0__inst_mult_21_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_26 (
// Equation(s):
// Xd_0__inst_mult_18_82  = SUM(( (din_a[110] & din_b[110]) ) + ( Xd_0__inst_mult_18_76  ) + ( Xd_0__inst_mult_18_75  ))
// Xd_0__inst_mult_18_83  = CARRY(( (din_a[110] & din_b[110]) ) + ( Xd_0__inst_mult_18_76  ) + ( Xd_0__inst_mult_18_75  ))
// Xd_0__inst_mult_18_84  = SHARE((din_a[110] & din_b[111]))

	.dataa(!din_a[110]),
	.datab(!din_b[110]),
	.datac(!din_b[111]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_75 ),
	.sharein(Xd_0__inst_mult_18_76 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_82 ),
	.cout(Xd_0__inst_mult_18_83 ),
	.shareout(Xd_0__inst_mult_18_84 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_27 (
// Equation(s):
// Xd_0__inst_mult_18_86  = SUM(( (!din_a[112] & (((din_a[111] & din_b[109])))) # (din_a[112] & (!din_b[108] $ (((!din_a[111]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_18_112  ) + ( Xd_0__inst_mult_18_111  ))
// Xd_0__inst_mult_18_87  = CARRY(( (!din_a[112] & (((din_a[111] & din_b[109])))) # (din_a[112] & (!din_b[108] $ (((!din_a[111]) # (!din_b[109]))))) ) + ( Xd_0__inst_mult_18_112  ) + ( Xd_0__inst_mult_18_111  ))
// Xd_0__inst_mult_18_88  = SHARE((din_a[112] & (din_b[108] & (din_a[111] & din_b[109]))))

	.dataa(!din_a[112]),
	.datab(!din_b[108]),
	.datac(!din_a[111]),
	.datad(!din_b[109]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_111 ),
	.sharein(Xd_0__inst_mult_18_112 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_86 ),
	.cout(Xd_0__inst_mult_18_87 ),
	.shareout(Xd_0__inst_mult_18_88 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_31 (
// Equation(s):
// Xd_0__inst_mult_19_103  = SUM(( (din_a[116] & din_b[116]) ) + ( Xd_0__inst_mult_19_101  ) + ( Xd_0__inst_mult_19_100  ))
// Xd_0__inst_mult_19_104  = CARRY(( (din_a[116] & din_b[116]) ) + ( Xd_0__inst_mult_19_101  ) + ( Xd_0__inst_mult_19_100  ))
// Xd_0__inst_mult_19_105  = SHARE((din_a[116] & din_b[117]))

	.dataa(!din_a[116]),
	.datab(!din_b[116]),
	.datac(!din_b[117]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_100 ),
	.sharein(Xd_0__inst_mult_19_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_103 ),
	.cout(Xd_0__inst_mult_19_104 ),
	.shareout(Xd_0__inst_mult_19_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_28 (
// Equation(s):
// Xd_0__inst_mult_16_90  = SUM(( (!din_a[100] & (((din_a[99] & din_b[98])))) # (din_a[100] & (!din_b[97] $ (((!din_a[99]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_16_84  ) + ( Xd_0__inst_mult_16_83  ))
// Xd_0__inst_mult_16_91  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[98])))) # (din_a[100] & (!din_b[97] $ (((!din_a[99]) # (!din_b[98]))))) ) + ( Xd_0__inst_mult_16_84  ) + ( Xd_0__inst_mult_16_83  ))
// Xd_0__inst_mult_16_92  = SHARE((din_a[100] & (din_b[97] & (din_a[99] & din_b[98]))))

	.dataa(!din_a[100]),
	.datab(!din_b[97]),
	.datac(!din_a[99]),
	.datad(!din_b[98]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_83 ),
	.sharein(Xd_0__inst_mult_16_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_90 ),
	.cout(Xd_0__inst_mult_16_91 ),
	.shareout(Xd_0__inst_mult_16_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_29 (
// Equation(s):
// Xd_0__inst_mult_16_94  = SUM(( GND ) + ( Xd_0__inst_mult_16_88  ) + ( Xd_0__inst_mult_16_87  ))
// Xd_0__inst_mult_16_95  = CARRY(( GND ) + ( Xd_0__inst_mult_16_88  ) + ( Xd_0__inst_mult_16_87  ))
// Xd_0__inst_mult_16_96  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_87 ),
	.sharein(Xd_0__inst_mult_16_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_94 ),
	.cout(Xd_0__inst_mult_16_95 ),
	.shareout(Xd_0__inst_mult_16_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_30 (
// Equation(s):
// Xd_0__inst_mult_17_99  = SUM(( (!din_a[106] & (((din_a[105] & din_b[104])))) # (din_a[106] & (!din_b[103] $ (((!din_a[105]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_17_93  ) + ( Xd_0__inst_mult_17_92  ))
// Xd_0__inst_mult_17_100  = CARRY(( (!din_a[106] & (((din_a[105] & din_b[104])))) # (din_a[106] & (!din_b[103] $ (((!din_a[105]) # (!din_b[104]))))) ) + ( Xd_0__inst_mult_17_93  ) + ( Xd_0__inst_mult_17_92  ))
// Xd_0__inst_mult_17_101  = SHARE((din_a[106] & (din_b[103] & (din_a[105] & din_b[104]))))

	.dataa(!din_a[106]),
	.datab(!din_b[103]),
	.datac(!din_a[105]),
	.datad(!din_b[104]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_92 ),
	.sharein(Xd_0__inst_mult_17_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_99 ),
	.cout(Xd_0__inst_mult_17_100 ),
	.shareout(Xd_0__inst_mult_17_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_31 (
// Equation(s):
// Xd_0__inst_mult_17_103  = SUM(( GND ) + ( Xd_0__inst_mult_17_97  ) + ( Xd_0__inst_mult_17_96  ))
// Xd_0__inst_mult_17_104  = CARRY(( GND ) + ( Xd_0__inst_mult_17_97  ) + ( Xd_0__inst_mult_17_96  ))
// Xd_0__inst_mult_17_105  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_96 ),
	.sharein(Xd_0__inst_mult_17_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_103 ),
	.cout(Xd_0__inst_mult_17_104 ),
	.shareout(Xd_0__inst_mult_17_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_28 (
// Equation(s):
// Xd_0__inst_mult_14_90  = SUM(( (!din_a[88] & (((din_a[87] & din_b[86])))) # (din_a[88] & (!din_b[85] $ (((!din_a[87]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_14_84  ) + ( Xd_0__inst_mult_14_83  ))
// Xd_0__inst_mult_14_91  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[86])))) # (din_a[88] & (!din_b[85] $ (((!din_a[87]) # (!din_b[86]))))) ) + ( Xd_0__inst_mult_14_84  ) + ( Xd_0__inst_mult_14_83  ))
// Xd_0__inst_mult_14_92  = SHARE((din_a[88] & (din_b[85] & (din_a[87] & din_b[86]))))

	.dataa(!din_a[88]),
	.datab(!din_b[85]),
	.datac(!din_a[87]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_83 ),
	.sharein(Xd_0__inst_mult_14_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_90 ),
	.cout(Xd_0__inst_mult_14_91 ),
	.shareout(Xd_0__inst_mult_14_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_29 (
// Equation(s):
// Xd_0__inst_mult_14_94  = SUM(( GND ) + ( Xd_0__inst_mult_14_88  ) + ( Xd_0__inst_mult_14_87  ))
// Xd_0__inst_mult_14_95  = CARRY(( GND ) + ( Xd_0__inst_mult_14_88  ) + ( Xd_0__inst_mult_14_87  ))
// Xd_0__inst_mult_14_96  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_87 ),
	.sharein(Xd_0__inst_mult_14_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_94 ),
	.cout(Xd_0__inst_mult_14_95 ),
	.shareout(Xd_0__inst_mult_14_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_30 (
// Equation(s):
// Xd_0__inst_mult_15_99  = SUM(( (!din_a[94] & (((din_a[93] & din_b[92])))) # (din_a[94] & (!din_b[91] $ (((!din_a[93]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_15_93  ) + ( Xd_0__inst_mult_15_92  ))
// Xd_0__inst_mult_15_100  = CARRY(( (!din_a[94] & (((din_a[93] & din_b[92])))) # (din_a[94] & (!din_b[91] $ (((!din_a[93]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_15_93  ) + ( Xd_0__inst_mult_15_92  ))
// Xd_0__inst_mult_15_101  = SHARE((din_a[94] & (din_b[91] & (din_a[93] & din_b[92]))))

	.dataa(!din_a[94]),
	.datab(!din_b[91]),
	.datac(!din_a[93]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_92 ),
	.sharein(Xd_0__inst_mult_15_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_99 ),
	.cout(Xd_0__inst_mult_15_100 ),
	.shareout(Xd_0__inst_mult_15_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_31 (
// Equation(s):
// Xd_0__inst_mult_15_103  = SUM(( GND ) + ( Xd_0__inst_mult_15_97  ) + ( Xd_0__inst_mult_15_96  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_96 ),
	.sharein(Xd_0__inst_mult_15_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_103 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_29 (
// Equation(s):
// Xd_0__inst_mult_12_94  = SUM(( (!din_a[76] & (((din_a[75] & din_b[74])))) # (din_a[76] & (!din_b[73] $ (((!din_a[75]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_12_88  ) + ( Xd_0__inst_mult_12_87  ))
// Xd_0__inst_mult_12_95  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[74])))) # (din_a[76] & (!din_b[73] $ (((!din_a[75]) # (!din_b[74]))))) ) + ( Xd_0__inst_mult_12_88  ) + ( Xd_0__inst_mult_12_87  ))
// Xd_0__inst_mult_12_96  = SHARE((din_a[76] & (din_b[73] & (din_a[75] & din_b[74]))))

	.dataa(!din_a[76]),
	.datab(!din_b[73]),
	.datac(!din_a[75]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_87 ),
	.sharein(Xd_0__inst_mult_12_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_94 ),
	.cout(Xd_0__inst_mult_12_95 ),
	.shareout(Xd_0__inst_mult_12_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_30 (
// Equation(s):
// Xd_0__inst_mult_12_98  = SUM(( GND ) + ( Xd_0__inst_mult_12_92  ) + ( Xd_0__inst_mult_12_91  ))
// Xd_0__inst_mult_12_99  = CARRY(( GND ) + ( Xd_0__inst_mult_12_92  ) + ( Xd_0__inst_mult_12_91  ))
// Xd_0__inst_mult_12_100  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_91 ),
	.sharein(Xd_0__inst_mult_12_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_98 ),
	.cout(Xd_0__inst_mult_12_99 ),
	.shareout(Xd_0__inst_mult_12_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_29 (
// Equation(s):
// Xd_0__inst_mult_13_95  = SUM(( (!din_a[82] & (((din_a[81] & din_b[80])))) # (din_a[82] & (!din_b[79] $ (((!din_a[81]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_13_89  ) + ( Xd_0__inst_mult_13_88  ))
// Xd_0__inst_mult_13_96  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[80])))) # (din_a[82] & (!din_b[79] $ (((!din_a[81]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_13_89  ) + ( Xd_0__inst_mult_13_88  ))
// Xd_0__inst_mult_13_97  = SHARE((din_a[82] & (din_b[79] & (din_a[81] & din_b[80]))))

	.dataa(!din_a[82]),
	.datab(!din_b[79]),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_88 ),
	.sharein(Xd_0__inst_mult_13_89 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_95 ),
	.cout(Xd_0__inst_mult_13_96 ),
	.shareout(Xd_0__inst_mult_13_97 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_30 (
// Equation(s):
// Xd_0__inst_mult_13_99  = SUM(( GND ) + ( Xd_0__inst_mult_13_93  ) + ( Xd_0__inst_mult_13_92  ))
// Xd_0__inst_mult_13_100  = CARRY(( GND ) + ( Xd_0__inst_mult_13_93  ) + ( Xd_0__inst_mult_13_92  ))
// Xd_0__inst_mult_13_101  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_92 ),
	.sharein(Xd_0__inst_mult_13_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_99 ),
	.cout(Xd_0__inst_mult_13_100 ),
	.shareout(Xd_0__inst_mult_13_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_28 (
// Equation(s):
// Xd_0__inst_mult_10_90  = SUM(( (!din_a[64] & (((din_a[63] & din_b[62])))) # (din_a[64] & (!din_b[61] $ (((!din_a[63]) # (!din_b[62]))))) ) + ( Xd_0__inst_mult_10_84  ) + ( Xd_0__inst_mult_10_83  ))
// Xd_0__inst_mult_10_91  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[62])))) # (din_a[64] & (!din_b[61] $ (((!din_a[63]) # (!din_b[62]))))) ) + ( Xd_0__inst_mult_10_84  ) + ( Xd_0__inst_mult_10_83  ))
// Xd_0__inst_mult_10_92  = SHARE((din_a[64] & (din_b[61] & (din_a[63] & din_b[62]))))

	.dataa(!din_a[64]),
	.datab(!din_b[61]),
	.datac(!din_a[63]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_83 ),
	.sharein(Xd_0__inst_mult_10_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_90 ),
	.cout(Xd_0__inst_mult_10_91 ),
	.shareout(Xd_0__inst_mult_10_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_29 (
// Equation(s):
// Xd_0__inst_mult_10_94  = SUM(( GND ) + ( Xd_0__inst_mult_10_88  ) + ( Xd_0__inst_mult_10_87  ))
// Xd_0__inst_mult_10_95  = CARRY(( GND ) + ( Xd_0__inst_mult_10_88  ) + ( Xd_0__inst_mult_10_87  ))
// Xd_0__inst_mult_10_96  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_87 ),
	.sharein(Xd_0__inst_mult_10_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_94 ),
	.cout(Xd_0__inst_mult_10_95 ),
	.shareout(Xd_0__inst_mult_10_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_32 (
// Equation(s):
// Xd_0__inst_mult_11_107  = SUM(( (!din_a[70] & (((din_a[69] & din_b[68])))) # (din_a[70] & (!din_b[67] $ (((!din_a[69]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_11_105  ) + ( Xd_0__inst_mult_11_104  ))
// Xd_0__inst_mult_11_108  = CARRY(( (!din_a[70] & (((din_a[69] & din_b[68])))) # (din_a[70] & (!din_b[67] $ (((!din_a[69]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_11_105  ) + ( Xd_0__inst_mult_11_104  ))
// Xd_0__inst_mult_11_109  = SHARE((din_a[70] & (din_b[67] & (din_a[69] & din_b[68]))))

	.dataa(!din_a[70]),
	.datab(!din_b[67]),
	.datac(!din_a[69]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_104 ),
	.sharein(Xd_0__inst_mult_11_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_107 ),
	.cout(Xd_0__inst_mult_11_108 ),
	.shareout(Xd_0__inst_mult_11_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_29 (
// Equation(s):
// Xd_0__inst_mult_8_94  = SUM(( (!din_a[52] & (((din_a[51] & din_b[50])))) # (din_a[52] & (!din_b[49] $ (((!din_a[51]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_8_88  ) + ( Xd_0__inst_mult_8_87  ))
// Xd_0__inst_mult_8_95  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[50])))) # (din_a[52] & (!din_b[49] $ (((!din_a[51]) # (!din_b[50]))))) ) + ( Xd_0__inst_mult_8_88  ) + ( Xd_0__inst_mult_8_87  ))
// Xd_0__inst_mult_8_96  = SHARE((din_a[52] & (din_b[49] & (din_a[51] & din_b[50]))))

	.dataa(!din_a[52]),
	.datab(!din_b[49]),
	.datac(!din_a[51]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_87 ),
	.sharein(Xd_0__inst_mult_8_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_94 ),
	.cout(Xd_0__inst_mult_8_95 ),
	.shareout(Xd_0__inst_mult_8_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_30 (
// Equation(s):
// Xd_0__inst_mult_8_98  = SUM(( GND ) + ( Xd_0__inst_mult_8_92  ) + ( Xd_0__inst_mult_8_91  ))
// Xd_0__inst_mult_8_99  = CARRY(( GND ) + ( Xd_0__inst_mult_8_92  ) + ( Xd_0__inst_mult_8_91  ))
// Xd_0__inst_mult_8_100  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_91 ),
	.sharein(Xd_0__inst_mult_8_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_98 ),
	.cout(Xd_0__inst_mult_8_99 ),
	.shareout(Xd_0__inst_mult_8_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_30 (
// Equation(s):
// Xd_0__inst_mult_9_99  = SUM(( (!din_a[58] & (((din_a[57] & din_b[56])))) # (din_a[58] & (!din_b[55] $ (((!din_a[57]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_9_93  ) + ( Xd_0__inst_mult_9_92  ))
// Xd_0__inst_mult_9_100  = CARRY(( (!din_a[58] & (((din_a[57] & din_b[56])))) # (din_a[58] & (!din_b[55] $ (((!din_a[57]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_9_93  ) + ( Xd_0__inst_mult_9_92  ))
// Xd_0__inst_mult_9_101  = SHARE((din_a[58] & (din_b[55] & (din_a[57] & din_b[56]))))

	.dataa(!din_a[58]),
	.datab(!din_b[55]),
	.datac(!din_a[57]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_92 ),
	.sharein(Xd_0__inst_mult_9_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_99 ),
	.cout(Xd_0__inst_mult_9_100 ),
	.shareout(Xd_0__inst_mult_9_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_31 (
// Equation(s):
// Xd_0__inst_mult_9_103  = SUM(( GND ) + ( Xd_0__inst_mult_9_97  ) + ( Xd_0__inst_mult_9_96  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_96 ),
	.sharein(Xd_0__inst_mult_9_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_103 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_28 (
// Equation(s):
// Xd_0__inst_mult_6_89  = SUM(( (!din_a[40] & (((din_a[39] & din_b[38])))) # (din_a[40] & (!din_b[37] $ (((!din_a[39]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_6_83  ) + ( Xd_0__inst_mult_6_82  ))
// Xd_0__inst_mult_6_90  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[38])))) # (din_a[40] & (!din_b[37] $ (((!din_a[39]) # (!din_b[38]))))) ) + ( Xd_0__inst_mult_6_83  ) + ( Xd_0__inst_mult_6_82  ))
// Xd_0__inst_mult_6_91  = SHARE((din_a[40] & (din_b[37] & (din_a[39] & din_b[38]))))

	.dataa(!din_a[40]),
	.datab(!din_b[37]),
	.datac(!din_a[39]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_82 ),
	.sharein(Xd_0__inst_mult_6_83 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_89 ),
	.cout(Xd_0__inst_mult_6_90 ),
	.shareout(Xd_0__inst_mult_6_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_30 (
// Equation(s):
// Xd_0__inst_mult_7_98  = SUM(( (!din_a[46] & (((din_a[45] & din_b[44])))) # (din_a[46] & (!din_b[43] $ (((!din_a[45]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_7_92  ) + ( Xd_0__inst_mult_7_91  ))
// Xd_0__inst_mult_7_99  = CARRY(( (!din_a[46] & (((din_a[45] & din_b[44])))) # (din_a[46] & (!din_b[43] $ (((!din_a[45]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_7_92  ) + ( Xd_0__inst_mult_7_91  ))
// Xd_0__inst_mult_7_100  = SHARE((din_a[46] & (din_b[43] & (din_a[45] & din_b[44]))))

	.dataa(!din_a[46]),
	.datab(!din_b[43]),
	.datac(!din_a[45]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_91 ),
	.sharein(Xd_0__inst_mult_7_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_98 ),
	.cout(Xd_0__inst_mult_7_99 ),
	.shareout(Xd_0__inst_mult_7_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_28 (
// Equation(s):
// Xd_0__inst_mult_4_89  = SUM(( (!din_a[28] & (((din_a[27] & din_b[26])))) # (din_a[28] & (!din_b[25] $ (((!din_a[27]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_4_83  ) + ( Xd_0__inst_mult_4_82  ))
// Xd_0__inst_mult_4_90  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[26])))) # (din_a[28] & (!din_b[25] $ (((!din_a[27]) # (!din_b[26]))))) ) + ( Xd_0__inst_mult_4_83  ) + ( Xd_0__inst_mult_4_82  ))
// Xd_0__inst_mult_4_91  = SHARE((din_a[28] & (din_b[25] & (din_a[27] & din_b[26]))))

	.dataa(!din_a[28]),
	.datab(!din_b[25]),
	.datac(!din_a[27]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_82 ),
	.sharein(Xd_0__inst_mult_4_83 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_89 ),
	.cout(Xd_0__inst_mult_4_90 ),
	.shareout(Xd_0__inst_mult_4_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_29 (
// Equation(s):
// Xd_0__inst_mult_5_94  = SUM(( (!din_a[34] & (((din_a[33] & din_b[32])))) # (din_a[34] & (!din_b[31] $ (((!din_a[33]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_5_88  ) + ( Xd_0__inst_mult_5_87  ))
// Xd_0__inst_mult_5_95  = CARRY(( (!din_a[34] & (((din_a[33] & din_b[32])))) # (din_a[34] & (!din_b[31] $ (((!din_a[33]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_5_88  ) + ( Xd_0__inst_mult_5_87  ))
// Xd_0__inst_mult_5_96  = SHARE((din_a[34] & (din_b[31] & (din_a[33] & din_b[32]))))

	.dataa(!din_a[34]),
	.datab(!din_b[31]),
	.datac(!din_a[33]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_87 ),
	.sharein(Xd_0__inst_mult_5_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_94 ),
	.cout(Xd_0__inst_mult_5_95 ),
	.shareout(Xd_0__inst_mult_5_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_30 (
// Equation(s):
// Xd_0__inst_mult_2_98  = SUM(( (!din_a[16] & (((din_a[15] & din_b[14])))) # (din_a[16] & (!din_b[13] $ (((!din_a[15]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_92  ) + ( Xd_0__inst_mult_2_91  ))
// Xd_0__inst_mult_2_99  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[14])))) # (din_a[16] & (!din_b[13] $ (((!din_a[15]) # (!din_b[14]))))) ) + ( Xd_0__inst_mult_2_92  ) + ( Xd_0__inst_mult_2_91  ))
// Xd_0__inst_mult_2_100  = SHARE((din_a[16] & (din_b[13] & (din_a[15] & din_b[14]))))

	.dataa(!din_a[16]),
	.datab(!din_b[13]),
	.datac(!din_a[15]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_91 ),
	.sharein(Xd_0__inst_mult_2_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_98 ),
	.cout(Xd_0__inst_mult_2_99 ),
	.shareout(Xd_0__inst_mult_2_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_29 (
// Equation(s):
// Xd_0__inst_mult_3_94  = SUM(( (!din_a[22] & (((din_a[21] & din_b[20])))) # (din_a[22] & (!din_b[19] $ (((!din_a[21]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_3_88  ) + ( Xd_0__inst_mult_3_87  ))
// Xd_0__inst_mult_3_95  = CARRY(( (!din_a[22] & (((din_a[21] & din_b[20])))) # (din_a[22] & (!din_b[19] $ (((!din_a[21]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_3_88  ) + ( Xd_0__inst_mult_3_87  ))
// Xd_0__inst_mult_3_96  = SHARE((din_a[22] & (din_b[19] & (din_a[21] & din_b[20]))))

	.dataa(!din_a[22]),
	.datab(!din_b[19]),
	.datac(!din_a[21]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_87 ),
	.sharein(Xd_0__inst_mult_3_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_94 ),
	.cout(Xd_0__inst_mult_3_95 ),
	.shareout(Xd_0__inst_mult_3_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_30 (
// Equation(s):
// Xd_0__inst_mult_0_98  = SUM(( (!din_a[4] & (((din_a[3] & din_b[2])))) # (din_a[4] & (!din_b[1] $ (((!din_a[3]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_92  ) + ( Xd_0__inst_mult_0_91  ))
// Xd_0__inst_mult_0_99  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[2])))) # (din_a[4] & (!din_b[1] $ (((!din_a[3]) # (!din_b[2]))))) ) + ( Xd_0__inst_mult_0_92  ) + ( Xd_0__inst_mult_0_91  ))
// Xd_0__inst_mult_0_100  = SHARE((din_a[4] & (din_b[1] & (din_a[3] & din_b[2]))))

	.dataa(!din_a[4]),
	.datab(!din_b[1]),
	.datac(!din_a[3]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_91 ),
	.sharein(Xd_0__inst_mult_0_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_98 ),
	.cout(Xd_0__inst_mult_0_99 ),
	.shareout(Xd_0__inst_mult_0_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_29 (
// Equation(s):
// Xd_0__inst_mult_1_94  = SUM(( (!din_a[10] & (((din_a[9] & din_b[8])))) # (din_a[10] & (!din_b[7] $ (((!din_a[9]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_88  ) + ( Xd_0__inst_mult_1_87  ))
// Xd_0__inst_mult_1_95  = CARRY(( (!din_a[10] & (((din_a[9] & din_b[8])))) # (din_a[10] & (!din_b[7] $ (((!din_a[9]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_1_88  ) + ( Xd_0__inst_mult_1_87  ))
// Xd_0__inst_mult_1_96  = SHARE((din_a[10] & (din_b[7] & (din_a[9] & din_b[8]))))

	.dataa(!din_a[10]),
	.datab(!din_b[7]),
	.datac(!din_a[9]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_87 ),
	.sharein(Xd_0__inst_mult_1_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_94 ),
	.cout(Xd_0__inst_mult_1_95 ),
	.shareout(Xd_0__inst_mult_1_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_31 (
// Equation(s):
// Xd_0__inst_mult_28_103  = SUM(( (!din_a[172] & (((din_a[171] & din_b[170])))) # (din_a[172] & (!din_b[169] $ (((!din_a[171]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_28_101  ) + ( Xd_0__inst_mult_28_100  ))
// Xd_0__inst_mult_28_104  = CARRY(( (!din_a[172] & (((din_a[171] & din_b[170])))) # (din_a[172] & (!din_b[169] $ (((!din_a[171]) # (!din_b[170]))))) ) + ( Xd_0__inst_mult_28_101  ) + ( Xd_0__inst_mult_28_100  ))
// Xd_0__inst_mult_28_105  = SHARE((din_a[172] & (din_b[169] & (din_a[171] & din_b[170]))))

	.dataa(!din_a[172]),
	.datab(!din_b[169]),
	.datac(!din_a[171]),
	.datad(!din_b[170]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_100 ),
	.sharein(Xd_0__inst_mult_28_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_103 ),
	.cout(Xd_0__inst_mult_28_104 ),
	.shareout(Xd_0__inst_mult_28_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_32 (
// Equation(s):
// Xd_0__inst_mult_29_107  = SUM(( (!din_a[178] & (((din_a[177] & din_b[176])))) # (din_a[178] & (!din_b[175] $ (((!din_a[177]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_29_105  ) + ( Xd_0__inst_mult_29_104  ))
// Xd_0__inst_mult_29_108  = CARRY(( (!din_a[178] & (((din_a[177] & din_b[176])))) # (din_a[178] & (!din_b[175] $ (((!din_a[177]) # (!din_b[176]))))) ) + ( Xd_0__inst_mult_29_105  ) + ( Xd_0__inst_mult_29_104  ))
// Xd_0__inst_mult_29_109  = SHARE((din_a[178] & (din_b[175] & (din_a[177] & din_b[176]))))

	.dataa(!din_a[178]),
	.datab(!din_b[175]),
	.datac(!din_a[177]),
	.datad(!din_b[176]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_104 ),
	.sharein(Xd_0__inst_mult_29_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_107 ),
	.cout(Xd_0__inst_mult_29_108 ),
	.shareout(Xd_0__inst_mult_29_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_32 (
// Equation(s):
// Xd_0__inst_mult_26_107  = SUM(( (!din_a[160] & (((din_a[159] & din_b[158])))) # (din_a[160] & (!din_b[157] $ (((!din_a[159]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_26_105  ) + ( Xd_0__inst_mult_26_104  ))
// Xd_0__inst_mult_26_108  = CARRY(( (!din_a[160] & (((din_a[159] & din_b[158])))) # (din_a[160] & (!din_b[157] $ (((!din_a[159]) # (!din_b[158]))))) ) + ( Xd_0__inst_mult_26_105  ) + ( Xd_0__inst_mult_26_104  ))
// Xd_0__inst_mult_26_109  = SHARE((din_a[160] & (din_b[157] & (din_a[159] & din_b[158]))))

	.dataa(!din_a[160]),
	.datab(!din_b[157]),
	.datac(!din_a[159]),
	.datad(!din_b[158]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_104 ),
	.sharein(Xd_0__inst_mult_26_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_107 ),
	.cout(Xd_0__inst_mult_26_108 ),
	.shareout(Xd_0__inst_mult_26_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_31 (
// Equation(s):
// Xd_0__inst_mult_27_103  = SUM(( (!din_a[166] & (((din_a[165] & din_b[164])))) # (din_a[166] & (!din_b[163] $ (((!din_a[165]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_27_101  ) + ( Xd_0__inst_mult_27_100  ))
// Xd_0__inst_mult_27_104  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[164])))) # (din_a[166] & (!din_b[163] $ (((!din_a[165]) # (!din_b[164]))))) ) + ( Xd_0__inst_mult_27_101  ) + ( Xd_0__inst_mult_27_100  ))
// Xd_0__inst_mult_27_105  = SHARE((din_a[166] & (din_b[163] & (din_a[165] & din_b[164]))))

	.dataa(!din_a[166]),
	.datab(!din_b[163]),
	.datac(!din_a[165]),
	.datad(!din_b[164]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_100 ),
	.sharein(Xd_0__inst_mult_27_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_103 ),
	.cout(Xd_0__inst_mult_27_104 ),
	.shareout(Xd_0__inst_mult_27_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_32 (
// Equation(s):
// Xd_0__inst_mult_24_107  = SUM(( (!din_a[148] & (((din_a[147] & din_b[146])))) # (din_a[148] & (!din_b[145] $ (((!din_a[147]) # (!din_b[146]))))) ) + ( Xd_0__inst_mult_24_105  ) + ( Xd_0__inst_mult_24_104  ))
// Xd_0__inst_mult_24_108  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[146])))) # (din_a[148] & (!din_b[145] $ (((!din_a[147]) # (!din_b[146]))))) ) + ( Xd_0__inst_mult_24_105  ) + ( Xd_0__inst_mult_24_104  ))
// Xd_0__inst_mult_24_109  = SHARE((din_a[148] & (din_b[145] & (din_a[147] & din_b[146]))))

	.dataa(!din_a[148]),
	.datab(!din_b[145]),
	.datac(!din_a[147]),
	.datad(!din_b[146]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_104 ),
	.sharein(Xd_0__inst_mult_24_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_107 ),
	.cout(Xd_0__inst_mult_24_108 ),
	.shareout(Xd_0__inst_mult_24_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_31 (
// Equation(s):
// Xd_0__inst_mult_25_103  = SUM(( (!din_a[154] & (((din_a[153] & din_b[152])))) # (din_a[154] & (!din_b[151] $ (((!din_a[153]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_25_101  ) + ( Xd_0__inst_mult_25_100  ))
// Xd_0__inst_mult_25_104  = CARRY(( (!din_a[154] & (((din_a[153] & din_b[152])))) # (din_a[154] & (!din_b[151] $ (((!din_a[153]) # (!din_b[152]))))) ) + ( Xd_0__inst_mult_25_101  ) + ( Xd_0__inst_mult_25_100  ))
// Xd_0__inst_mult_25_105  = SHARE((din_a[154] & (din_b[151] & (din_a[153] & din_b[152]))))

	.dataa(!din_a[154]),
	.datab(!din_b[151]),
	.datac(!din_a[153]),
	.datad(!din_b[152]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_100 ),
	.sharein(Xd_0__inst_mult_25_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_103 ),
	.cout(Xd_0__inst_mult_25_104 ),
	.shareout(Xd_0__inst_mult_25_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_32 (
// Equation(s):
// Xd_0__inst_mult_22_107  = SUM(( (!din_a[136] & (((din_a[135] & din_b[134])))) # (din_a[136] & (!din_b[133] $ (((!din_a[135]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_22_105  ) + ( Xd_0__inst_mult_22_104  ))
// Xd_0__inst_mult_22_108  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[134])))) # (din_a[136] & (!din_b[133] $ (((!din_a[135]) # (!din_b[134]))))) ) + ( Xd_0__inst_mult_22_105  ) + ( Xd_0__inst_mult_22_104  ))
// Xd_0__inst_mult_22_109  = SHARE((din_a[136] & (din_b[133] & (din_a[135] & din_b[134]))))

	.dataa(!din_a[136]),
	.datab(!din_b[133]),
	.datac(!din_a[135]),
	.datad(!din_b[134]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_104 ),
	.sharein(Xd_0__inst_mult_22_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_107 ),
	.cout(Xd_0__inst_mult_22_108 ),
	.shareout(Xd_0__inst_mult_22_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_31 (
// Equation(s):
// Xd_0__inst_mult_23_103  = SUM(( (!din_a[142] & (((din_a[141] & din_b[140])))) # (din_a[142] & (!din_b[139] $ (((!din_a[141]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_23_101  ) + ( Xd_0__inst_mult_23_100  ))
// Xd_0__inst_mult_23_104  = CARRY(( (!din_a[142] & (((din_a[141] & din_b[140])))) # (din_a[142] & (!din_b[139] $ (((!din_a[141]) # (!din_b[140]))))) ) + ( Xd_0__inst_mult_23_101  ) + ( Xd_0__inst_mult_23_100  ))
// Xd_0__inst_mult_23_105  = SHARE((din_a[142] & (din_b[139] & (din_a[141] & din_b[140]))))

	.dataa(!din_a[142]),
	.datab(!din_b[139]),
	.datac(!din_a[141]),
	.datad(!din_b[140]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_100 ),
	.sharein(Xd_0__inst_mult_23_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_103 ),
	.cout(Xd_0__inst_mult_23_104 ),
	.shareout(Xd_0__inst_mult_23_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_31 (
// Equation(s):
// Xd_0__inst_mult_20_103  = SUM(( (!din_a[124] & (((din_a[123] & din_b[122])))) # (din_a[124] & (!din_b[121] $ (((!din_a[123]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_20_101  ) + ( Xd_0__inst_mult_20_100  ))
// Xd_0__inst_mult_20_104  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[122])))) # (din_a[124] & (!din_b[121] $ (((!din_a[123]) # (!din_b[122]))))) ) + ( Xd_0__inst_mult_20_101  ) + ( Xd_0__inst_mult_20_100  ))
// Xd_0__inst_mult_20_105  = SHARE((din_a[124] & (din_b[121] & (din_a[123] & din_b[122]))))

	.dataa(!din_a[124]),
	.datab(!din_b[121]),
	.datac(!din_a[123]),
	.datad(!din_b[122]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_100 ),
	.sharein(Xd_0__inst_mult_20_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_103 ),
	.cout(Xd_0__inst_mult_20_104 ),
	.shareout(Xd_0__inst_mult_20_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_30 (
// Equation(s):
// Xd_0__inst_mult_21_99  = SUM(( (!din_a[130] & (((din_a[129] & din_b[128])))) # (din_a[130] & (!din_b[127] $ (((!din_a[129]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_21_93  ) + ( Xd_0__inst_mult_21_92  ))
// Xd_0__inst_mult_21_100  = CARRY(( (!din_a[130] & (((din_a[129] & din_b[128])))) # (din_a[130] & (!din_b[127] $ (((!din_a[129]) # (!din_b[128]))))) ) + ( Xd_0__inst_mult_21_93  ) + ( Xd_0__inst_mult_21_92  ))
// Xd_0__inst_mult_21_101  = SHARE((din_a[130] & (din_b[127] & (din_a[129] & din_b[128]))))

	.dataa(!din_a[130]),
	.datab(!din_b[127]),
	.datac(!din_a[129]),
	.datad(!din_b[128]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_92 ),
	.sharein(Xd_0__inst_mult_21_93 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_99 ),
	.cout(Xd_0__inst_mult_21_100 ),
	.shareout(Xd_0__inst_mult_21_101 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_31 (
// Equation(s):
// Xd_0__inst_mult_21_103  = SUM(( GND ) + ( Xd_0__inst_mult_21_97  ) + ( Xd_0__inst_mult_21_96  ))
// Xd_0__inst_mult_21_104  = CARRY(( GND ) + ( Xd_0__inst_mult_21_97  ) + ( Xd_0__inst_mult_21_96  ))
// Xd_0__inst_mult_21_105  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_96 ),
	.sharein(Xd_0__inst_mult_21_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_103 ),
	.cout(Xd_0__inst_mult_21_104 ),
	.shareout(Xd_0__inst_mult_21_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_28 (
// Equation(s):
// Xd_0__inst_mult_18_90  = SUM(( (!din_a[112] & (((din_a[111] & din_b[110])))) # (din_a[112] & (!din_b[109] $ (((!din_a[111]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_18_84  ) + ( Xd_0__inst_mult_18_83  ))
// Xd_0__inst_mult_18_91  = CARRY(( (!din_a[112] & (((din_a[111] & din_b[110])))) # (din_a[112] & (!din_b[109] $ (((!din_a[111]) # (!din_b[110]))))) ) + ( Xd_0__inst_mult_18_84  ) + ( Xd_0__inst_mult_18_83  ))
// Xd_0__inst_mult_18_92  = SHARE((din_a[112] & (din_b[109] & (din_a[111] & din_b[110]))))

	.dataa(!din_a[112]),
	.datab(!din_b[109]),
	.datac(!din_a[111]),
	.datad(!din_b[110]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_83 ),
	.sharein(Xd_0__inst_mult_18_84 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_90 ),
	.cout(Xd_0__inst_mult_18_91 ),
	.shareout(Xd_0__inst_mult_18_92 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_29 (
// Equation(s):
// Xd_0__inst_mult_18_94  = SUM(( GND ) + ( Xd_0__inst_mult_18_88  ) + ( Xd_0__inst_mult_18_87  ))
// Xd_0__inst_mult_18_95  = CARRY(( GND ) + ( Xd_0__inst_mult_18_88  ) + ( Xd_0__inst_mult_18_87  ))
// Xd_0__inst_mult_18_96  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_87 ),
	.sharein(Xd_0__inst_mult_18_88 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_94 ),
	.cout(Xd_0__inst_mult_18_95 ),
	.shareout(Xd_0__inst_mult_18_96 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_32 (
// Equation(s):
// Xd_0__inst_mult_19_107  = SUM(( (!din_a[118] & (((din_a[117] & din_b[116])))) # (din_a[118] & (!din_b[115] $ (((!din_a[117]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_19_105  ) + ( Xd_0__inst_mult_19_104  ))
// Xd_0__inst_mult_19_108  = CARRY(( (!din_a[118] & (((din_a[117] & din_b[116])))) # (din_a[118] & (!din_b[115] $ (((!din_a[117]) # (!din_b[116]))))) ) + ( Xd_0__inst_mult_19_105  ) + ( Xd_0__inst_mult_19_104  ))
// Xd_0__inst_mult_19_109  = SHARE((din_a[118] & (din_b[115] & (din_a[117] & din_b[116]))))

	.dataa(!din_a[118]),
	.datab(!din_b[115]),
	.datac(!din_a[117]),
	.datad(!din_b[116]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_104 ),
	.sharein(Xd_0__inst_mult_19_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_107 ),
	.cout(Xd_0__inst_mult_19_108 ),
	.shareout(Xd_0__inst_mult_19_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_16_30 (
// Equation(s):
// Xd_0__inst_mult_16_98  = SUM(( (!din_a[100] & (((din_a[99] & din_b[99])))) # (din_a[100] & (!din_b[98] $ (((!din_a[99]) # (!din_b[99]))))) ) + ( Xd_0__inst_mult_16_92  ) + ( Xd_0__inst_mult_16_91  ))
// Xd_0__inst_mult_16_99  = CARRY(( (!din_a[100] & (((din_a[99] & din_b[99])))) # (din_a[100] & (!din_b[98] $ (((!din_a[99]) # (!din_b[99]))))) ) + ( Xd_0__inst_mult_16_92  ) + ( Xd_0__inst_mult_16_91  ))
// Xd_0__inst_mult_16_100  = SHARE((din_a[100] & (din_b[98] & (din_a[99] & din_b[99]))))

	.dataa(!din_a[100]),
	.datab(!din_b[98]),
	.datac(!din_a[99]),
	.datad(!din_b[99]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_91 ),
	.sharein(Xd_0__inst_mult_16_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_98 ),
	.cout(Xd_0__inst_mult_16_99 ),
	.shareout(Xd_0__inst_mult_16_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_17_32 (
// Equation(s):
// Xd_0__inst_mult_17_107  = SUM(( (!din_a[106] & (((din_a[105] & din_b[105])))) # (din_a[106] & (!din_b[104] $ (((!din_a[105]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_17_101  ) + ( Xd_0__inst_mult_17_100  ))
// Xd_0__inst_mult_17_108  = CARRY(( (!din_a[106] & (((din_a[105] & din_b[105])))) # (din_a[106] & (!din_b[104] $ (((!din_a[105]) # (!din_b[105]))))) ) + ( Xd_0__inst_mult_17_101  ) + ( Xd_0__inst_mult_17_100  ))
// Xd_0__inst_mult_17_109  = SHARE((din_a[106] & (din_b[104] & (din_a[105] & din_b[105]))))

	.dataa(!din_a[106]),
	.datab(!din_b[104]),
	.datac(!din_a[105]),
	.datad(!din_b[105]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_100 ),
	.sharein(Xd_0__inst_mult_17_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_107 ),
	.cout(Xd_0__inst_mult_17_108 ),
	.shareout(Xd_0__inst_mult_17_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_14_30 (
// Equation(s):
// Xd_0__inst_mult_14_98  = SUM(( (!din_a[88] & (((din_a[87] & din_b[87])))) # (din_a[88] & (!din_b[86] $ (((!din_a[87]) # (!din_b[87]))))) ) + ( Xd_0__inst_mult_14_92  ) + ( Xd_0__inst_mult_14_91  ))
// Xd_0__inst_mult_14_99  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[87])))) # (din_a[88] & (!din_b[86] $ (((!din_a[87]) # (!din_b[87]))))) ) + ( Xd_0__inst_mult_14_92  ) + ( Xd_0__inst_mult_14_91  ))
// Xd_0__inst_mult_14_100  = SHARE((din_a[88] & (din_b[86] & (din_a[87] & din_b[87]))))

	.dataa(!din_a[88]),
	.datab(!din_b[86]),
	.datac(!din_a[87]),
	.datad(!din_b[87]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_91 ),
	.sharein(Xd_0__inst_mult_14_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_98 ),
	.cout(Xd_0__inst_mult_14_99 ),
	.shareout(Xd_0__inst_mult_14_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_15_32 (
// Equation(s):
// Xd_0__inst_mult_15_107  = SUM(( (!din_a[94] & (((din_a[93] & din_b[93])))) # (din_a[94] & (!din_b[92] $ (((!din_a[93]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_15_101  ) + ( Xd_0__inst_mult_15_100  ))
// Xd_0__inst_mult_15_108  = CARRY(( (!din_a[94] & (((din_a[93] & din_b[93])))) # (din_a[94] & (!din_b[92] $ (((!din_a[93]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_15_101  ) + ( Xd_0__inst_mult_15_100  ))
// Xd_0__inst_mult_15_109  = SHARE((din_a[94] & (din_b[92] & (din_a[93] & din_b[93]))))

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(!din_a[93]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_100 ),
	.sharein(Xd_0__inst_mult_15_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_107 ),
	.cout(Xd_0__inst_mult_15_108 ),
	.shareout(Xd_0__inst_mult_15_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_12_31 (
// Equation(s):
// Xd_0__inst_mult_12_102  = SUM(( (!din_a[76] & (((din_a[75] & din_b[75])))) # (din_a[76] & (!din_b[74] $ (((!din_a[75]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_12_96  ) + ( Xd_0__inst_mult_12_95  ))
// Xd_0__inst_mult_12_103  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[75])))) # (din_a[76] & (!din_b[74] $ (((!din_a[75]) # (!din_b[75]))))) ) + ( Xd_0__inst_mult_12_96  ) + ( Xd_0__inst_mult_12_95  ))
// Xd_0__inst_mult_12_104  = SHARE((din_a[76] & (din_b[74] & (din_a[75] & din_b[75]))))

	.dataa(!din_a[76]),
	.datab(!din_b[74]),
	.datac(!din_a[75]),
	.datad(!din_b[75]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_95 ),
	.sharein(Xd_0__inst_mult_12_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_102 ),
	.cout(Xd_0__inst_mult_12_103 ),
	.shareout(Xd_0__inst_mult_12_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_13_31 (
// Equation(s):
// Xd_0__inst_mult_13_103  = SUM(( (!din_a[82] & (((din_a[81] & din_b[81])))) # (din_a[82] & (!din_b[80] $ (((!din_a[81]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_13_97  ) + ( Xd_0__inst_mult_13_96  ))
// Xd_0__inst_mult_13_104  = CARRY(( (!din_a[82] & (((din_a[81] & din_b[81])))) # (din_a[82] & (!din_b[80] $ (((!din_a[81]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_13_97  ) + ( Xd_0__inst_mult_13_96  ))
// Xd_0__inst_mult_13_105  = SHARE((din_a[82] & (din_b[80] & (din_a[81] & din_b[81]))))

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(!din_a[81]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_96 ),
	.sharein(Xd_0__inst_mult_13_97 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_103 ),
	.cout(Xd_0__inst_mult_13_104 ),
	.shareout(Xd_0__inst_mult_13_105 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_10_30 (
// Equation(s):
// Xd_0__inst_mult_10_98  = SUM(( (!din_a[64] & (((din_a[63] & din_b[63])))) # (din_a[64] & (!din_b[62] $ (((!din_a[63]) # (!din_b[63]))))) ) + ( Xd_0__inst_mult_10_92  ) + ( Xd_0__inst_mult_10_91  ))
// Xd_0__inst_mult_10_99  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[63])))) # (din_a[64] & (!din_b[62] $ (((!din_a[63]) # (!din_b[63]))))) ) + ( Xd_0__inst_mult_10_92  ) + ( Xd_0__inst_mult_10_91  ))
// Xd_0__inst_mult_10_100  = SHARE((din_a[64] & (din_b[62] & (din_a[63] & din_b[63]))))

	.dataa(!din_a[64]),
	.datab(!din_b[62]),
	.datac(!din_a[63]),
	.datad(!din_b[63]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_91 ),
	.sharein(Xd_0__inst_mult_10_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_98 ),
	.cout(Xd_0__inst_mult_10_99 ),
	.shareout(Xd_0__inst_mult_10_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_11_33 (
// Equation(s):
// Xd_0__inst_mult_11_111  = SUM(( (!din_a[70] & (((din_a[69] & din_b[69])))) # (din_a[70] & (!din_b[68] $ (((!din_a[69]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_11_109  ) + ( Xd_0__inst_mult_11_108  ))
// Xd_0__inst_mult_11_112  = CARRY(( (!din_a[70] & (((din_a[69] & din_b[69])))) # (din_a[70] & (!din_b[68] $ (((!din_a[69]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_11_109  ) + ( Xd_0__inst_mult_11_108  ))
// Xd_0__inst_mult_11_113  = SHARE((din_a[70] & (din_b[68] & (din_a[69] & din_b[69]))))

	.dataa(!din_a[70]),
	.datab(!din_b[68]),
	.datac(!din_a[69]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_108 ),
	.sharein(Xd_0__inst_mult_11_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_111 ),
	.cout(Xd_0__inst_mult_11_112 ),
	.shareout(Xd_0__inst_mult_11_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_8_31 (
// Equation(s):
// Xd_0__inst_mult_8_102  = SUM(( (!din_a[52] & (((din_a[51] & din_b[51])))) # (din_a[52] & (!din_b[50] $ (((!din_a[51]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_8_96  ) + ( Xd_0__inst_mult_8_95  ))
// Xd_0__inst_mult_8_103  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[51])))) # (din_a[52] & (!din_b[50] $ (((!din_a[51]) # (!din_b[51]))))) ) + ( Xd_0__inst_mult_8_96  ) + ( Xd_0__inst_mult_8_95  ))
// Xd_0__inst_mult_8_104  = SHARE((din_a[52] & (din_b[50] & (din_a[51] & din_b[51]))))

	.dataa(!din_a[52]),
	.datab(!din_b[50]),
	.datac(!din_a[51]),
	.datad(!din_b[51]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_95 ),
	.sharein(Xd_0__inst_mult_8_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_102 ),
	.cout(Xd_0__inst_mult_8_103 ),
	.shareout(Xd_0__inst_mult_8_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_9_32 (
// Equation(s):
// Xd_0__inst_mult_9_107  = SUM(( (!din_a[58] & (((din_a[57] & din_b[57])))) # (din_a[58] & (!din_b[56] $ (((!din_a[57]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_9_101  ) + ( Xd_0__inst_mult_9_100  ))
// Xd_0__inst_mult_9_108  = CARRY(( (!din_a[58] & (((din_a[57] & din_b[57])))) # (din_a[58] & (!din_b[56] $ (((!din_a[57]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_9_101  ) + ( Xd_0__inst_mult_9_100  ))
// Xd_0__inst_mult_9_109  = SHARE((din_a[58] & (din_b[56] & (din_a[57] & din_b[57]))))

	.dataa(!din_a[58]),
	.datab(!din_b[56]),
	.datac(!din_a[57]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_100 ),
	.sharein(Xd_0__inst_mult_9_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_107 ),
	.cout(Xd_0__inst_mult_9_108 ),
	.shareout(Xd_0__inst_mult_9_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_29 (
// Equation(s):
// Xd_0__inst_mult_6_93  = SUM(( (!din_a[40] & (((din_a[39] & din_b[39])))) # (din_a[40] & (!din_b[38] $ (((!din_a[39]) # (!din_b[39]))))) ) + ( Xd_0__inst_mult_6_91  ) + ( Xd_0__inst_mult_6_90  ))
// Xd_0__inst_mult_6_94  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[39])))) # (din_a[40] & (!din_b[38] $ (((!din_a[39]) # (!din_b[39]))))) ) + ( Xd_0__inst_mult_6_91  ) + ( Xd_0__inst_mult_6_90  ))
// Xd_0__inst_mult_6_95  = SHARE((din_a[40] & (din_b[38] & (din_a[39] & din_b[39]))))

	.dataa(!din_a[40]),
	.datab(!din_b[38]),
	.datac(!din_a[39]),
	.datad(!din_b[39]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_90 ),
	.sharein(Xd_0__inst_mult_6_91 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_93 ),
	.cout(Xd_0__inst_mult_6_94 ),
	.shareout(Xd_0__inst_mult_6_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_31 (
// Equation(s):
// Xd_0__inst_mult_7_102  = SUM(( (!din_a[46] & (((din_a[45] & din_b[45])))) # (din_a[46] & (!din_b[44] $ (((!din_a[45]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_7_100  ) + ( Xd_0__inst_mult_7_99  ))
// Xd_0__inst_mult_7_103  = CARRY(( (!din_a[46] & (((din_a[45] & din_b[45])))) # (din_a[46] & (!din_b[44] $ (((!din_a[45]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_7_100  ) + ( Xd_0__inst_mult_7_99  ))
// Xd_0__inst_mult_7_104  = SHARE((din_a[46] & (din_b[44] & (din_a[45] & din_b[45]))))

	.dataa(!din_a[46]),
	.datab(!din_b[44]),
	.datac(!din_a[45]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_99 ),
	.sharein(Xd_0__inst_mult_7_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_102 ),
	.cout(Xd_0__inst_mult_7_103 ),
	.shareout(Xd_0__inst_mult_7_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_29 (
// Equation(s):
// Xd_0__inst_mult_4_93  = SUM(( (!din_a[28] & (((din_a[27] & din_b[27])))) # (din_a[28] & (!din_b[26] $ (((!din_a[27]) # (!din_b[27]))))) ) + ( Xd_0__inst_mult_4_91  ) + ( Xd_0__inst_mult_4_90  ))
// Xd_0__inst_mult_4_94  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[27])))) # (din_a[28] & (!din_b[26] $ (((!din_a[27]) # (!din_b[27]))))) ) + ( Xd_0__inst_mult_4_91  ) + ( Xd_0__inst_mult_4_90  ))
// Xd_0__inst_mult_4_95  = SHARE((din_a[28] & (din_b[26] & (din_a[27] & din_b[27]))))

	.dataa(!din_a[28]),
	.datab(!din_b[26]),
	.datac(!din_a[27]),
	.datad(!din_b[27]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_90 ),
	.sharein(Xd_0__inst_mult_4_91 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_93 ),
	.cout(Xd_0__inst_mult_4_94 ),
	.shareout(Xd_0__inst_mult_4_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_30 (
// Equation(s):
// Xd_0__inst_mult_5_98  = SUM(( (!din_a[34] & (((din_a[33] & din_b[33])))) # (din_a[34] & (!din_b[32] $ (((!din_a[33]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_5_96  ) + ( Xd_0__inst_mult_5_95  ))
// Xd_0__inst_mult_5_99  = CARRY(( (!din_a[34] & (((din_a[33] & din_b[33])))) # (din_a[34] & (!din_b[32] $ (((!din_a[33]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_5_96  ) + ( Xd_0__inst_mult_5_95  ))
// Xd_0__inst_mult_5_100  = SHARE((din_a[34] & (din_b[32] & (din_a[33] & din_b[33]))))

	.dataa(!din_a[34]),
	.datab(!din_b[32]),
	.datac(!din_a[33]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_95 ),
	.sharein(Xd_0__inst_mult_5_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_98 ),
	.cout(Xd_0__inst_mult_5_99 ),
	.shareout(Xd_0__inst_mult_5_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_31 (
// Equation(s):
// Xd_0__inst_mult_2_102  = SUM(( (!din_a[16] & (((din_a[15] & din_b[15])))) # (din_a[16] & (!din_b[14] $ (((!din_a[15]) # (!din_b[15]))))) ) + ( Xd_0__inst_mult_2_100  ) + ( Xd_0__inst_mult_2_99  ))
// Xd_0__inst_mult_2_103  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[15])))) # (din_a[16] & (!din_b[14] $ (((!din_a[15]) # (!din_b[15]))))) ) + ( Xd_0__inst_mult_2_100  ) + ( Xd_0__inst_mult_2_99  ))
// Xd_0__inst_mult_2_104  = SHARE((din_a[16] & (din_b[14] & (din_a[15] & din_b[15]))))

	.dataa(!din_a[16]),
	.datab(!din_b[14]),
	.datac(!din_a[15]),
	.datad(!din_b[15]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_99 ),
	.sharein(Xd_0__inst_mult_2_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_102 ),
	.cout(Xd_0__inst_mult_2_103 ),
	.shareout(Xd_0__inst_mult_2_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_30 (
// Equation(s):
// Xd_0__inst_mult_3_98  = SUM(( (!din_a[22] & (((din_a[21] & din_b[21])))) # (din_a[22] & (!din_b[20] $ (((!din_a[21]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_3_96  ) + ( Xd_0__inst_mult_3_95  ))
// Xd_0__inst_mult_3_99  = CARRY(( (!din_a[22] & (((din_a[21] & din_b[21])))) # (din_a[22] & (!din_b[20] $ (((!din_a[21]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_3_96  ) + ( Xd_0__inst_mult_3_95  ))
// Xd_0__inst_mult_3_100  = SHARE((din_a[22] & (din_b[20] & (din_a[21] & din_b[21]))))

	.dataa(!din_a[22]),
	.datab(!din_b[20]),
	.datac(!din_a[21]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_95 ),
	.sharein(Xd_0__inst_mult_3_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_98 ),
	.cout(Xd_0__inst_mult_3_99 ),
	.shareout(Xd_0__inst_mult_3_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_31 (
// Equation(s):
// Xd_0__inst_mult_0_102  = SUM(( (!din_a[4] & (((din_a[3] & din_b[3])))) # (din_a[4] & (!din_b[2] $ (((!din_a[3]) # (!din_b[3]))))) ) + ( Xd_0__inst_mult_0_100  ) + ( Xd_0__inst_mult_0_99  ))
// Xd_0__inst_mult_0_103  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[3])))) # (din_a[4] & (!din_b[2] $ (((!din_a[3]) # (!din_b[3]))))) ) + ( Xd_0__inst_mult_0_100  ) + ( Xd_0__inst_mult_0_99  ))
// Xd_0__inst_mult_0_104  = SHARE((din_a[4] & (din_b[2] & (din_a[3] & din_b[3]))))

	.dataa(!din_a[4]),
	.datab(!din_b[2]),
	.datac(!din_a[3]),
	.datad(!din_b[3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_99 ),
	.sharein(Xd_0__inst_mult_0_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_102 ),
	.cout(Xd_0__inst_mult_0_103 ),
	.shareout(Xd_0__inst_mult_0_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_30 (
// Equation(s):
// Xd_0__inst_mult_1_98  = SUM(( (!din_a[10] & (((din_a[9] & din_b[9])))) # (din_a[10] & (!din_b[8] $ (((!din_a[9]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_96  ) + ( Xd_0__inst_mult_1_95  ))
// Xd_0__inst_mult_1_99  = CARRY(( (!din_a[10] & (((din_a[9] & din_b[9])))) # (din_a[10] & (!din_b[8] $ (((!din_a[9]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_1_96  ) + ( Xd_0__inst_mult_1_95  ))
// Xd_0__inst_mult_1_100  = SHARE((din_a[10] & (din_b[8] & (din_a[9] & din_b[9]))))

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(!din_a[9]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_95 ),
	.sharein(Xd_0__inst_mult_1_96 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_98 ),
	.cout(Xd_0__inst_mult_1_99 ),
	.shareout(Xd_0__inst_mult_1_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_28_32 (
// Equation(s):
// Xd_0__inst_mult_28_107  = SUM(( (!din_a[172] & (((din_a[171] & din_b[171])))) # (din_a[172] & (!din_b[170] $ (((!din_a[171]) # (!din_b[171]))))) ) + ( Xd_0__inst_mult_28_105  ) + ( Xd_0__inst_mult_28_104  ))
// Xd_0__inst_mult_28_108  = CARRY(( (!din_a[172] & (((din_a[171] & din_b[171])))) # (din_a[172] & (!din_b[170] $ (((!din_a[171]) # (!din_b[171]))))) ) + ( Xd_0__inst_mult_28_105  ) + ( Xd_0__inst_mult_28_104  ))
// Xd_0__inst_mult_28_109  = SHARE((din_a[172] & (din_b[170] & (din_a[171] & din_b[171]))))

	.dataa(!din_a[172]),
	.datab(!din_b[170]),
	.datac(!din_a[171]),
	.datad(!din_b[171]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_104 ),
	.sharein(Xd_0__inst_mult_28_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_107 ),
	.cout(Xd_0__inst_mult_28_108 ),
	.shareout(Xd_0__inst_mult_28_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_29_33 (
// Equation(s):
// Xd_0__inst_mult_29_111  = SUM(( (!din_a[178] & (((din_a[177] & din_b[177])))) # (din_a[178] & (!din_b[176] $ (((!din_a[177]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_29_109  ) + ( Xd_0__inst_mult_29_108  ))
// Xd_0__inst_mult_29_112  = CARRY(( (!din_a[178] & (((din_a[177] & din_b[177])))) # (din_a[178] & (!din_b[176] $ (((!din_a[177]) # (!din_b[177]))))) ) + ( Xd_0__inst_mult_29_109  ) + ( Xd_0__inst_mult_29_108  ))
// Xd_0__inst_mult_29_113  = SHARE((din_a[178] & (din_b[176] & (din_a[177] & din_b[177]))))

	.dataa(!din_a[178]),
	.datab(!din_b[176]),
	.datac(!din_a[177]),
	.datad(!din_b[177]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_108 ),
	.sharein(Xd_0__inst_mult_29_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_111 ),
	.cout(Xd_0__inst_mult_29_112 ),
	.shareout(Xd_0__inst_mult_29_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_26_33 (
// Equation(s):
// Xd_0__inst_mult_26_111  = SUM(( (!din_a[160] & (((din_a[159] & din_b[159])))) # (din_a[160] & (!din_b[158] $ (((!din_a[159]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_26_109  ) + ( Xd_0__inst_mult_26_108  ))
// Xd_0__inst_mult_26_112  = CARRY(( (!din_a[160] & (((din_a[159] & din_b[159])))) # (din_a[160] & (!din_b[158] $ (((!din_a[159]) # (!din_b[159]))))) ) + ( Xd_0__inst_mult_26_109  ) + ( Xd_0__inst_mult_26_108  ))
// Xd_0__inst_mult_26_113  = SHARE((din_a[160] & (din_b[158] & (din_a[159] & din_b[159]))))

	.dataa(!din_a[160]),
	.datab(!din_b[158]),
	.datac(!din_a[159]),
	.datad(!din_b[159]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_108 ),
	.sharein(Xd_0__inst_mult_26_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_111 ),
	.cout(Xd_0__inst_mult_26_112 ),
	.shareout(Xd_0__inst_mult_26_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_27_32 (
// Equation(s):
// Xd_0__inst_mult_27_107  = SUM(( (!din_a[166] & (((din_a[165] & din_b[165])))) # (din_a[166] & (!din_b[164] $ (((!din_a[165]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_27_105  ) + ( Xd_0__inst_mult_27_104  ))
// Xd_0__inst_mult_27_108  = CARRY(( (!din_a[166] & (((din_a[165] & din_b[165])))) # (din_a[166] & (!din_b[164] $ (((!din_a[165]) # (!din_b[165]))))) ) + ( Xd_0__inst_mult_27_105  ) + ( Xd_0__inst_mult_27_104  ))
// Xd_0__inst_mult_27_109  = SHARE((din_a[166] & (din_b[164] & (din_a[165] & din_b[165]))))

	.dataa(!din_a[166]),
	.datab(!din_b[164]),
	.datac(!din_a[165]),
	.datad(!din_b[165]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_104 ),
	.sharein(Xd_0__inst_mult_27_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_107 ),
	.cout(Xd_0__inst_mult_27_108 ),
	.shareout(Xd_0__inst_mult_27_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_24_33 (
// Equation(s):
// Xd_0__inst_mult_24_111  = SUM(( (!din_a[148] & (((din_a[147] & din_b[147])))) # (din_a[148] & (!din_b[146] $ (((!din_a[147]) # (!din_b[147]))))) ) + ( Xd_0__inst_mult_24_109  ) + ( Xd_0__inst_mult_24_108  ))
// Xd_0__inst_mult_24_112  = CARRY(( (!din_a[148] & (((din_a[147] & din_b[147])))) # (din_a[148] & (!din_b[146] $ (((!din_a[147]) # (!din_b[147]))))) ) + ( Xd_0__inst_mult_24_109  ) + ( Xd_0__inst_mult_24_108  ))
// Xd_0__inst_mult_24_113  = SHARE((din_a[148] & (din_b[146] & (din_a[147] & din_b[147]))))

	.dataa(!din_a[148]),
	.datab(!din_b[146]),
	.datac(!din_a[147]),
	.datad(!din_b[147]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_108 ),
	.sharein(Xd_0__inst_mult_24_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_111 ),
	.cout(Xd_0__inst_mult_24_112 ),
	.shareout(Xd_0__inst_mult_24_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_25_32 (
// Equation(s):
// Xd_0__inst_mult_25_107  = SUM(( (!din_a[154] & (((din_a[153] & din_b[153])))) # (din_a[154] & (!din_b[152] $ (((!din_a[153]) # (!din_b[153]))))) ) + ( Xd_0__inst_mult_25_105  ) + ( Xd_0__inst_mult_25_104  ))
// Xd_0__inst_mult_25_108  = CARRY(( (!din_a[154] & (((din_a[153] & din_b[153])))) # (din_a[154] & (!din_b[152] $ (((!din_a[153]) # (!din_b[153]))))) ) + ( Xd_0__inst_mult_25_105  ) + ( Xd_0__inst_mult_25_104  ))
// Xd_0__inst_mult_25_109  = SHARE((din_a[154] & (din_b[152] & (din_a[153] & din_b[153]))))

	.dataa(!din_a[154]),
	.datab(!din_b[152]),
	.datac(!din_a[153]),
	.datad(!din_b[153]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_104 ),
	.sharein(Xd_0__inst_mult_25_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_107 ),
	.cout(Xd_0__inst_mult_25_108 ),
	.shareout(Xd_0__inst_mult_25_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_22_33 (
// Equation(s):
// Xd_0__inst_mult_22_111  = SUM(( (!din_a[136] & (((din_a[135] & din_b[135])))) # (din_a[136] & (!din_b[134] $ (((!din_a[135]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_22_109  ) + ( Xd_0__inst_mult_22_108  ))
// Xd_0__inst_mult_22_112  = CARRY(( (!din_a[136] & (((din_a[135] & din_b[135])))) # (din_a[136] & (!din_b[134] $ (((!din_a[135]) # (!din_b[135]))))) ) + ( Xd_0__inst_mult_22_109  ) + ( Xd_0__inst_mult_22_108  ))
// Xd_0__inst_mult_22_113  = SHARE((din_a[136] & (din_b[134] & (din_a[135] & din_b[135]))))

	.dataa(!din_a[136]),
	.datab(!din_b[134]),
	.datac(!din_a[135]),
	.datad(!din_b[135]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_108 ),
	.sharein(Xd_0__inst_mult_22_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_111 ),
	.cout(Xd_0__inst_mult_22_112 ),
	.shareout(Xd_0__inst_mult_22_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_23_32 (
// Equation(s):
// Xd_0__inst_mult_23_107  = SUM(( (!din_a[142] & (((din_a[141] & din_b[141])))) # (din_a[142] & (!din_b[140] $ (((!din_a[141]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_23_105  ) + ( Xd_0__inst_mult_23_104  ))
// Xd_0__inst_mult_23_108  = CARRY(( (!din_a[142] & (((din_a[141] & din_b[141])))) # (din_a[142] & (!din_b[140] $ (((!din_a[141]) # (!din_b[141]))))) ) + ( Xd_0__inst_mult_23_105  ) + ( Xd_0__inst_mult_23_104  ))
// Xd_0__inst_mult_23_109  = SHARE((din_a[142] & (din_b[140] & (din_a[141] & din_b[141]))))

	.dataa(!din_a[142]),
	.datab(!din_b[140]),
	.datac(!din_a[141]),
	.datad(!din_b[141]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_104 ),
	.sharein(Xd_0__inst_mult_23_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_107 ),
	.cout(Xd_0__inst_mult_23_108 ),
	.shareout(Xd_0__inst_mult_23_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_20_32 (
// Equation(s):
// Xd_0__inst_mult_20_107  = SUM(( (!din_a[124] & (((din_a[123] & din_b[123])))) # (din_a[124] & (!din_b[122] $ (((!din_a[123]) # (!din_b[123]))))) ) + ( Xd_0__inst_mult_20_105  ) + ( Xd_0__inst_mult_20_104  ))
// Xd_0__inst_mult_20_108  = CARRY(( (!din_a[124] & (((din_a[123] & din_b[123])))) # (din_a[124] & (!din_b[122] $ (((!din_a[123]) # (!din_b[123]))))) ) + ( Xd_0__inst_mult_20_105  ) + ( Xd_0__inst_mult_20_104  ))
// Xd_0__inst_mult_20_109  = SHARE((din_a[124] & (din_b[122] & (din_a[123] & din_b[123]))))

	.dataa(!din_a[124]),
	.datab(!din_b[122]),
	.datac(!din_a[123]),
	.datad(!din_b[123]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_104 ),
	.sharein(Xd_0__inst_mult_20_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_107 ),
	.cout(Xd_0__inst_mult_20_108 ),
	.shareout(Xd_0__inst_mult_20_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_21_32 (
// Equation(s):
// Xd_0__inst_mult_21_107  = SUM(( (!din_a[130] & (((din_a[129] & din_b[129])))) # (din_a[130] & (!din_b[128] $ (((!din_a[129]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_21_101  ) + ( Xd_0__inst_mult_21_100  ))
// Xd_0__inst_mult_21_108  = CARRY(( (!din_a[130] & (((din_a[129] & din_b[129])))) # (din_a[130] & (!din_b[128] $ (((!din_a[129]) # (!din_b[129]))))) ) + ( Xd_0__inst_mult_21_101  ) + ( Xd_0__inst_mult_21_100  ))
// Xd_0__inst_mult_21_109  = SHARE((din_a[130] & (din_b[128] & (din_a[129] & din_b[129]))))

	.dataa(!din_a[130]),
	.datab(!din_b[128]),
	.datac(!din_a[129]),
	.datad(!din_b[129]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_100 ),
	.sharein(Xd_0__inst_mult_21_101 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_107 ),
	.cout(Xd_0__inst_mult_21_108 ),
	.shareout(Xd_0__inst_mult_21_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_18_30 (
// Equation(s):
// Xd_0__inst_mult_18_98  = SUM(( (!din_a[112] & (((din_a[111] & din_b[111])))) # (din_a[112] & (!din_b[110] $ (((!din_a[111]) # (!din_b[111]))))) ) + ( Xd_0__inst_mult_18_92  ) + ( Xd_0__inst_mult_18_91  ))
// Xd_0__inst_mult_18_99  = CARRY(( (!din_a[112] & (((din_a[111] & din_b[111])))) # (din_a[112] & (!din_b[110] $ (((!din_a[111]) # (!din_b[111]))))) ) + ( Xd_0__inst_mult_18_92  ) + ( Xd_0__inst_mult_18_91  ))
// Xd_0__inst_mult_18_100  = SHARE((din_a[112] & (din_b[110] & (din_a[111] & din_b[111]))))

	.dataa(!din_a[112]),
	.datab(!din_b[110]),
	.datac(!din_a[111]),
	.datad(!din_b[111]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_91 ),
	.sharein(Xd_0__inst_mult_18_92 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_98 ),
	.cout(Xd_0__inst_mult_18_99 ),
	.shareout(Xd_0__inst_mult_18_100 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_19_33 (
// Equation(s):
// Xd_0__inst_mult_19_111  = SUM(( (!din_a[118] & (((din_a[117] & din_b[117])))) # (din_a[118] & (!din_b[116] $ (((!din_a[117]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_19_109  ) + ( Xd_0__inst_mult_19_108  ))
// Xd_0__inst_mult_19_112  = CARRY(( (!din_a[118] & (((din_a[117] & din_b[117])))) # (din_a[118] & (!din_b[116] $ (((!din_a[117]) # (!din_b[117]))))) ) + ( Xd_0__inst_mult_19_109  ) + ( Xd_0__inst_mult_19_108  ))
// Xd_0__inst_mult_19_113  = SHARE((din_a[118] & (din_b[116] & (din_a[117] & din_b[117]))))

	.dataa(!din_a[118]),
	.datab(!din_b[116]),
	.datac(!din_a[117]),
	.datad(!din_b[117]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_108 ),
	.sharein(Xd_0__inst_mult_19_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_111 ),
	.cout(Xd_0__inst_mult_19_112 ),
	.shareout(Xd_0__inst_mult_19_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_16_31 (
// Equation(s):
// Xd_0__inst_mult_16_102  = SUM(( (din_a[100] & din_b[99]) ) + ( Xd_0__inst_mult_16_100  ) + ( Xd_0__inst_mult_16_99  ))
// Xd_0__inst_mult_16_103  = CARRY(( (din_a[100] & din_b[99]) ) + ( Xd_0__inst_mult_16_100  ) + ( Xd_0__inst_mult_16_99  ))
// Xd_0__inst_mult_16_104  = SHARE(GND)

	.dataa(!din_a[100]),
	.datab(!din_b[99]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_99 ),
	.sharein(Xd_0__inst_mult_16_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_102 ),
	.cout(Xd_0__inst_mult_16_103 ),
	.shareout(Xd_0__inst_mult_16_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_17_33 (
// Equation(s):
// Xd_0__inst_mult_17_111  = SUM(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_17_109  ) + ( Xd_0__inst_mult_17_108  ))
// Xd_0__inst_mult_17_112  = CARRY(( (din_a[106] & din_b[105]) ) + ( Xd_0__inst_mult_17_109  ) + ( Xd_0__inst_mult_17_108  ))
// Xd_0__inst_mult_17_113  = SHARE(GND)

	.dataa(!din_a[106]),
	.datab(!din_b[105]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_108 ),
	.sharein(Xd_0__inst_mult_17_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_17_111 ),
	.cout(Xd_0__inst_mult_17_112 ),
	.shareout(Xd_0__inst_mult_17_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_14_31 (
// Equation(s):
// Xd_0__inst_mult_14_102  = SUM(( (din_a[88] & din_b[87]) ) + ( Xd_0__inst_mult_14_100  ) + ( Xd_0__inst_mult_14_99  ))
// Xd_0__inst_mult_14_103  = CARRY(( (din_a[88] & din_b[87]) ) + ( Xd_0__inst_mult_14_100  ) + ( Xd_0__inst_mult_14_99  ))
// Xd_0__inst_mult_14_104  = SHARE(GND)

	.dataa(!din_a[88]),
	.datab(!din_b[87]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_99 ),
	.sharein(Xd_0__inst_mult_14_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_102 ),
	.cout(Xd_0__inst_mult_14_103 ),
	.shareout(Xd_0__inst_mult_14_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_15_33 (
// Equation(s):
// Xd_0__inst_mult_15_111  = SUM(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_15_109  ) + ( Xd_0__inst_mult_15_108  ))
// Xd_0__inst_mult_15_112  = CARRY(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_15_109  ) + ( Xd_0__inst_mult_15_108  ))
// Xd_0__inst_mult_15_113  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_15_108 ),
	.sharein(Xd_0__inst_mult_15_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_15_111 ),
	.cout(Xd_0__inst_mult_15_112 ),
	.shareout(Xd_0__inst_mult_15_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_12_32 (
// Equation(s):
// Xd_0__inst_mult_12_106  = SUM(( (din_a[76] & din_b[75]) ) + ( Xd_0__inst_mult_12_104  ) + ( Xd_0__inst_mult_12_103  ))
// Xd_0__inst_mult_12_107  = CARRY(( (din_a[76] & din_b[75]) ) + ( Xd_0__inst_mult_12_104  ) + ( Xd_0__inst_mult_12_103  ))
// Xd_0__inst_mult_12_108  = SHARE(GND)

	.dataa(!din_a[76]),
	.datab(!din_b[75]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_103 ),
	.sharein(Xd_0__inst_mult_12_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_12_106 ),
	.cout(Xd_0__inst_mult_12_107 ),
	.shareout(Xd_0__inst_mult_12_108 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_13_32 (
// Equation(s):
// Xd_0__inst_mult_13_107  = SUM(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_13_105  ) + ( Xd_0__inst_mult_13_104  ))
// Xd_0__inst_mult_13_108  = CARRY(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_13_105  ) + ( Xd_0__inst_mult_13_104  ))
// Xd_0__inst_mult_13_109  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_104 ),
	.sharein(Xd_0__inst_mult_13_105 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_107 ),
	.cout(Xd_0__inst_mult_13_108 ),
	.shareout(Xd_0__inst_mult_13_109 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_10_31 (
// Equation(s):
// Xd_0__inst_mult_10_102  = SUM(( (din_a[64] & din_b[63]) ) + ( Xd_0__inst_mult_10_100  ) + ( Xd_0__inst_mult_10_99  ))
// Xd_0__inst_mult_10_103  = CARRY(( (din_a[64] & din_b[63]) ) + ( Xd_0__inst_mult_10_100  ) + ( Xd_0__inst_mult_10_99  ))
// Xd_0__inst_mult_10_104  = SHARE(GND)

	.dataa(!din_a[64]),
	.datab(!din_b[63]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_99 ),
	.sharein(Xd_0__inst_mult_10_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_102 ),
	.cout(Xd_0__inst_mult_10_103 ),
	.shareout(Xd_0__inst_mult_10_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_11_34 (
// Equation(s):
// Xd_0__inst_mult_11_115  = SUM(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_11_113  ) + ( Xd_0__inst_mult_11_112  ))
// Xd_0__inst_mult_11_116  = CARRY(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_11_113  ) + ( Xd_0__inst_mult_11_112  ))
// Xd_0__inst_mult_11_117  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_11_112 ),
	.sharein(Xd_0__inst_mult_11_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_11_115 ),
	.cout(Xd_0__inst_mult_11_116 ),
	.shareout(Xd_0__inst_mult_11_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_8_32 (
// Equation(s):
// Xd_0__inst_mult_8_106  = SUM(( (din_a[52] & din_b[51]) ) + ( Xd_0__inst_mult_8_104  ) + ( Xd_0__inst_mult_8_103  ))
// Xd_0__inst_mult_8_107  = CARRY(( (din_a[52] & din_b[51]) ) + ( Xd_0__inst_mult_8_104  ) + ( Xd_0__inst_mult_8_103  ))
// Xd_0__inst_mult_8_108  = SHARE(GND)

	.dataa(!din_a[52]),
	.datab(!din_b[51]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_103 ),
	.sharein(Xd_0__inst_mult_8_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_8_106 ),
	.cout(Xd_0__inst_mult_8_107 ),
	.shareout(Xd_0__inst_mult_8_108 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_9_33 (
// Equation(s):
// Xd_0__inst_mult_9_111  = SUM(( (din_a[58] & din_b[57]) ) + ( Xd_0__inst_mult_9_109  ) + ( Xd_0__inst_mult_9_108  ))
// Xd_0__inst_mult_9_112  = CARRY(( (din_a[58] & din_b[57]) ) + ( Xd_0__inst_mult_9_109  ) + ( Xd_0__inst_mult_9_108  ))
// Xd_0__inst_mult_9_113  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_9_108 ),
	.sharein(Xd_0__inst_mult_9_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_9_111 ),
	.cout(Xd_0__inst_mult_9_112 ),
	.shareout(Xd_0__inst_mult_9_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_30 (
// Equation(s):
// Xd_0__inst_mult_6_97  = SUM(( (din_a[40] & din_b[39]) ) + ( Xd_0__inst_mult_6_95  ) + ( Xd_0__inst_mult_6_94  ))
// Xd_0__inst_mult_6_98  = CARRY(( (din_a[40] & din_b[39]) ) + ( Xd_0__inst_mult_6_95  ) + ( Xd_0__inst_mult_6_94  ))
// Xd_0__inst_mult_6_99  = SHARE(GND)

	.dataa(!din_a[40]),
	.datab(!din_b[39]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_94 ),
	.sharein(Xd_0__inst_mult_6_95 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_97 ),
	.cout(Xd_0__inst_mult_6_98 ),
	.shareout(Xd_0__inst_mult_6_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_32 (
// Equation(s):
// Xd_0__inst_mult_7_106  = SUM(( (din_a[46] & din_b[45]) ) + ( Xd_0__inst_mult_7_104  ) + ( Xd_0__inst_mult_7_103  ))
// Xd_0__inst_mult_7_107  = CARRY(( (din_a[46] & din_b[45]) ) + ( Xd_0__inst_mult_7_104  ) + ( Xd_0__inst_mult_7_103  ))
// Xd_0__inst_mult_7_108  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_103 ),
	.sharein(Xd_0__inst_mult_7_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_106 ),
	.cout(Xd_0__inst_mult_7_107 ),
	.shareout(Xd_0__inst_mult_7_108 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_30 (
// Equation(s):
// Xd_0__inst_mult_4_97  = SUM(( (din_a[28] & din_b[27]) ) + ( Xd_0__inst_mult_4_95  ) + ( Xd_0__inst_mult_4_94  ))
// Xd_0__inst_mult_4_98  = CARRY(( (din_a[28] & din_b[27]) ) + ( Xd_0__inst_mult_4_95  ) + ( Xd_0__inst_mult_4_94  ))
// Xd_0__inst_mult_4_99  = SHARE(GND)

	.dataa(!din_a[28]),
	.datab(!din_b[27]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_94 ),
	.sharein(Xd_0__inst_mult_4_95 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_97 ),
	.cout(Xd_0__inst_mult_4_98 ),
	.shareout(Xd_0__inst_mult_4_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_31 (
// Equation(s):
// Xd_0__inst_mult_5_102  = SUM(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_5_100  ) + ( Xd_0__inst_mult_5_99  ))
// Xd_0__inst_mult_5_103  = CARRY(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_5_100  ) + ( Xd_0__inst_mult_5_99  ))
// Xd_0__inst_mult_5_104  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_99 ),
	.sharein(Xd_0__inst_mult_5_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_102 ),
	.cout(Xd_0__inst_mult_5_103 ),
	.shareout(Xd_0__inst_mult_5_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_32 (
// Equation(s):
// Xd_0__inst_mult_2_106  = SUM(( (din_a[16] & din_b[15]) ) + ( Xd_0__inst_mult_2_104  ) + ( Xd_0__inst_mult_2_103  ))
// Xd_0__inst_mult_2_107  = CARRY(( (din_a[16] & din_b[15]) ) + ( Xd_0__inst_mult_2_104  ) + ( Xd_0__inst_mult_2_103  ))
// Xd_0__inst_mult_2_108  = SHARE(GND)

	.dataa(!din_a[16]),
	.datab(!din_b[15]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_103 ),
	.sharein(Xd_0__inst_mult_2_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_106 ),
	.cout(Xd_0__inst_mult_2_107 ),
	.shareout(Xd_0__inst_mult_2_108 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_31 (
// Equation(s):
// Xd_0__inst_mult_3_102  = SUM(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_3_100  ) + ( Xd_0__inst_mult_3_99  ))
// Xd_0__inst_mult_3_103  = CARRY(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_3_100  ) + ( Xd_0__inst_mult_3_99  ))
// Xd_0__inst_mult_3_104  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_99 ),
	.sharein(Xd_0__inst_mult_3_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_102 ),
	.cout(Xd_0__inst_mult_3_103 ),
	.shareout(Xd_0__inst_mult_3_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_32 (
// Equation(s):
// Xd_0__inst_mult_0_106  = SUM(( (din_a[4] & din_b[3]) ) + ( Xd_0__inst_mult_0_104  ) + ( Xd_0__inst_mult_0_103  ))
// Xd_0__inst_mult_0_107  = CARRY(( (din_a[4] & din_b[3]) ) + ( Xd_0__inst_mult_0_104  ) + ( Xd_0__inst_mult_0_103  ))
// Xd_0__inst_mult_0_108  = SHARE(GND)

	.dataa(!din_a[4]),
	.datab(!din_b[3]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_103 ),
	.sharein(Xd_0__inst_mult_0_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_106 ),
	.cout(Xd_0__inst_mult_0_107 ),
	.shareout(Xd_0__inst_mult_0_108 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_31 (
// Equation(s):
// Xd_0__inst_mult_1_102  = SUM(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_1_100  ) + ( Xd_0__inst_mult_1_99  ))
// Xd_0__inst_mult_1_103  = CARRY(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_1_100  ) + ( Xd_0__inst_mult_1_99  ))
// Xd_0__inst_mult_1_104  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_99 ),
	.sharein(Xd_0__inst_mult_1_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_102 ),
	.cout(Xd_0__inst_mult_1_103 ),
	.shareout(Xd_0__inst_mult_1_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_28_33 (
// Equation(s):
// Xd_0__inst_mult_28_111  = SUM(( (din_a[172] & din_b[171]) ) + ( Xd_0__inst_mult_28_109  ) + ( Xd_0__inst_mult_28_108  ))
// Xd_0__inst_mult_28_112  = CARRY(( (din_a[172] & din_b[171]) ) + ( Xd_0__inst_mult_28_109  ) + ( Xd_0__inst_mult_28_108  ))
// Xd_0__inst_mult_28_113  = SHARE(GND)

	.dataa(!din_a[172]),
	.datab(!din_b[171]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_108 ),
	.sharein(Xd_0__inst_mult_28_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_111 ),
	.cout(Xd_0__inst_mult_28_112 ),
	.shareout(Xd_0__inst_mult_28_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_29_34 (
// Equation(s):
// Xd_0__inst_mult_29_115  = SUM(( (din_a[178] & din_b[177]) ) + ( Xd_0__inst_mult_29_113  ) + ( Xd_0__inst_mult_29_112  ))
// Xd_0__inst_mult_29_116  = CARRY(( (din_a[178] & din_b[177]) ) + ( Xd_0__inst_mult_29_113  ) + ( Xd_0__inst_mult_29_112  ))
// Xd_0__inst_mult_29_117  = SHARE(GND)

	.dataa(!din_a[178]),
	.datab(!din_b[177]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_29_112 ),
	.sharein(Xd_0__inst_mult_29_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_29_115 ),
	.cout(Xd_0__inst_mult_29_116 ),
	.shareout(Xd_0__inst_mult_29_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_26_34 (
// Equation(s):
// Xd_0__inst_mult_26_115  = SUM(( (din_a[160] & din_b[159]) ) + ( Xd_0__inst_mult_26_113  ) + ( Xd_0__inst_mult_26_112  ))
// Xd_0__inst_mult_26_116  = CARRY(( (din_a[160] & din_b[159]) ) + ( Xd_0__inst_mult_26_113  ) + ( Xd_0__inst_mult_26_112  ))
// Xd_0__inst_mult_26_117  = SHARE(GND)

	.dataa(!din_a[160]),
	.datab(!din_b[159]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_26_112 ),
	.sharein(Xd_0__inst_mult_26_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_26_115 ),
	.cout(Xd_0__inst_mult_26_116 ),
	.shareout(Xd_0__inst_mult_26_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_27_33 (
// Equation(s):
// Xd_0__inst_mult_27_111  = SUM(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_27_109  ) + ( Xd_0__inst_mult_27_108  ))
// Xd_0__inst_mult_27_112  = CARRY(( (din_a[166] & din_b[165]) ) + ( Xd_0__inst_mult_27_109  ) + ( Xd_0__inst_mult_27_108  ))
// Xd_0__inst_mult_27_113  = SHARE(GND)

	.dataa(!din_a[166]),
	.datab(!din_b[165]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_108 ),
	.sharein(Xd_0__inst_mult_27_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_111 ),
	.cout(Xd_0__inst_mult_27_112 ),
	.shareout(Xd_0__inst_mult_27_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_24_34 (
// Equation(s):
// Xd_0__inst_mult_24_115  = SUM(( (din_a[148] & din_b[147]) ) + ( Xd_0__inst_mult_24_113  ) + ( Xd_0__inst_mult_24_112  ))
// Xd_0__inst_mult_24_116  = CARRY(( (din_a[148] & din_b[147]) ) + ( Xd_0__inst_mult_24_113  ) + ( Xd_0__inst_mult_24_112  ))
// Xd_0__inst_mult_24_117  = SHARE(GND)

	.dataa(!din_a[148]),
	.datab(!din_b[147]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_24_112 ),
	.sharein(Xd_0__inst_mult_24_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_24_115 ),
	.cout(Xd_0__inst_mult_24_116 ),
	.shareout(Xd_0__inst_mult_24_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_25_33 (
// Equation(s):
// Xd_0__inst_mult_25_111  = SUM(( (din_a[154] & din_b[153]) ) + ( Xd_0__inst_mult_25_109  ) + ( Xd_0__inst_mult_25_108  ))
// Xd_0__inst_mult_25_112  = CARRY(( (din_a[154] & din_b[153]) ) + ( Xd_0__inst_mult_25_109  ) + ( Xd_0__inst_mult_25_108  ))
// Xd_0__inst_mult_25_113  = SHARE(GND)

	.dataa(!din_a[154]),
	.datab(!din_b[153]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_108 ),
	.sharein(Xd_0__inst_mult_25_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_111 ),
	.cout(Xd_0__inst_mult_25_112 ),
	.shareout(Xd_0__inst_mult_25_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_22_34 (
// Equation(s):
// Xd_0__inst_mult_22_115  = SUM(( (din_a[136] & din_b[135]) ) + ( Xd_0__inst_mult_22_113  ) + ( Xd_0__inst_mult_22_112  ))
// Xd_0__inst_mult_22_116  = CARRY(( (din_a[136] & din_b[135]) ) + ( Xd_0__inst_mult_22_113  ) + ( Xd_0__inst_mult_22_112  ))
// Xd_0__inst_mult_22_117  = SHARE(GND)

	.dataa(!din_a[136]),
	.datab(!din_b[135]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_22_112 ),
	.sharein(Xd_0__inst_mult_22_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_22_115 ),
	.cout(Xd_0__inst_mult_22_116 ),
	.shareout(Xd_0__inst_mult_22_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_23_33 (
// Equation(s):
// Xd_0__inst_mult_23_111  = SUM(( (din_a[142] & din_b[141]) ) + ( Xd_0__inst_mult_23_109  ) + ( Xd_0__inst_mult_23_108  ))
// Xd_0__inst_mult_23_112  = CARRY(( (din_a[142] & din_b[141]) ) + ( Xd_0__inst_mult_23_109  ) + ( Xd_0__inst_mult_23_108  ))
// Xd_0__inst_mult_23_113  = SHARE(GND)

	.dataa(!din_a[142]),
	.datab(!din_b[141]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_108 ),
	.sharein(Xd_0__inst_mult_23_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_111 ),
	.cout(Xd_0__inst_mult_23_112 ),
	.shareout(Xd_0__inst_mult_23_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_20_33 (
// Equation(s):
// Xd_0__inst_mult_20_111  = SUM(( (din_a[124] & din_b[123]) ) + ( Xd_0__inst_mult_20_109  ) + ( Xd_0__inst_mult_20_108  ))
// Xd_0__inst_mult_20_112  = CARRY(( (din_a[124] & din_b[123]) ) + ( Xd_0__inst_mult_20_109  ) + ( Xd_0__inst_mult_20_108  ))
// Xd_0__inst_mult_20_113  = SHARE(GND)

	.dataa(!din_a[124]),
	.datab(!din_b[123]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_108 ),
	.sharein(Xd_0__inst_mult_20_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_111 ),
	.cout(Xd_0__inst_mult_20_112 ),
	.shareout(Xd_0__inst_mult_20_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_21_33 (
// Equation(s):
// Xd_0__inst_mult_21_111  = SUM(( (din_a[130] & din_b[129]) ) + ( Xd_0__inst_mult_21_109  ) + ( Xd_0__inst_mult_21_108  ))
// Xd_0__inst_mult_21_112  = CARRY(( (din_a[130] & din_b[129]) ) + ( Xd_0__inst_mult_21_109  ) + ( Xd_0__inst_mult_21_108  ))
// Xd_0__inst_mult_21_113  = SHARE(GND)

	.dataa(!din_a[130]),
	.datab(!din_b[129]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_108 ),
	.sharein(Xd_0__inst_mult_21_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_21_111 ),
	.cout(Xd_0__inst_mult_21_112 ),
	.shareout(Xd_0__inst_mult_21_113 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_18_31 (
// Equation(s):
// Xd_0__inst_mult_18_102  = SUM(( (din_a[112] & din_b[111]) ) + ( Xd_0__inst_mult_18_100  ) + ( Xd_0__inst_mult_18_99  ))
// Xd_0__inst_mult_18_103  = CARRY(( (din_a[112] & din_b[111]) ) + ( Xd_0__inst_mult_18_100  ) + ( Xd_0__inst_mult_18_99  ))
// Xd_0__inst_mult_18_104  = SHARE(GND)

	.dataa(!din_a[112]),
	.datab(!din_b[111]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_99 ),
	.sharein(Xd_0__inst_mult_18_100 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_102 ),
	.cout(Xd_0__inst_mult_18_103 ),
	.shareout(Xd_0__inst_mult_18_104 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_19_34 (
// Equation(s):
// Xd_0__inst_mult_19_115  = SUM(( (din_a[118] & din_b[117]) ) + ( Xd_0__inst_mult_19_113  ) + ( Xd_0__inst_mult_19_112  ))
// Xd_0__inst_mult_19_116  = CARRY(( (din_a[118] & din_b[117]) ) + ( Xd_0__inst_mult_19_113  ) + ( Xd_0__inst_mult_19_112  ))
// Xd_0__inst_mult_19_117  = SHARE(GND)

	.dataa(!din_a[118]),
	.datab(!din_b[117]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_19_112 ),
	.sharein(Xd_0__inst_mult_19_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_19_115 ),
	.cout(Xd_0__inst_mult_19_116 ),
	.shareout(Xd_0__inst_mult_19_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_32 (
// Equation(s):
// Xd_0__inst_mult_16_106  = SUM(( GND ) + ( Xd_0__inst_mult_16_104  ) + ( Xd_0__inst_mult_16_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_103 ),
	.sharein(Xd_0__inst_mult_16_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_16_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_32 (
// Equation(s):
// Xd_0__inst_mult_14_106  = SUM(( GND ) + ( Xd_0__inst_mult_14_104  ) + ( Xd_0__inst_mult_14_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_103 ),
	.sharein(Xd_0__inst_mult_14_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_14_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_33 (
// Equation(s):
// Xd_0__inst_mult_13_111  = SUM(( GND ) + ( Xd_0__inst_mult_13_109  ) + ( Xd_0__inst_mult_13_108  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_108 ),
	.sharein(Xd_0__inst_mult_13_109 ),
	.combout(),
	.sumout(Xd_0__inst_mult_13_111 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_32 (
// Equation(s):
// Xd_0__inst_mult_10_106  = SUM(( GND ) + ( Xd_0__inst_mult_10_104  ) + ( Xd_0__inst_mult_10_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_103 ),
	.sharein(Xd_0__inst_mult_10_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_10_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_31 (
// Equation(s):
// Xd_0__inst_mult_6_101  = SUM(( GND ) + ( Xd_0__inst_mult_6_99  ) + ( Xd_0__inst_mult_6_98  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_98 ),
	.sharein(Xd_0__inst_mult_6_99 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_101 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_31 (
// Equation(s):
// Xd_0__inst_mult_4_101  = SUM(( GND ) + ( Xd_0__inst_mult_4_99  ) + ( Xd_0__inst_mult_4_98  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_98 ),
	.sharein(Xd_0__inst_mult_4_99 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_101 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_32 (
// Equation(s):
// Xd_0__inst_mult_5_106  = SUM(( GND ) + ( Xd_0__inst_mult_5_104  ) + ( Xd_0__inst_mult_5_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_103 ),
	.sharein(Xd_0__inst_mult_5_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_32 (
// Equation(s):
// Xd_0__inst_mult_3_106  = SUM(( GND ) + ( Xd_0__inst_mult_3_104  ) + ( Xd_0__inst_mult_3_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_103 ),
	.sharein(Xd_0__inst_mult_3_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_32 (
// Equation(s):
// Xd_0__inst_mult_1_106  = SUM(( GND ) + ( Xd_0__inst_mult_1_104  ) + ( Xd_0__inst_mult_1_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_103 ),
	.sharein(Xd_0__inst_mult_1_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_28_34 (
// Equation(s):
// Xd_0__inst_mult_28_115  = SUM(( GND ) + ( Xd_0__inst_mult_28_113  ) + ( Xd_0__inst_mult_28_112  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_28_112 ),
	.sharein(Xd_0__inst_mult_28_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_28_115 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_27_34 (
// Equation(s):
// Xd_0__inst_mult_27_115  = SUM(( GND ) + ( Xd_0__inst_mult_27_113  ) + ( Xd_0__inst_mult_27_112  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_27_112 ),
	.sharein(Xd_0__inst_mult_27_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_27_115 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_25_34 (
// Equation(s):
// Xd_0__inst_mult_25_115  = SUM(( GND ) + ( Xd_0__inst_mult_25_113  ) + ( Xd_0__inst_mult_25_112  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_25_112 ),
	.sharein(Xd_0__inst_mult_25_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_25_115 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_23_34 (
// Equation(s):
// Xd_0__inst_mult_23_115  = SUM(( GND ) + ( Xd_0__inst_mult_23_113  ) + ( Xd_0__inst_mult_23_112  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_23_112 ),
	.sharein(Xd_0__inst_mult_23_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_23_115 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_20_34 (
// Equation(s):
// Xd_0__inst_mult_20_115  = SUM(( GND ) + ( Xd_0__inst_mult_20_113  ) + ( Xd_0__inst_mult_20_112  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_20_112 ),
	.sharein(Xd_0__inst_mult_20_113 ),
	.combout(),
	.sumout(Xd_0__inst_mult_20_115 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_32 (
// Equation(s):
// Xd_0__inst_mult_18_106  = SUM(( GND ) + ( Xd_0__inst_mult_18_104  ) + ( Xd_0__inst_mult_18_103  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_103 ),
	.sharein(Xd_0__inst_mult_18_104 ),
	.combout(),
	.sumout(Xd_0__inst_mult_18_106 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_16_33 (
// Equation(s):
// Xd_0__inst_mult_16_111  = CARRY(( GND ) + ( Xd_0__inst_mult_18_96  ) + ( Xd_0__inst_mult_18_95  ))
// Xd_0__inst_mult_16_112  = SHARE((din_b[99] & din_a[97]))

	.dataa(!din_b[99]),
	.datab(!din_a[97]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_18_95 ),
	.sharein(Xd_0__inst_mult_18_96 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_16_111 ),
	.shareout(Xd_0__inst_mult_16_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_17_34 (
// Equation(s):
// Xd_0__inst_mult_17_116  = CARRY(( GND ) + ( Xd_0__inst_mult_16_96  ) + ( Xd_0__inst_mult_16_95  ))
// Xd_0__inst_mult_17_117  = SHARE((din_b[105] & din_a[103]))

	.dataa(!din_b[105]),
	.datab(!din_a[103]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_16_95 ),
	.sharein(Xd_0__inst_mult_16_96 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_17_116 ),
	.shareout(Xd_0__inst_mult_17_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_14_33 (
// Equation(s):
// Xd_0__inst_mult_14_111  = CARRY(( GND ) + ( Xd_0__inst_mult_17_105  ) + ( Xd_0__inst_mult_17_104  ))
// Xd_0__inst_mult_14_112  = SHARE((din_b[87] & din_a[85]))

	.dataa(!din_b[87]),
	.datab(!din_a[85]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_17_104 ),
	.sharein(Xd_0__inst_mult_17_105 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_14_111 ),
	.shareout(Xd_0__inst_mult_14_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_15_34 (
// Equation(s):
// Xd_0__inst_mult_15_116  = CARRY(( GND ) + ( Xd_0__inst_mult_14_96  ) + ( Xd_0__inst_mult_14_95  ))
// Xd_0__inst_mult_15_117  = SHARE((din_b[93] & din_a[91]))

	.dataa(!din_b[93]),
	.datab(!din_a[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_14_95 ),
	.sharein(Xd_0__inst_mult_14_96 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_15_116 ),
	.shareout(Xd_0__inst_mult_15_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_12_33 (
// Equation(s):
// Xd_0__inst_mult_12_111  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_12_112  = SHARE((din_b[75] & din_a[73]))

	.dataa(!din_b[75]),
	.datab(!din_a[73]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_12_111 ),
	.shareout(Xd_0__inst_mult_12_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_13_34 (
// Equation(s):
// Xd_0__inst_mult_13_116  = CARRY(( GND ) + ( Xd_0__inst_mult_12_100  ) + ( Xd_0__inst_mult_12_99  ))
// Xd_0__inst_mult_13_117  = SHARE((din_b[81] & din_a[79]))

	.dataa(!din_b[81]),
	.datab(!din_a[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_12_99 ),
	.sharein(Xd_0__inst_mult_12_100 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_13_116 ),
	.shareout(Xd_0__inst_mult_13_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_10_33 (
// Equation(s):
// Xd_0__inst_mult_10_111  = CARRY(( GND ) + ( Xd_0__inst_mult_13_101  ) + ( Xd_0__inst_mult_13_100  ))
// Xd_0__inst_mult_10_112  = SHARE((din_b[63] & din_a[61]))

	.dataa(!din_b[63]),
	.datab(!din_a[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_13_100 ),
	.sharein(Xd_0__inst_mult_13_101 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_10_111 ),
	.shareout(Xd_0__inst_mult_10_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_8_33 (
// Equation(s):
// Xd_0__inst_mult_8_111  = CARRY(( GND ) + ( Xd_0__inst_mult_21_105  ) + ( Xd_0__inst_mult_21_104  ))
// Xd_0__inst_mult_8_112  = SHARE((din_b[51] & din_a[49]))

	.dataa(!din_b[51]),
	.datab(!din_a[49]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_21_104 ),
	.sharein(Xd_0__inst_mult_21_105 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_8_111 ),
	.shareout(Xd_0__inst_mult_8_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_9_34 (
// Equation(s):
// Xd_0__inst_mult_9_116  = CARRY(( GND ) + ( Xd_0__inst_mult_8_100  ) + ( Xd_0__inst_mult_8_99  ))
// Xd_0__inst_mult_9_117  = SHARE((din_b[57] & din_a[55]))

	.dataa(!din_b[57]),
	.datab(!din_a[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_8_99 ),
	.sharein(Xd_0__inst_mult_8_100 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_9_116 ),
	.shareout(Xd_0__inst_mult_9_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_32 (
// Equation(s):
// Xd_0__inst_mult_6_106  = CARRY(( GND ) + ( Xd_0__inst_i17_123  ) + ( Xd_0__inst_i17_122  ))
// Xd_0__inst_mult_6_107  = SHARE((din_b[39] & din_a[37]))

	.dataa(!din_b[39]),
	.datab(!din_a[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_122 ),
	.sharein(Xd_0__inst_i17_123 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_106 ),
	.shareout(Xd_0__inst_mult_6_107 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_33 (
// Equation(s):
// Xd_0__inst_mult_7_111  = CARRY(( GND ) + ( Xd_0__inst_i17_127  ) + ( Xd_0__inst_i17_126  ))
// Xd_0__inst_mult_7_112  = SHARE((din_b[45] & din_a[43]))

	.dataa(!din_b[45]),
	.datab(!din_a[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_126 ),
	.sharein(Xd_0__inst_i17_127 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_111 ),
	.shareout(Xd_0__inst_mult_7_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_32 (
// Equation(s):
// Xd_0__inst_mult_4_106  = CARRY(( GND ) + ( Xd_0__inst_i17_23  ) + ( Xd_0__inst_i17_22  ))
// Xd_0__inst_mult_4_107  = SHARE((din_b[27] & din_a[25]))

	.dataa(!din_b[27]),
	.datab(!din_a[25]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_22 ),
	.sharein(Xd_0__inst_i17_23 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_106 ),
	.shareout(Xd_0__inst_mult_4_107 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_33 (
// Equation(s):
// Xd_0__inst_mult_5_111  = CARRY(( GND ) + ( Xd_0__inst_i17_15  ) + ( Xd_0__inst_i17_14  ))
// Xd_0__inst_mult_5_112  = SHARE((din_b[33] & din_a[31]))

	.dataa(!din_b[33]),
	.datab(!din_a[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_14 ),
	.sharein(Xd_0__inst_i17_15 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_111 ),
	.shareout(Xd_0__inst_mult_5_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_33 (
// Equation(s):
// Xd_0__inst_mult_2_111  = CARRY(( GND ) + ( Xd_0__inst_i17_83  ) + ( Xd_0__inst_i17_82  ))
// Xd_0__inst_mult_2_112  = SHARE((din_b[15] & din_a[13]))

	.dataa(!din_b[15]),
	.datab(!din_a[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_82 ),
	.sharein(Xd_0__inst_i17_83 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_111 ),
	.shareout(Xd_0__inst_mult_2_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_33 (
// Equation(s):
// Xd_0__inst_mult_3_111  = CARRY(( GND ) + ( Xd_0__inst_i17_79  ) + ( Xd_0__inst_i17_78  ))
// Xd_0__inst_mult_3_112  = SHARE((din_b[21] & din_a[19]))

	.dataa(!din_b[21]),
	.datab(!din_a[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_78 ),
	.sharein(Xd_0__inst_i17_79 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_111 ),
	.shareout(Xd_0__inst_mult_3_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_33 (
// Equation(s):
// Xd_0__inst_mult_0_111  = CARRY(( GND ) + ( Xd_0__inst_i17_75  ) + ( Xd_0__inst_i17_74  ))
// Xd_0__inst_mult_0_112  = SHARE((din_b[3] & din_a[1]))

	.dataa(!din_b[3]),
	.datab(!din_a[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_74 ),
	.sharein(Xd_0__inst_i17_75 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_111 ),
	.shareout(Xd_0__inst_mult_0_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_33 (
// Equation(s):
// Xd_0__inst_mult_1_111  = CARRY(( GND ) + ( Xd_0__inst_i17_71  ) + ( Xd_0__inst_i17_70  ))
// Xd_0__inst_mult_1_112  = SHARE((din_b[9] & din_a[7]))

	.dataa(!din_b[9]),
	.datab(!din_a[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i17_70 ),
	.sharein(Xd_0__inst_i17_71 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_111 ),
	.shareout(Xd_0__inst_mult_1_112 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_21_34 (
// Equation(s):
// Xd_0__inst_mult_21_116  = CARRY(( GND ) + ( Xd_0__inst_mult_10_96  ) + ( Xd_0__inst_mult_10_95  ))
// Xd_0__inst_mult_21_117  = SHARE((din_b[129] & din_a[127]))

	.dataa(!din_b[129]),
	.datab(!din_a[127]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_10_95 ),
	.sharein(Xd_0__inst_mult_10_96 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_21_116 ),
	.shareout(Xd_0__inst_mult_21_117 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_18_33 (
// Equation(s):
// Xd_0__inst_mult_18_111  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_18_112  = SHARE((din_b[111] & din_a[109]))

	.dataa(!din_b[111]),
	.datab(!din_a[109]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_18_111 ),
	.shareout(Xd_0__inst_mult_18_112 ));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_inst_dout [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_3_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_first_level_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__5__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__6__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__7__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__8__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__9__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__10__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_15__11__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_5__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_4_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_2_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_8_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_6_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_15__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_15__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_15__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_8__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_7__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_6__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_5__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_4__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_14__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_13__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_12__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_11__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_10__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_9__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_8__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_8__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_14__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_14__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_13__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_13__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_12__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_12__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_11__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_11__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_10__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_10__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_9__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_9__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_30_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [30]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_31_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [31]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_30__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_31__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_30__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_30__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_31__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_31__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(din_a[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(din_b[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_16_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_17_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_14_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_15_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_12_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_13_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_10_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_11_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_8_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_9_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_28_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [28]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_29_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [29]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_26_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [26]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_27_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [27]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_24_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_25_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_22_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_23_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_20_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_21_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_18_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_19_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_30_ (
	.clk(clk),
	.d(Xd_0__inst_i17_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [30]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_31_ (
	.clk(clk),
	.d(Xd_0__inst_i17_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [31]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_16__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_17__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_14__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_15__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_12__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_13__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_10__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_11__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_8__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_9__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_28__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_29__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_26__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_27__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_24__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_25__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_22__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_23__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_20__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_21__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_18__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_19__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_30__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_30_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_30__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_31__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_31_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_31__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_34 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_34 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_35 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_38 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_38 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_39 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_41 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_41 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_43 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_42 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_45 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_45 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_47 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_46 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_49 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_51 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_50 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_53 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_55 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_54 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_16__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_16__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_17__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_17__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_14__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_14__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_15__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_15__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_12__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_12__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_13__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_13__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_10__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_10__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_11__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_11__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_8__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_59 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_8__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_9__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_9__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_28__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_28__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_29__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_29__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_26__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_26__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_27__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_27__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_24__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_24__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_25__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_25__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_22__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_22__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_23__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_23__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_20__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_20__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_21__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_63 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_21__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_18__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_18__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_19__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_19__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(din_a[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(din_b[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_0 (
	.clk(clk),
	.d(din_a[153]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_1 (
	.clk(clk),
	.d(din_b[150]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_0 (
	.clk(clk),
	.d(din_a[147]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_1 (
	.clk(clk),
	.d(din_b[144]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_0 (
	.clk(clk),
	.d(din_a[165]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_1 (
	.clk(clk),
	.d(din_b[162]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_0 (
	.clk(clk),
	.d(din_a[159]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_1 (
	.clk(clk),
	.d(din_b[156]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_0 (
	.clk(clk),
	.d(din_a[177]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_1 (
	.clk(clk),
	.d(din_b[174]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_0 (
	.clk(clk),
	.d(din_a[171]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_1 (
	.clk(clk),
	.d(din_b[168]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_0 (
	.clk(clk),
	.d(din_a[189]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_1 (
	.clk(clk),
	.d(din_b[186]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_0 (
	.clk(clk),
	.d(din_a[123]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_1 (
	.clk(clk),
	.d(din_b[120]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(din_a[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(din_b[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(din_a[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(din_b[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_0 (
	.clk(clk),
	.d(din_a[69]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_1 (
	.clk(clk),
	.d(din_b[66]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_0 (
	.clk(clk),
	.d(din_a[183]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_1 (
	.clk(clk),
	.d(din_b[180]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_0 (
	.clk(clk),
	.d(din_a[141]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_1 (
	.clk(clk),
	.d(din_b[138]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_0 (
	.clk(clk),
	.d(din_a[135]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_1 (
	.clk(clk),
	.d(din_b[132]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_16_ (
	.clk(clk),
	.d(Xd_0__inst_i17_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_17_ (
	.clk(clk),
	.d(Xd_0__inst_i17_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_14_ (
	.clk(clk),
	.d(Xd_0__inst_i17_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_15_ (
	.clk(clk),
	.d(Xd_0__inst_i17_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_12_ (
	.clk(clk),
	.d(Xd_0__inst_i17_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_13_ (
	.clk(clk),
	.d(Xd_0__inst_i17_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_10_ (
	.clk(clk),
	.d(Xd_0__inst_i17_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_11_ (
	.clk(clk),
	.d(Xd_0__inst_i17_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_8_ (
	.clk(clk),
	.d(Xd_0__inst_i17_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_9_ (
	.clk(clk),
	.d(Xd_0__inst_i17_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_57 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i17_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i17_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_57 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i17_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i17_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i17_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i17_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i17_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i17_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_28_ (
	.clk(clk),
	.d(Xd_0__inst_i17_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [28]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_29_ (
	.clk(clk),
	.d(Xd_0__inst_i17_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [29]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_26_ (
	.clk(clk),
	.d(Xd_0__inst_i17_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [26]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_27_ (
	.clk(clk),
	.d(Xd_0__inst_i17_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [27]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_24_ (
	.clk(clk),
	.d(Xd_0__inst_i17_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_25_ (
	.clk(clk),
	.d(Xd_0__inst_i17_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_22_ (
	.clk(clk),
	.d(Xd_0__inst_i17_105_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_23_ (
	.clk(clk),
	.d(Xd_0__inst_i17_109_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_20_ (
	.clk(clk),
	.d(Xd_0__inst_i17_113_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_21_ (
	.clk(clk),
	.d(Xd_0__inst_i17_117_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_58 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_18_ (
	.clk(clk),
	.d(Xd_0__inst_i17_121_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_19_ (
	.clk(clk),
	.d(Xd_0__inst_i17_125_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_61 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_61 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_70 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_79 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_62 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_16__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_16_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_16__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_17__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_17_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_17__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_14__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_14_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_14__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_15__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_15_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_15__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_12__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_12_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_12__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_13__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_13_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_13__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_10__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_10_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_10__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_11__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_11_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_11__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_8__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_8_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_8__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_9__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_9_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_9__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_65 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_65 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_28__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_28_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_28__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_29__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_29_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_29__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_26__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_26_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_26__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_27__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_27_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_27__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_24__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_24_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_24__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_25__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_25_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_25__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_22__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_22_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_22__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_23__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_23_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_23__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_20__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_20_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_20__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_21__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_21_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_21__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_18__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_18_66 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_18__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_19__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_19_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_19__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_4 (
	.clk(clk),
	.d(din_b[184]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_2 (
	.clk(clk),
	.d(din_a[180]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_4 (
	.clk(clk),
	.d(din_b[190]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_2 (
	.clk(clk),
	.d(din_a[186]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_10 (
	.clk(clk),
	.d(din_a[181]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_67 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_10 (
	.clk(clk),
	.d(din_a[187]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_11 (
	.clk(clk),
	.d(din_a[182]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_11 (
	.clk(clk),
	.d(din_a[188]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_14 (
	.clk(clk),
	.d(din_a[184]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_30_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_14 (
	.clk(clk),
	.d(din_a[190]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_31_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_4 (
	.clk(clk),
	.d(din_b[100]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_2 (
	.clk(clk),
	.d(din_a[96]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_4 (
	.clk(clk),
	.d(din_b[106]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_2 (
	.clk(clk),
	.d(din_a[102]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_4 (
	.clk(clk),
	.d(din_b[88]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_2 (
	.clk(clk),
	.d(din_a[84]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_4 (
	.clk(clk),
	.d(din_b[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_2 (
	.clk(clk),
	.d(din_a[90]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_4 (
	.clk(clk),
	.d(din_b[76]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_2 (
	.clk(clk),
	.d(din_a[72]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_4 (
	.clk(clk),
	.d(din_b[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_2 (
	.clk(clk),
	.d(din_a[78]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_4 (
	.clk(clk),
	.d(din_b[64]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_2 (
	.clk(clk),
	.d(din_a[60]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_4 (
	.clk(clk),
	.d(din_b[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_2 (
	.clk(clk),
	.d(din_a[66]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_4 (
	.clk(clk),
	.d(din_b[52]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_2 (
	.clk(clk),
	.d(din_a[48]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_4 (
	.clk(clk),
	.d(din_b[58]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_2 (
	.clk(clk),
	.d(din_a[54]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(din_b[40]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(din_a[36]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_73 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(din_b[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(din_a[42]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(din_b[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(din_a[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_73 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(din_b[34]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(din_a[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(din_b[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(din_a[12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(din_b[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(din_a[18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(din_b[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(din_a[0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(din_b[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(din_a[6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_4 (
	.clk(clk),
	.d(din_b[172]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_2 (
	.clk(clk),
	.d(din_a[168]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_4 (
	.clk(clk),
	.d(din_b[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_2 (
	.clk(clk),
	.d(din_a[174]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_4 (
	.clk(clk),
	.d(din_b[160]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_2 (
	.clk(clk),
	.d(din_a[156]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_4 (
	.clk(clk),
	.d(din_b[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_2 (
	.clk(clk),
	.d(din_a[162]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_4 (
	.clk(clk),
	.d(din_b[148]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_2 (
	.clk(clk),
	.d(din_a[144]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_4 (
	.clk(clk),
	.d(din_b[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_2 (
	.clk(clk),
	.d(din_a[150]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_4 (
	.clk(clk),
	.d(din_b[136]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_2 (
	.clk(clk),
	.d(din_a[132]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_4 (
	.clk(clk),
	.d(din_b[142]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_2 (
	.clk(clk),
	.d(din_a[138]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_4 (
	.clk(clk),
	.d(din_b[124]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_2 (
	.clk(clk),
	.d(din_a[120]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_4 (
	.clk(clk),
	.d(din_b[130]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_2 (
	.clk(clk),
	.d(din_a[126]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_4 (
	.clk(clk),
	.d(din_b[112]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_2 (
	.clk(clk),
	.d(din_a[108]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_4 (
	.clk(clk),
	.d(din_b[118]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_2 (
	.clk(clk),
	.d(din_a[114]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_30_3 (
	.clk(clk),
	.d(din_b[183]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_30_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_31_3 (
	.clk(clk),
	.d(din_b[189]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_31_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_87 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_81 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_81 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_85 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_71 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_75 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_86 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_10 (
	.clk(clk),
	.d(din_a[97]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_10 (
	.clk(clk),
	.d(din_a[103]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_10 (
	.clk(clk),
	.d(din_a[85]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_10 (
	.clk(clk),
	.d(din_a[91]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_10 (
	.clk(clk),
	.d(din_a[73]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_10 (
	.clk(clk),
	.d(din_a[79]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_10 (
	.clk(clk),
	.d(din_a[61]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_10 (
	.clk(clk),
	.d(din_a[67]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_10 (
	.clk(clk),
	.d(din_a[49]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_10 (
	.clk(clk),
	.d(din_a[55]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(din_a[37]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(din_a[43]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_89 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(din_a[25]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(din_a[31]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_78 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(din_a[13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(din_a[19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_77 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(din_a[1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_77 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(din_a[7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_10 (
	.clk(clk),
	.d(din_a[169]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_10 (
	.clk(clk),
	.d(din_a[175]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_10 (
	.clk(clk),
	.d(din_a[157]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_10 (
	.clk(clk),
	.d(din_a[163]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_10 (
	.clk(clk),
	.d(din_a[145]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_40 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_10 (
	.clk(clk),
	.d(din_a[151]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_10 (
	.clk(clk),
	.d(din_a[133]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_10 (
	.clk(clk),
	.d(din_a[139]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_10 (
	.clk(clk),
	.d(din_a[121]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_99 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_10 (
	.clk(clk),
	.d(din_a[127]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_90 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_94 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_10 (
	.clk(clk),
	.d(din_a[109]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_36 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_10 (
	.clk(clk),
	.d(din_a[115]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_11 (
	.clk(clk),
	.d(din_a[98]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_11 (
	.clk(clk),
	.d(din_a[104]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_11 (
	.clk(clk),
	.d(din_a[86]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_11 (
	.clk(clk),
	.d(din_a[92]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_11 (
	.clk(clk),
	.d(din_a[74]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_11 (
	.clk(clk),
	.d(din_a[80]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_103 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_11 (
	.clk(clk),
	.d(din_a[62]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_11 (
	.clk(clk),
	.d(din_a[68]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_11 (
	.clk(clk),
	.d(din_a[50]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_11 (
	.clk(clk),
	.d(din_a[56]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(din_a[38]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(din_a[44]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(din_a[26]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_93 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(din_a[32]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(din_a[14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(din_a[20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(din_a[2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(din_a[8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_11 (
	.clk(clk),
	.d(din_a[170]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_11 (
	.clk(clk),
	.d(din_a[176]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_11 (
	.clk(clk),
	.d(din_a[158]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_11 (
	.clk(clk),
	.d(din_a[164]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_11 (
	.clk(clk),
	.d(din_a[146]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_11 (
	.clk(clk),
	.d(din_a[152]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_11 (
	.clk(clk),
	.d(din_a[134]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_11 (
	.clk(clk),
	.d(din_a[140]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_11 (
	.clk(clk),
	.d(din_a[122]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_11 (
	.clk(clk),
	.d(din_a[128]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_11 (
	.clk(clk),
	.d(din_a[110]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_98 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_11 (
	.clk(clk),
	.d(din_a[116]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_0 (
	.clk(clk),
	.d(din_a[99]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_0 (
	.clk(clk),
	.d(din_a[105]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_0 (
	.clk(clk),
	.d(din_a[87]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_0 (
	.clk(clk),
	.d(din_a[93]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_0 (
	.clk(clk),
	.d(din_a[75]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_0 (
	.clk(clk),
	.d(din_a[81]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_107 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_0 (
	.clk(clk),
	.d(din_a[63]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_0 (
	.clk(clk),
	.d(din_a[51]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_0 (
	.clk(clk),
	.d(din_a[57]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(din_a[39]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_97 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(din_a[45]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(din_a[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_97 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(din_a[33]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_0 (
	.clk(clk),
	.d(din_a[129]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_0 (
	.clk(clk),
	.d(din_a[111]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_102 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_0 (
	.clk(clk),
	.d(din_a[117]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_14 (
	.clk(clk),
	.d(din_a[100]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_16_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_14 (
	.clk(clk),
	.d(din_a[106]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_17_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_14 (
	.clk(clk),
	.d(din_a[88]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_14_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_14 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_15_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_14 (
	.clk(clk),
	.d(din_a[76]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_12_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_14 (
	.clk(clk),
	.d(din_a[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_13_111 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_14 (
	.clk(clk),
	.d(din_a[64]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_10_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_14 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_11_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_14 (
	.clk(clk),
	.d(din_a[52]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_8_74 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_14 (
	.clk(clk),
	.d(din_a[58]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_9_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(din_a[40]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_101 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(din_a[28]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_101 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(din_a[34]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(din_a[16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(din_a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(din_a[4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_82 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(din_a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_14 (
	.clk(clk),
	.d(din_a[172]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_28_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_14 (
	.clk(clk),
	.d(din_a[178]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_29_91 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_14 (
	.clk(clk),
	.d(din_a[160]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_26_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_14 (
	.clk(clk),
	.d(din_a[166]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_27_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_14 (
	.clk(clk),
	.d(din_a[148]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_24_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_14 (
	.clk(clk),
	.d(din_a[154]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_25_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_14 (
	.clk(clk),
	.d(din_a[136]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_22_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_14 (
	.clk(clk),
	.d(din_a[142]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_23_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_14 (
	.clk(clk),
	.d(din_a[124]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_20_115 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_14 (
	.clk(clk),
	.d(din_a[130]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_21_83 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_14 (
	.clk(clk),
	.d(din_a[112]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_18_106 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_14 (
	.clk(clk),
	.d(din_a[118]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_19_95 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_1 (
	.clk(clk),
	.d(din_b[102]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_1 (
	.clk(clk),
	.d(din_b[90]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_1 (
	.clk(clk),
	.d(din_b[78]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_1 (
	.clk(clk),
	.d(din_b[126]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_1 (
	.clk(clk),
	.d(din_b[54]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(din_b[42]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(din_b[30]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_1 (
	.clk(clk),
	.d(din_b[114]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_1 (
	.clk(clk),
	.d(din_b[96]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_16_3 (
	.clk(clk),
	.d(din_b[99]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_16_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_17_3 (
	.clk(clk),
	.d(din_b[105]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_17_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_1 (
	.clk(clk),
	.d(din_b[84]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_14_3 (
	.clk(clk),
	.d(din_b[87]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_14_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_15_3 (
	.clk(clk),
	.d(din_b[93]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_15_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_1 (
	.clk(clk),
	.d(din_b[72]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_12_3 (
	.clk(clk),
	.d(din_b[75]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_12_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_13_3 (
	.clk(clk),
	.d(din_b[81]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_13_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_1 (
	.clk(clk),
	.d(din_b[60]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_10_3 (
	.clk(clk),
	.d(din_b[63]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_10_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_11_3 (
	.clk(clk),
	.d(din_b[69]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_11_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_1 (
	.clk(clk),
	.d(din_b[48]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_8_3 (
	.clk(clk),
	.d(din_b[51]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_8_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_9_3 (
	.clk(clk),
	.d(din_b[57]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_9_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(din_b[36]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(din_b[39]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(din_b[45]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(din_b[24]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(din_b[27]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(din_b[33]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(din_b[15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(din_b[21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(din_b[3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(din_b[9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_28_3 (
	.clk(clk),
	.d(din_b[171]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_28_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_29_3 (
	.clk(clk),
	.d(din_b[177]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_29_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_26_3 (
	.clk(clk),
	.d(din_b[159]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_26_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_27_3 (
	.clk(clk),
	.d(din_b[165]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_27_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_24_3 (
	.clk(clk),
	.d(din_b[147]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_24_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_25_3 (
	.clk(clk),
	.d(din_b[153]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_25_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_22_3 (
	.clk(clk),
	.d(din_b[135]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_22_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_23_3 (
	.clk(clk),
	.d(din_b[141]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_23_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_20_3 (
	.clk(clk),
	.d(din_b[123]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_20_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_21_3 (
	.clk(clk),
	.d(din_b[129]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_21_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_1 (
	.clk(clk),
	.d(din_b[108]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_18_3 (
	.clk(clk),
	.d(din_b[111]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_18_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_19_3 (
	.clk(clk),
	.d(din_b[117]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_19_3_q ),
	.prn(vcc));

assign dout[0] = Xd_0__inst_inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_inst_dout [15];

endmodule
