// Copyright (C) 2018  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// VENDOR "Altera"
// PROGRAM "Quartus Prime"
// VERSION "Version 18.1.1 Internal Build 259 12/02/2018 SJ Pro Edition"

// DATE "12/08/2018 22:18:14"

// 
// Device: Altera 10AX115S2F45I1SG Package FBGA1932
// 

// 
// This Verilog file should be used for ModelSim (Verilog) only
// 

`timescale 1 ps/ 1 ps

module pe_dot_alm_a10_12x12x8 (
	dout,
	clk,
	din_a,
	din_b);
output 	[25:0] dout;
input 	clk;
input 	[95:0] din_a;
input 	[95:0] din_b;

wire gnd;
wire vcc;
wire unknown;

assign gnd = 1'b0;
assign vcc = 1'b1;
assign unknown = 1'bx;

tri1 devclrn;
tri1 devpor;
tri1 devoe;
wire Xd_0__inst_inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_inst_add_0_2 ;
wire Xd_0__inst_inst_inst_add_0_3 ;
wire Xd_0__inst_inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_inst_add_0_6 ;
wire Xd_0__inst_inst_inst_add_0_7 ;
wire Xd_0__inst_inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_inst_add_0_10 ;
wire Xd_0__inst_inst_inst_add_0_11 ;
wire Xd_0__inst_inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_inst_add_0_14 ;
wire Xd_0__inst_inst_inst_add_0_15 ;
wire Xd_0__inst_inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_inst_add_0_18 ;
wire Xd_0__inst_inst_inst_add_0_19 ;
wire Xd_0__inst_inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_inst_add_0_22 ;
wire Xd_0__inst_inst_inst_add_0_23 ;
wire Xd_0__inst_inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_inst_add_0_26 ;
wire Xd_0__inst_inst_inst_add_0_27 ;
wire Xd_0__inst_inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_inst_add_0_30 ;
wire Xd_0__inst_inst_inst_add_0_31 ;
wire Xd_0__inst_inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_inst_add_0_34 ;
wire Xd_0__inst_inst_inst_add_0_35 ;
wire Xd_0__inst_inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_inst_add_0_38 ;
wire Xd_0__inst_inst_inst_add_0_39 ;
wire Xd_0__inst_inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_inst_add_0_42 ;
wire Xd_0__inst_inst_inst_add_0_43 ;
wire Xd_0__inst_inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_inst_add_0_46 ;
wire Xd_0__inst_inst_inst_add_0_47 ;
wire Xd_0__inst_inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_inst_add_0_50 ;
wire Xd_0__inst_inst_inst_add_0_51 ;
wire Xd_0__inst_inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_inst_add_0_54 ;
wire Xd_0__inst_inst_inst_add_0_55 ;
wire Xd_0__inst_inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_inst_add_0_58 ;
wire Xd_0__inst_inst_inst_add_0_59 ;
wire Xd_0__inst_inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_inst_add_0_62 ;
wire Xd_0__inst_inst_inst_add_0_63 ;
wire Xd_0__inst_inst_inst_add_0_65_sumout ;
wire Xd_0__inst_inst_inst_add_0_66 ;
wire Xd_0__inst_inst_inst_add_0_67 ;
wire Xd_0__inst_inst_inst_add_0_69_sumout ;
wire Xd_0__inst_inst_inst_add_0_70 ;
wire Xd_0__inst_inst_inst_add_0_71 ;
wire Xd_0__inst_inst_inst_add_0_73_sumout ;
wire Xd_0__inst_inst_inst_add_0_74 ;
wire Xd_0__inst_inst_inst_add_0_75 ;
wire Xd_0__inst_inst_inst_add_0_77_sumout ;
wire Xd_0__inst_inst_inst_add_0_78 ;
wire Xd_0__inst_inst_inst_add_0_79 ;
wire Xd_0__inst_inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_inst_add_0_82 ;
wire Xd_0__inst_inst_inst_add_0_83 ;
wire Xd_0__inst_inst_inst_add_0_85_sumout ;
wire Xd_0__inst_inst_inst_add_0_86 ;
wire Xd_0__inst_inst_inst_add_0_87 ;
wire Xd_0__inst_inst_inst_add_0_89_sumout ;
wire Xd_0__inst_inst_inst_add_0_90 ;
wire Xd_0__inst_inst_inst_add_0_91 ;
wire Xd_0__inst_inst_inst_add_0_93_sumout ;
wire Xd_0__inst_inst_inst_add_0_94 ;
wire Xd_0__inst_inst_inst_add_0_95 ;
wire Xd_0__inst_inst_inst_add_0_97_sumout ;
wire Xd_0__inst_inst_inst_add_0_98 ;
wire Xd_0__inst_inst_inst_add_0_99 ;
wire Xd_0__inst_mult_1_169 ;
wire Xd_0__inst_mult_1_170 ;
wire Xd_0__inst_mult_1_171 ;
wire Xd_0__inst_mult_1_173 ;
wire Xd_0__inst_mult_1_174 ;
wire Xd_0__inst_mult_1_175 ;
wire Xd_0__inst_inst_add_0_1_sumout ;
wire Xd_0__inst_inst_add_0_2 ;
wire Xd_0__inst_inst_add_0_3 ;
wire Xd_0__inst_inst_add_0_5_sumout ;
wire Xd_0__inst_inst_add_0_6 ;
wire Xd_0__inst_inst_add_0_7 ;
wire Xd_0__inst_inst_add_0_9_sumout ;
wire Xd_0__inst_inst_add_0_10 ;
wire Xd_0__inst_inst_add_0_11 ;
wire Xd_0__inst_inst_add_0_13_sumout ;
wire Xd_0__inst_inst_add_0_14 ;
wire Xd_0__inst_inst_add_0_15 ;
wire Xd_0__inst_inst_add_0_17_sumout ;
wire Xd_0__inst_inst_add_0_18 ;
wire Xd_0__inst_inst_add_0_19 ;
wire Xd_0__inst_inst_add_0_21_sumout ;
wire Xd_0__inst_inst_add_0_22 ;
wire Xd_0__inst_inst_add_0_23 ;
wire Xd_0__inst_inst_add_0_25_sumout ;
wire Xd_0__inst_inst_add_0_26 ;
wire Xd_0__inst_inst_add_0_27 ;
wire Xd_0__inst_inst_add_0_29_sumout ;
wire Xd_0__inst_inst_add_0_30 ;
wire Xd_0__inst_inst_add_0_31 ;
wire Xd_0__inst_inst_add_0_33_sumout ;
wire Xd_0__inst_inst_add_0_34 ;
wire Xd_0__inst_inst_add_0_35 ;
wire Xd_0__inst_inst_add_0_37_sumout ;
wire Xd_0__inst_inst_add_0_38 ;
wire Xd_0__inst_inst_add_0_39 ;
wire Xd_0__inst_inst_add_0_41_sumout ;
wire Xd_0__inst_inst_add_0_42 ;
wire Xd_0__inst_inst_add_0_43 ;
wire Xd_0__inst_inst_add_0_45_sumout ;
wire Xd_0__inst_inst_add_0_46 ;
wire Xd_0__inst_inst_add_0_47 ;
wire Xd_0__inst_inst_add_0_49_sumout ;
wire Xd_0__inst_inst_add_0_50 ;
wire Xd_0__inst_inst_add_0_51 ;
wire Xd_0__inst_inst_add_0_53_sumout ;
wire Xd_0__inst_inst_add_0_54 ;
wire Xd_0__inst_inst_add_0_55 ;
wire Xd_0__inst_inst_add_0_57_sumout ;
wire Xd_0__inst_inst_add_0_58 ;
wire Xd_0__inst_inst_add_0_59 ;
wire Xd_0__inst_inst_add_0_61_sumout ;
wire Xd_0__inst_inst_add_0_62 ;
wire Xd_0__inst_inst_add_0_63 ;
wire Xd_0__inst_inst_add_0_65_sumout ;
wire Xd_0__inst_inst_add_0_66 ;
wire Xd_0__inst_inst_add_0_67 ;
wire Xd_0__inst_inst_add_0_69_sumout ;
wire Xd_0__inst_inst_add_0_70 ;
wire Xd_0__inst_inst_add_0_71 ;
wire Xd_0__inst_inst_add_0_73_sumout ;
wire Xd_0__inst_inst_add_0_74 ;
wire Xd_0__inst_inst_add_0_75 ;
wire Xd_0__inst_inst_add_0_77_sumout ;
wire Xd_0__inst_inst_add_0_78 ;
wire Xd_0__inst_inst_add_0_79 ;
wire Xd_0__inst_inst_add_0_81_sumout ;
wire Xd_0__inst_inst_add_0_82 ;
wire Xd_0__inst_inst_add_0_83 ;
wire Xd_0__inst_inst_add_0_85_sumout ;
wire Xd_0__inst_inst_add_0_86 ;
wire Xd_0__inst_inst_add_0_87 ;
wire Xd_0__inst_inst_add_0_89_sumout ;
wire Xd_0__inst_inst_add_0_90 ;
wire Xd_0__inst_inst_add_0_91 ;
wire Xd_0__inst_inst_add_0_93_sumout ;
wire Xd_0__inst_inst_add_0_94 ;
wire Xd_0__inst_inst_add_0_95 ;
wire Xd_0__inst_inst_add_0_97_sumout ;
wire Xd_0__inst_inst_add_0_98 ;
wire Xd_0__inst_inst_add_0_99 ;
wire Xd_0__inst_inst_add_0_101_sumout ;
wire Xd_0__inst_mult_1_176 ;
wire Xd_0__inst_mult_1_177 ;
wire Xd_0__inst_mult_1_178 ;
wire Xd_0__inst_mult_3_169 ;
wire Xd_0__inst_mult_3_170 ;
wire Xd_0__inst_mult_3_171 ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_mult_1_180 ;
wire Xd_0__inst_mult_1_181 ;
wire Xd_0__inst_mult_1_182 ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ;
wire Xd_0__inst_mult_3_173 ;
wire Xd_0__inst_mult_3_174 ;
wire Xd_0__inst_mult_3_175 ;
wire Xd_0__inst_mult_7_173 ;
wire Xd_0__inst_mult_7_174 ;
wire Xd_0__inst_mult_7_175 ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ;
wire Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ;
wire Xd_0__inst_mult_1_184 ;
wire Xd_0__inst_mult_1_185 ;
wire Xd_0__inst_mult_1_186 ;
wire Xd_0__inst_mult_3_176 ;
wire Xd_0__inst_mult_3_177 ;
wire Xd_0__inst_mult_3_178 ;
wire Xd_0__inst_mult_6_173 ;
wire Xd_0__inst_mult_6_174 ;
wire Xd_0__inst_mult_6_175 ;
wire Xd_0__inst_mult_0_169 ;
wire Xd_0__inst_mult_0_170 ;
wire Xd_0__inst_mult_0_171 ;
wire Xd_0__inst_mult_3_180 ;
wire Xd_0__inst_mult_3_181 ;
wire Xd_0__inst_mult_3_182 ;
wire Xd_0__inst_mult_7_177 ;
wire Xd_0__inst_mult_7_178 ;
wire Xd_0__inst_mult_7_179 ;
wire Xd_0__inst_mult_6_177 ;
wire Xd_0__inst_mult_6_178 ;
wire Xd_0__inst_mult_6_179 ;
wire Xd_0__inst_mult_7_180 ;
wire Xd_0__inst_mult_7_181 ;
wire Xd_0__inst_mult_7_182 ;
wire Xd_0__inst_mult_6_180 ;
wire Xd_0__inst_mult_6_181 ;
wire Xd_0__inst_mult_6_182 ;
wire Xd_0__inst_mult_7_184 ;
wire Xd_0__inst_mult_7_185 ;
wire Xd_0__inst_mult_7_186 ;
wire Xd_0__inst_mult_6_184 ;
wire Xd_0__inst_mult_6_185 ;
wire Xd_0__inst_mult_6_186 ;
wire Xd_0__inst_mult_7_188 ;
wire Xd_0__inst_mult_7_189 ;
wire Xd_0__inst_mult_7_190 ;
wire Xd_0__inst_mult_6_188 ;
wire Xd_0__inst_mult_6_189 ;
wire Xd_0__inst_mult_6_190 ;
wire Xd_0__inst_mult_7_192 ;
wire Xd_0__inst_mult_7_193 ;
wire Xd_0__inst_mult_7_194 ;
wire Xd_0__inst_mult_6_192 ;
wire Xd_0__inst_mult_6_193 ;
wire Xd_0__inst_mult_6_194 ;
wire Xd_0__inst_mult_7_196 ;
wire Xd_0__inst_mult_7_197 ;
wire Xd_0__inst_mult_7_198 ;
wire Xd_0__inst_mult_6_196 ;
wire Xd_0__inst_mult_6_197 ;
wire Xd_0__inst_mult_6_198 ;
wire Xd_0__inst_mult_7_200 ;
wire Xd_0__inst_mult_7_201 ;
wire Xd_0__inst_mult_7_202 ;
wire Xd_0__inst_mult_6_200 ;
wire Xd_0__inst_mult_6_201 ;
wire Xd_0__inst_mult_6_202 ;
wire Xd_0__inst_mult_7_204 ;
wire Xd_0__inst_mult_7_205 ;
wire Xd_0__inst_mult_7_206 ;
wire Xd_0__inst_mult_6_204 ;
wire Xd_0__inst_mult_6_205 ;
wire Xd_0__inst_mult_6_206 ;
wire Xd_0__inst_mult_7_208 ;
wire Xd_0__inst_mult_7_209 ;
wire Xd_0__inst_mult_7_210 ;
wire Xd_0__inst_mult_6_208 ;
wire Xd_0__inst_mult_6_209 ;
wire Xd_0__inst_mult_6_210 ;
wire Xd_0__inst_mult_7_212 ;
wire Xd_0__inst_mult_7_213 ;
wire Xd_0__inst_mult_7_214 ;
wire Xd_0__inst_mult_6_212 ;
wire Xd_0__inst_mult_6_213 ;
wire Xd_0__inst_mult_6_214 ;
wire Xd_0__inst_mult_7_216 ;
wire Xd_0__inst_mult_7_217 ;
wire Xd_0__inst_mult_7_218 ;
wire Xd_0__inst_mult_6_216 ;
wire Xd_0__inst_mult_6_217 ;
wire Xd_0__inst_mult_6_218 ;
wire Xd_0__inst_mult_7_220 ;
wire Xd_0__inst_mult_7_221 ;
wire Xd_0__inst_mult_7_222 ;
wire Xd_0__inst_mult_6_220 ;
wire Xd_0__inst_mult_6_221 ;
wire Xd_0__inst_mult_6_222 ;
wire Xd_0__inst_mult_7_224 ;
wire Xd_0__inst_mult_7_225 ;
wire Xd_0__inst_mult_7_226 ;
wire Xd_0__inst_mult_6_224 ;
wire Xd_0__inst_mult_6_225 ;
wire Xd_0__inst_mult_6_226 ;
wire Xd_0__inst_mult_7_228 ;
wire Xd_0__inst_mult_7_229 ;
wire Xd_0__inst_mult_7_230 ;
wire Xd_0__inst_mult_6_228 ;
wire Xd_0__inst_mult_6_229 ;
wire Xd_0__inst_mult_6_230 ;
wire Xd_0__inst_mult_7_232 ;
wire Xd_0__inst_mult_7_233 ;
wire Xd_0__inst_mult_7_234 ;
wire Xd_0__inst_mult_6_232 ;
wire Xd_0__inst_mult_6_233 ;
wire Xd_0__inst_mult_6_234 ;
wire Xd_0__inst_mult_7_236 ;
wire Xd_0__inst_mult_7_237 ;
wire Xd_0__inst_mult_7_238 ;
wire Xd_0__inst_mult_6_236 ;
wire Xd_0__inst_mult_6_237 ;
wire Xd_0__inst_mult_6_238 ;
wire Xd_0__inst_mult_7_240 ;
wire Xd_0__inst_mult_7_241 ;
wire Xd_0__inst_mult_7_242 ;
wire Xd_0__inst_mult_6_240 ;
wire Xd_0__inst_mult_7_244 ;
wire Xd_0__inst_mult_3_184 ;
wire Xd_0__inst_mult_3_185 ;
wire Xd_0__inst_mult_3_186 ;
wire Xd_0__inst_mult_6_244 ;
wire Xd_0__inst_mult_6_245 ;
wire Xd_0__inst_mult_6_246 ;
wire Xd_0__inst_mult_0_173 ;
wire Xd_0__inst_mult_0_174 ;
wire Xd_0__inst_mult_0_175 ;
wire Xd_0__inst_mult_3_188 ;
wire Xd_0__inst_mult_3_189 ;
wire Xd_0__inst_mult_3_190 ;
wire Xd_0__inst_mult_6_248 ;
wire Xd_0__inst_mult_6_249 ;
wire Xd_0__inst_mult_6_250 ;
wire Xd_0__inst_mult_7_248 ;
wire Xd_0__inst_mult_7_249 ;
wire Xd_0__inst_mult_7_250 ;
wire Xd_0__inst_i29_1_sumout ;
wire Xd_0__inst_i29_2 ;
wire Xd_0__inst_i29_3 ;
wire Xd_0__inst_i29_5_sumout ;
wire Xd_0__inst_i29_6 ;
wire Xd_0__inst_i29_7 ;
wire Xd_0__inst_mult_7_252 ;
wire Xd_0__inst_mult_7_256 ;
wire Xd_0__inst_mult_7_257 ;
wire Xd_0__inst_mult_7_258 ;
wire Xd_0__inst_mult_6_252 ;
wire Xd_0__inst_mult_6_253 ;
wire Xd_0__inst_mult_6_254 ;
wire Xd_0__inst_mult_7_260 ;
wire Xd_0__inst_mult_7_261 ;
wire Xd_0__inst_mult_7_262 ;
wire Xd_0__inst_mult_6_256 ;
wire Xd_0__inst_mult_6_257 ;
wire Xd_0__inst_mult_6_258 ;
wire Xd_0__inst_mult_7_264 ;
wire Xd_0__inst_mult_7_265 ;
wire Xd_0__inst_mult_7_266 ;
wire Xd_0__inst_mult_6_260 ;
wire Xd_0__inst_mult_6_261 ;
wire Xd_0__inst_mult_6_262 ;
wire Xd_0__inst_mult_7_268 ;
wire Xd_0__inst_mult_7_269 ;
wire Xd_0__inst_mult_7_270 ;
wire Xd_0__inst_mult_6_264 ;
wire Xd_0__inst_mult_6_265 ;
wire Xd_0__inst_mult_6_266 ;
wire Xd_0__inst_mult_7_272 ;
wire Xd_0__inst_mult_7_273 ;
wire Xd_0__inst_mult_7_274 ;
wire Xd_0__inst_mult_4_173 ;
wire Xd_0__inst_mult_4_174 ;
wire Xd_0__inst_mult_4_175 ;
wire Xd_0__inst_mult_5_173 ;
wire Xd_0__inst_mult_5_174 ;
wire Xd_0__inst_mult_5_175 ;
wire Xd_0__inst_mult_2_173 ;
wire Xd_0__inst_mult_2_174 ;
wire Xd_0__inst_mult_2_175 ;
wire Xd_0__inst_mult_3_192 ;
wire Xd_0__inst_mult_3_193 ;
wire Xd_0__inst_mult_3_194 ;
wire Xd_0__inst_mult_0_176 ;
wire Xd_0__inst_mult_0_177 ;
wire Xd_0__inst_mult_0_178 ;
wire Xd_0__inst_mult_1_188 ;
wire Xd_0__inst_mult_1_189 ;
wire Xd_0__inst_mult_1_190 ;
wire Xd_0__inst_mult_4_35_sumout ;
wire Xd_0__inst_mult_4_36 ;
wire Xd_0__inst_mult_4_37 ;
wire Xd_0__inst_mult_3_35_sumout ;
wire Xd_0__inst_mult_3_36 ;
wire Xd_0__inst_mult_3_37 ;
wire Xd_0__inst_mult_4_177 ;
wire Xd_0__inst_mult_4_178 ;
wire Xd_0__inst_mult_4_179 ;
wire Xd_0__inst_mult_5_177 ;
wire Xd_0__inst_mult_5_178 ;
wire Xd_0__inst_mult_5_179 ;
wire Xd_0__inst_mult_2_177 ;
wire Xd_0__inst_mult_2_178 ;
wire Xd_0__inst_mult_2_179 ;
wire Xd_0__inst_mult_3_196 ;
wire Xd_0__inst_mult_3_197 ;
wire Xd_0__inst_mult_3_198 ;
wire Xd_0__inst_mult_0_180 ;
wire Xd_0__inst_mult_0_181 ;
wire Xd_0__inst_mult_0_182 ;
wire Xd_0__inst_mult_1_192 ;
wire Xd_0__inst_mult_1_193 ;
wire Xd_0__inst_mult_1_194 ;
wire Xd_0__inst_mult_4_180 ;
wire Xd_0__inst_mult_4_181 ;
wire Xd_0__inst_mult_4_182 ;
wire Xd_0__inst_mult_5_180 ;
wire Xd_0__inst_mult_5_181 ;
wire Xd_0__inst_mult_5_182 ;
wire Xd_0__inst_mult_2_180 ;
wire Xd_0__inst_mult_2_181 ;
wire Xd_0__inst_mult_2_182 ;
wire Xd_0__inst_mult_3_200 ;
wire Xd_0__inst_mult_3_201 ;
wire Xd_0__inst_mult_3_202 ;
wire Xd_0__inst_mult_0_184 ;
wire Xd_0__inst_mult_0_185 ;
wire Xd_0__inst_mult_0_186 ;
wire Xd_0__inst_mult_1_196 ;
wire Xd_0__inst_mult_1_197 ;
wire Xd_0__inst_mult_1_198 ;
wire Xd_0__inst_mult_4_184 ;
wire Xd_0__inst_mult_4_185 ;
wire Xd_0__inst_mult_4_186 ;
wire Xd_0__inst_mult_5_184 ;
wire Xd_0__inst_mult_5_185 ;
wire Xd_0__inst_mult_5_186 ;
wire Xd_0__inst_mult_2_184 ;
wire Xd_0__inst_mult_2_185 ;
wire Xd_0__inst_mult_2_186 ;
wire Xd_0__inst_mult_3_204 ;
wire Xd_0__inst_mult_3_205 ;
wire Xd_0__inst_mult_3_206 ;
wire Xd_0__inst_mult_0_188 ;
wire Xd_0__inst_mult_0_189 ;
wire Xd_0__inst_mult_0_190 ;
wire Xd_0__inst_mult_1_200 ;
wire Xd_0__inst_mult_1_201 ;
wire Xd_0__inst_mult_1_202 ;
wire Xd_0__inst_mult_4_188 ;
wire Xd_0__inst_mult_4_189 ;
wire Xd_0__inst_mult_4_190 ;
wire Xd_0__inst_mult_5_188 ;
wire Xd_0__inst_mult_5_189 ;
wire Xd_0__inst_mult_5_190 ;
wire Xd_0__inst_mult_2_188 ;
wire Xd_0__inst_mult_2_189 ;
wire Xd_0__inst_mult_2_190 ;
wire Xd_0__inst_mult_3_208 ;
wire Xd_0__inst_mult_3_209 ;
wire Xd_0__inst_mult_3_210 ;
wire Xd_0__inst_mult_0_192 ;
wire Xd_0__inst_mult_0_193 ;
wire Xd_0__inst_mult_0_194 ;
wire Xd_0__inst_mult_1_204 ;
wire Xd_0__inst_mult_1_205 ;
wire Xd_0__inst_mult_1_206 ;
wire Xd_0__inst_mult_4_192 ;
wire Xd_0__inst_mult_4_193 ;
wire Xd_0__inst_mult_4_194 ;
wire Xd_0__inst_mult_5_192 ;
wire Xd_0__inst_mult_5_193 ;
wire Xd_0__inst_mult_5_194 ;
wire Xd_0__inst_mult_2_192 ;
wire Xd_0__inst_mult_2_193 ;
wire Xd_0__inst_mult_2_194 ;
wire Xd_0__inst_mult_3_212 ;
wire Xd_0__inst_mult_3_213 ;
wire Xd_0__inst_mult_3_214 ;
wire Xd_0__inst_mult_0_196 ;
wire Xd_0__inst_mult_0_197 ;
wire Xd_0__inst_mult_0_198 ;
wire Xd_0__inst_mult_1_208 ;
wire Xd_0__inst_mult_1_209 ;
wire Xd_0__inst_mult_1_210 ;
wire Xd_0__inst_mult_4_196 ;
wire Xd_0__inst_mult_4_197 ;
wire Xd_0__inst_mult_4_198 ;
wire Xd_0__inst_mult_5_196 ;
wire Xd_0__inst_mult_5_197 ;
wire Xd_0__inst_mult_5_198 ;
wire Xd_0__inst_mult_2_196 ;
wire Xd_0__inst_mult_2_197 ;
wire Xd_0__inst_mult_2_198 ;
wire Xd_0__inst_mult_3_216 ;
wire Xd_0__inst_mult_3_217 ;
wire Xd_0__inst_mult_3_218 ;
wire Xd_0__inst_mult_0_200 ;
wire Xd_0__inst_mult_0_201 ;
wire Xd_0__inst_mult_0_202 ;
wire Xd_0__inst_mult_1_212 ;
wire Xd_0__inst_mult_1_213 ;
wire Xd_0__inst_mult_1_214 ;
wire Xd_0__inst_mult_4_200 ;
wire Xd_0__inst_mult_4_201 ;
wire Xd_0__inst_mult_4_202 ;
wire Xd_0__inst_mult_5_200 ;
wire Xd_0__inst_mult_5_201 ;
wire Xd_0__inst_mult_5_202 ;
wire Xd_0__inst_mult_2_200 ;
wire Xd_0__inst_mult_2_201 ;
wire Xd_0__inst_mult_2_202 ;
wire Xd_0__inst_mult_3_220 ;
wire Xd_0__inst_mult_3_221 ;
wire Xd_0__inst_mult_3_222 ;
wire Xd_0__inst_mult_0_204 ;
wire Xd_0__inst_mult_0_205 ;
wire Xd_0__inst_mult_0_206 ;
wire Xd_0__inst_mult_1_216 ;
wire Xd_0__inst_mult_1_217 ;
wire Xd_0__inst_mult_1_218 ;
wire Xd_0__inst_mult_4_204 ;
wire Xd_0__inst_mult_4_205 ;
wire Xd_0__inst_mult_4_206 ;
wire Xd_0__inst_mult_5_204 ;
wire Xd_0__inst_mult_5_205 ;
wire Xd_0__inst_mult_5_206 ;
wire Xd_0__inst_mult_2_204 ;
wire Xd_0__inst_mult_2_205 ;
wire Xd_0__inst_mult_2_206 ;
wire Xd_0__inst_mult_3_224 ;
wire Xd_0__inst_mult_3_225 ;
wire Xd_0__inst_mult_3_226 ;
wire Xd_0__inst_mult_0_208 ;
wire Xd_0__inst_mult_0_209 ;
wire Xd_0__inst_mult_0_210 ;
wire Xd_0__inst_mult_1_220 ;
wire Xd_0__inst_mult_1_221 ;
wire Xd_0__inst_mult_1_222 ;
wire Xd_0__inst_mult_4_208 ;
wire Xd_0__inst_mult_4_209 ;
wire Xd_0__inst_mult_4_210 ;
wire Xd_0__inst_mult_5_208 ;
wire Xd_0__inst_mult_5_209 ;
wire Xd_0__inst_mult_5_210 ;
wire Xd_0__inst_mult_2_208 ;
wire Xd_0__inst_mult_2_209 ;
wire Xd_0__inst_mult_2_210 ;
wire Xd_0__inst_mult_3_228 ;
wire Xd_0__inst_mult_3_229 ;
wire Xd_0__inst_mult_3_230 ;
wire Xd_0__inst_mult_0_212 ;
wire Xd_0__inst_mult_0_213 ;
wire Xd_0__inst_mult_0_214 ;
wire Xd_0__inst_mult_1_224 ;
wire Xd_0__inst_mult_1_225 ;
wire Xd_0__inst_mult_1_226 ;
wire Xd_0__inst_mult_4_212 ;
wire Xd_0__inst_mult_4_213 ;
wire Xd_0__inst_mult_4_214 ;
wire Xd_0__inst_mult_5_212 ;
wire Xd_0__inst_mult_5_213 ;
wire Xd_0__inst_mult_5_214 ;
wire Xd_0__inst_mult_2_212 ;
wire Xd_0__inst_mult_2_213 ;
wire Xd_0__inst_mult_2_214 ;
wire Xd_0__inst_mult_3_232 ;
wire Xd_0__inst_mult_3_233 ;
wire Xd_0__inst_mult_3_234 ;
wire Xd_0__inst_mult_0_216 ;
wire Xd_0__inst_mult_0_217 ;
wire Xd_0__inst_mult_0_218 ;
wire Xd_0__inst_mult_1_228 ;
wire Xd_0__inst_mult_1_229 ;
wire Xd_0__inst_mult_1_230 ;
wire Xd_0__inst_mult_4_216 ;
wire Xd_0__inst_mult_4_217 ;
wire Xd_0__inst_mult_4_218 ;
wire Xd_0__inst_mult_5_216 ;
wire Xd_0__inst_mult_5_217 ;
wire Xd_0__inst_mult_5_218 ;
wire Xd_0__inst_mult_2_216 ;
wire Xd_0__inst_mult_2_217 ;
wire Xd_0__inst_mult_2_218 ;
wire Xd_0__inst_mult_3_236 ;
wire Xd_0__inst_mult_3_237 ;
wire Xd_0__inst_mult_3_238 ;
wire Xd_0__inst_mult_0_220 ;
wire Xd_0__inst_mult_0_221 ;
wire Xd_0__inst_mult_0_222 ;
wire Xd_0__inst_mult_1_232 ;
wire Xd_0__inst_mult_1_233 ;
wire Xd_0__inst_mult_1_234 ;
wire Xd_0__inst_mult_4_220 ;
wire Xd_0__inst_mult_4_221 ;
wire Xd_0__inst_mult_4_222 ;
wire Xd_0__inst_mult_5_220 ;
wire Xd_0__inst_mult_5_221 ;
wire Xd_0__inst_mult_5_222 ;
wire Xd_0__inst_mult_2_220 ;
wire Xd_0__inst_mult_2_221 ;
wire Xd_0__inst_mult_2_222 ;
wire Xd_0__inst_mult_3_240 ;
wire Xd_0__inst_mult_3_241 ;
wire Xd_0__inst_mult_3_242 ;
wire Xd_0__inst_mult_0_224 ;
wire Xd_0__inst_mult_0_225 ;
wire Xd_0__inst_mult_0_226 ;
wire Xd_0__inst_mult_1_236 ;
wire Xd_0__inst_mult_1_237 ;
wire Xd_0__inst_mult_1_238 ;
wire Xd_0__inst_mult_4_224 ;
wire Xd_0__inst_mult_4_225 ;
wire Xd_0__inst_mult_4_226 ;
wire Xd_0__inst_mult_5_224 ;
wire Xd_0__inst_mult_5_225 ;
wire Xd_0__inst_mult_5_226 ;
wire Xd_0__inst_mult_2_224 ;
wire Xd_0__inst_mult_2_225 ;
wire Xd_0__inst_mult_2_226 ;
wire Xd_0__inst_mult_3_244 ;
wire Xd_0__inst_mult_3_245 ;
wire Xd_0__inst_mult_3_246 ;
wire Xd_0__inst_mult_0_228 ;
wire Xd_0__inst_mult_0_229 ;
wire Xd_0__inst_mult_0_230 ;
wire Xd_0__inst_mult_1_240 ;
wire Xd_0__inst_mult_1_241 ;
wire Xd_0__inst_mult_1_242 ;
wire Xd_0__inst_mult_4_228 ;
wire Xd_0__inst_mult_4_229 ;
wire Xd_0__inst_mult_4_230 ;
wire Xd_0__inst_mult_5_228 ;
wire Xd_0__inst_mult_5_229 ;
wire Xd_0__inst_mult_5_230 ;
wire Xd_0__inst_mult_2_228 ;
wire Xd_0__inst_mult_2_229 ;
wire Xd_0__inst_mult_2_230 ;
wire Xd_0__inst_mult_3_248 ;
wire Xd_0__inst_mult_3_249 ;
wire Xd_0__inst_mult_3_250 ;
wire Xd_0__inst_mult_0_232 ;
wire Xd_0__inst_mult_0_233 ;
wire Xd_0__inst_mult_0_234 ;
wire Xd_0__inst_mult_1_244 ;
wire Xd_0__inst_mult_1_245 ;
wire Xd_0__inst_mult_1_246 ;
wire Xd_0__inst_mult_4_232 ;
wire Xd_0__inst_mult_4_233 ;
wire Xd_0__inst_mult_4_234 ;
wire Xd_0__inst_mult_5_232 ;
wire Xd_0__inst_mult_5_233 ;
wire Xd_0__inst_mult_5_234 ;
wire Xd_0__inst_mult_2_232 ;
wire Xd_0__inst_mult_2_233 ;
wire Xd_0__inst_mult_2_234 ;
wire Xd_0__inst_mult_3_252 ;
wire Xd_0__inst_mult_3_253 ;
wire Xd_0__inst_mult_3_254 ;
wire Xd_0__inst_mult_0_236 ;
wire Xd_0__inst_mult_0_237 ;
wire Xd_0__inst_mult_0_238 ;
wire Xd_0__inst_mult_1_248 ;
wire Xd_0__inst_mult_1_249 ;
wire Xd_0__inst_mult_1_250 ;
wire Xd_0__inst_mult_4_236 ;
wire Xd_0__inst_mult_5_236 ;
wire Xd_0__inst_mult_2_236 ;
wire Xd_0__inst_mult_3_256 ;
wire Xd_0__inst_mult_0_240 ;
wire Xd_0__inst_mult_1_252 ;
wire Xd_0__inst_mult_4_240 ;
wire Xd_0__inst_mult_4_241 ;
wire Xd_0__inst_mult_4_242 ;
wire Xd_0__inst_mult_5_240 ;
wire Xd_0__inst_mult_5_241 ;
wire Xd_0__inst_mult_5_242 ;
wire Xd_0__inst_i29_9_sumout ;
wire Xd_0__inst_i29_10 ;
wire Xd_0__inst_i29_11 ;
wire Xd_0__inst_i29_13_sumout ;
wire Xd_0__inst_i29_14 ;
wire Xd_0__inst_i29_15 ;
wire Xd_0__inst_mult_3_260 ;
wire Xd_0__inst_mult_3_264 ;
wire Xd_0__inst_mult_3_265 ;
wire Xd_0__inst_mult_3_266 ;
wire Xd_0__inst_mult_2_240 ;
wire Xd_0__inst_mult_2_241 ;
wire Xd_0__inst_mult_2_242 ;
wire Xd_0__inst_mult_3_268 ;
wire Xd_0__inst_mult_3_269 ;
wire Xd_0__inst_mult_3_270 ;
wire Xd_0__inst_i29_17_sumout ;
wire Xd_0__inst_i29_18 ;
wire Xd_0__inst_i29_19 ;
wire Xd_0__inst_i29_21_sumout ;
wire Xd_0__inst_i29_22 ;
wire Xd_0__inst_i29_23 ;
wire Xd_0__inst_mult_6_268 ;
wire Xd_0__inst_mult_6_272 ;
wire Xd_0__inst_mult_6_273 ;
wire Xd_0__inst_mult_6_274 ;
wire Xd_0__inst_mult_0_244 ;
wire Xd_0__inst_mult_0_245 ;
wire Xd_0__inst_mult_0_246 ;
wire Xd_0__inst_i29_25_sumout ;
wire Xd_0__inst_i29_26 ;
wire Xd_0__inst_i29_27 ;
wire Xd_0__inst_i29_29_sumout ;
wire Xd_0__inst_i29_30 ;
wire Xd_0__inst_i29_31 ;
wire Xd_0__inst_mult_0_248 ;
wire Xd_0__inst_mult_0_252 ;
wire Xd_0__inst_mult_0_253 ;
wire Xd_0__inst_mult_0_254 ;
wire Xd_0__inst_mult_3_272 ;
wire Xd_0__inst_mult_3_273 ;
wire Xd_0__inst_mult_3_274 ;
wire Xd_0__inst_mult_7_276 ;
wire Xd_0__inst_mult_7_277 ;
wire Xd_0__inst_mult_7_278 ;
wire Xd_0__inst_mult_7_280 ;
wire Xd_0__inst_mult_7_281 ;
wire Xd_0__inst_mult_7_282 ;
wire Xd_0__inst_mult_4_244 ;
wire Xd_0__inst_mult_4_245 ;
wire Xd_0__inst_mult_4_246 ;
wire Xd_0__inst_mult_5_244 ;
wire Xd_0__inst_mult_5_245 ;
wire Xd_0__inst_mult_5_246 ;
wire Xd_0__inst_mult_2_244 ;
wire Xd_0__inst_mult_2_245 ;
wire Xd_0__inst_mult_2_246 ;
wire Xd_0__inst_mult_3_276 ;
wire Xd_0__inst_mult_3_277 ;
wire Xd_0__inst_mult_3_278 ;
wire Xd_0__inst_mult_0_256 ;
wire Xd_0__inst_mult_0_257 ;
wire Xd_0__inst_mult_0_258 ;
wire Xd_0__inst_mult_4_248 ;
wire Xd_0__inst_mult_4_249 ;
wire Xd_0__inst_mult_4_250 ;
wire Xd_0__inst_mult_5_248 ;
wire Xd_0__inst_mult_5_249 ;
wire Xd_0__inst_mult_5_250 ;
wire Xd_0__inst_mult_2_248 ;
wire Xd_0__inst_mult_2_249 ;
wire Xd_0__inst_mult_2_250 ;
wire Xd_0__inst_mult_3_280 ;
wire Xd_0__inst_mult_3_281 ;
wire Xd_0__inst_mult_3_282 ;
wire Xd_0__inst_mult_0_260 ;
wire Xd_0__inst_mult_0_261 ;
wire Xd_0__inst_mult_0_262 ;
wire Xd_0__inst_mult_4_252 ;
wire Xd_0__inst_mult_4_253 ;
wire Xd_0__inst_mult_4_254 ;
wire Xd_0__inst_mult_5_252 ;
wire Xd_0__inst_mult_5_253 ;
wire Xd_0__inst_mult_5_254 ;
wire Xd_0__inst_mult_2_252 ;
wire Xd_0__inst_mult_2_253 ;
wire Xd_0__inst_mult_2_254 ;
wire Xd_0__inst_mult_3_284 ;
wire Xd_0__inst_mult_3_285 ;
wire Xd_0__inst_mult_3_286 ;
wire Xd_0__inst_mult_0_264 ;
wire Xd_0__inst_mult_0_265 ;
wire Xd_0__inst_mult_0_266 ;
wire Xd_0__inst_mult_1_256 ;
wire Xd_0__inst_mult_1_257 ;
wire Xd_0__inst_mult_1_258 ;
wire Xd_0__inst_mult_6_277 ;
wire Xd_0__inst_mult_6_278 ;
wire Xd_0__inst_mult_7_285 ;
wire Xd_0__inst_mult_7_286 ;
wire Xd_0__inst_mult_4_256 ;
wire Xd_0__inst_mult_4_257 ;
wire Xd_0__inst_mult_4_258 ;
wire Xd_0__inst_mult_5_256 ;
wire Xd_0__inst_mult_5_257 ;
wire Xd_0__inst_mult_5_258 ;
wire Xd_0__inst_mult_2_256 ;
wire Xd_0__inst_mult_2_257 ;
wire Xd_0__inst_mult_2_258 ;
wire Xd_0__inst_mult_3_288 ;
wire Xd_0__inst_mult_3_289 ;
wire Xd_0__inst_mult_3_290 ;
wire Xd_0__inst_mult_0_268 ;
wire Xd_0__inst_mult_0_269 ;
wire Xd_0__inst_mult_0_270 ;
wire Xd_0__inst_mult_1_260 ;
wire Xd_0__inst_mult_1_261 ;
wire Xd_0__inst_mult_1_262 ;
wire Xd_0__inst_mult_6_280 ;
wire Xd_0__inst_mult_6_281 ;
wire Xd_0__inst_mult_6_282 ;
wire Xd_0__inst_mult_6_284 ;
wire Xd_0__inst_mult_6_285 ;
wire Xd_0__inst_mult_6_286 ;
wire Xd_0__inst_mult_7_288 ;
wire Xd_0__inst_mult_7_289 ;
wire Xd_0__inst_mult_7_290 ;
wire Xd_0__inst_mult_7_292 ;
wire Xd_0__inst_mult_7_293 ;
wire Xd_0__inst_mult_7_294 ;
wire Xd_0__inst_mult_2_35_sumout ;
wire Xd_0__inst_mult_2_36 ;
wire Xd_0__inst_mult_2_37 ;
wire Xd_0__inst_mult_0_35_sumout ;
wire Xd_0__inst_mult_0_36 ;
wire Xd_0__inst_mult_0_37 ;
wire Xd_0__inst_mult_2_39_sumout ;
wire Xd_0__inst_mult_2_40 ;
wire Xd_0__inst_mult_2_41 ;
wire Xd_0__inst_mult_1_35_sumout ;
wire Xd_0__inst_mult_1_36 ;
wire Xd_0__inst_mult_1_37 ;
wire Xd_0__inst_mult_2_43_sumout ;
wire Xd_0__inst_mult_2_44 ;
wire Xd_0__inst_mult_2_45 ;
wire Xd_0__inst_mult_1_39_sumout ;
wire Xd_0__inst_mult_1_40 ;
wire Xd_0__inst_mult_1_41 ;
wire Xd_0__inst_mult_6_288 ;
wire Xd_0__inst_mult_6_289 ;
wire Xd_0__inst_mult_6_290 ;
wire Xd_0__inst_mult_6_292 ;
wire Xd_0__inst_mult_6_293 ;
wire Xd_0__inst_mult_6_294 ;
wire Xd_0__inst_mult_1_43_sumout ;
wire Xd_0__inst_mult_1_44 ;
wire Xd_0__inst_mult_1_45 ;
wire Xd_0__inst_mult_7_296 ;
wire Xd_0__inst_mult_7_297 ;
wire Xd_0__inst_mult_7_298 ;
wire Xd_0__inst_mult_7_300 ;
wire Xd_0__inst_mult_7_301 ;
wire Xd_0__inst_mult_7_302 ;
wire Xd_0__inst_mult_2_47_sumout ;
wire Xd_0__inst_mult_2_48 ;
wire Xd_0__inst_mult_2_49 ;
wire Xd_0__inst_mult_6_296 ;
wire Xd_0__inst_mult_6_297 ;
wire Xd_0__inst_mult_6_298 ;
wire Xd_0__inst_mult_6_300 ;
wire Xd_0__inst_mult_6_301 ;
wire Xd_0__inst_mult_6_302 ;
wire Xd_0__inst_mult_7_304 ;
wire Xd_0__inst_mult_7_305 ;
wire Xd_0__inst_mult_7_306 ;
wire Xd_0__inst_mult_7_308 ;
wire Xd_0__inst_mult_7_309 ;
wire Xd_0__inst_mult_7_310 ;
wire Xd_0__inst_mult_6_304 ;
wire Xd_0__inst_mult_6_305 ;
wire Xd_0__inst_mult_6_306 ;
wire Xd_0__inst_mult_6_308 ;
wire Xd_0__inst_mult_6_309 ;
wire Xd_0__inst_mult_6_310 ;
wire Xd_0__inst_mult_7_312 ;
wire Xd_0__inst_mult_7_313 ;
wire Xd_0__inst_mult_7_314 ;
wire Xd_0__inst_mult_7_316 ;
wire Xd_0__inst_mult_7_317 ;
wire Xd_0__inst_mult_7_318 ;
wire Xd_0__inst_mult_6_312 ;
wire Xd_0__inst_mult_6_313 ;
wire Xd_0__inst_mult_6_314 ;
wire Xd_0__inst_mult_6_316 ;
wire Xd_0__inst_mult_6_317 ;
wire Xd_0__inst_mult_6_318 ;
wire Xd_0__inst_mult_7_320 ;
wire Xd_0__inst_mult_7_321 ;
wire Xd_0__inst_mult_7_322 ;
wire Xd_0__inst_mult_7_324 ;
wire Xd_0__inst_mult_7_325 ;
wire Xd_0__inst_mult_7_326 ;
wire Xd_0__inst_mult_6_320 ;
wire Xd_0__inst_mult_6_321 ;
wire Xd_0__inst_mult_6_322 ;
wire Xd_0__inst_mult_6_324 ;
wire Xd_0__inst_mult_6_325 ;
wire Xd_0__inst_mult_6_326 ;
wire Xd_0__inst_mult_7_328 ;
wire Xd_0__inst_mult_7_329 ;
wire Xd_0__inst_mult_7_330 ;
wire Xd_0__inst_mult_7_332 ;
wire Xd_0__inst_mult_7_333 ;
wire Xd_0__inst_mult_7_334 ;
wire Xd_0__inst_mult_6_328 ;
wire Xd_0__inst_mult_6_329 ;
wire Xd_0__inst_mult_6_330 ;
wire Xd_0__inst_mult_6_332 ;
wire Xd_0__inst_mult_6_333 ;
wire Xd_0__inst_mult_6_334 ;
wire Xd_0__inst_mult_7_336 ;
wire Xd_0__inst_mult_7_337 ;
wire Xd_0__inst_mult_7_338 ;
wire Xd_0__inst_mult_7_340 ;
wire Xd_0__inst_mult_7_341 ;
wire Xd_0__inst_mult_7_342 ;
wire Xd_0__inst_mult_6_336 ;
wire Xd_0__inst_mult_6_337 ;
wire Xd_0__inst_mult_6_338 ;
wire Xd_0__inst_mult_6_340 ;
wire Xd_0__inst_mult_6_341 ;
wire Xd_0__inst_mult_6_342 ;
wire Xd_0__inst_mult_7_344 ;
wire Xd_0__inst_mult_7_345 ;
wire Xd_0__inst_mult_7_346 ;
wire Xd_0__inst_mult_7_348 ;
wire Xd_0__inst_mult_7_349 ;
wire Xd_0__inst_mult_7_350 ;
wire Xd_0__inst_mult_6_344 ;
wire Xd_0__inst_mult_6_345 ;
wire Xd_0__inst_mult_6_346 ;
wire Xd_0__inst_mult_6_348 ;
wire Xd_0__inst_mult_6_349 ;
wire Xd_0__inst_mult_6_350 ;
wire Xd_0__inst_mult_7_352 ;
wire Xd_0__inst_mult_7_353 ;
wire Xd_0__inst_mult_7_354 ;
wire Xd_0__inst_mult_6_352 ;
wire Xd_0__inst_mult_6_353 ;
wire Xd_0__inst_mult_6_354 ;
wire Xd_0__inst_mult_7_356 ;
wire Xd_0__inst_mult_7_357 ;
wire Xd_0__inst_mult_7_358 ;
wire Xd_0__inst_mult_6_356 ;
wire Xd_0__inst_mult_6_357 ;
wire Xd_0__inst_mult_6_358 ;
wire Xd_0__inst_mult_7_360 ;
wire Xd_0__inst_mult_7_361 ;
wire Xd_0__inst_mult_7_362 ;
wire Xd_0__inst_mult_6_360 ;
wire Xd_0__inst_mult_6_361 ;
wire Xd_0__inst_mult_6_362 ;
wire Xd_0__inst_mult_7_364 ;
wire Xd_0__inst_mult_7_365 ;
wire Xd_0__inst_mult_7_366 ;
wire Xd_0__inst_mult_6_364 ;
wire Xd_0__inst_mult_6_365 ;
wire Xd_0__inst_mult_6_366 ;
wire Xd_0__inst_mult_6_35_sumout ;
wire Xd_0__inst_mult_6_36 ;
wire Xd_0__inst_mult_6_37 ;
wire Xd_0__inst_mult_7_368 ;
wire Xd_0__inst_mult_7_369 ;
wire Xd_0__inst_mult_7_370 ;
wire Xd_0__inst_mult_7_35_sumout ;
wire Xd_0__inst_mult_7_36 ;
wire Xd_0__inst_mult_7_37 ;
wire Xd_0__inst_mult_6_368 ;
wire Xd_0__inst_mult_6_369 ;
wire Xd_0__inst_mult_6_370 ;
wire Xd_0__inst_mult_6_39_sumout ;
wire Xd_0__inst_mult_6_40 ;
wire Xd_0__inst_mult_6_41 ;
wire Xd_0__inst_mult_7_372 ;
wire Xd_0__inst_mult_7_373 ;
wire Xd_0__inst_mult_7_374 ;
wire Xd_0__inst_mult_7_39_sumout ;
wire Xd_0__inst_mult_7_40 ;
wire Xd_0__inst_mult_7_41 ;
wire Xd_0__inst_mult_6_372 ;
wire Xd_0__inst_mult_6_373 ;
wire Xd_0__inst_mult_6_374 ;
wire Xd_0__inst_mult_6_43_sumout ;
wire Xd_0__inst_mult_6_44 ;
wire Xd_0__inst_mult_6_45 ;
wire Xd_0__inst_mult_7_376 ;
wire Xd_0__inst_mult_7_377 ;
wire Xd_0__inst_mult_7_378 ;
wire Xd_0__inst_mult_7_43_sumout ;
wire Xd_0__inst_mult_7_44 ;
wire Xd_0__inst_mult_7_45 ;
wire Xd_0__inst_mult_6_376 ;
wire Xd_0__inst_mult_6_377 ;
wire Xd_0__inst_mult_6_378 ;
wire Xd_0__inst_mult_6_47_sumout ;
wire Xd_0__inst_mult_6_48 ;
wire Xd_0__inst_mult_6_49 ;
wire Xd_0__inst_mult_7_380 ;
wire Xd_0__inst_mult_7_381 ;
wire Xd_0__inst_mult_7_382 ;
wire Xd_0__inst_mult_7_47_sumout ;
wire Xd_0__inst_mult_7_48 ;
wire Xd_0__inst_mult_7_49 ;
wire Xd_0__inst_mult_6_380 ;
wire Xd_0__inst_mult_6_51_sumout ;
wire Xd_0__inst_mult_6_52 ;
wire Xd_0__inst_mult_6_53 ;
wire Xd_0__inst_mult_7_384 ;
wire Xd_0__inst_mult_7_51_sumout ;
wire Xd_0__inst_mult_7_52 ;
wire Xd_0__inst_mult_7_53 ;
wire Xd_0__inst_mult_3_292 ;
wire Xd_0__inst_mult_3_293 ;
wire Xd_0__inst_mult_3_294 ;
wire Xd_0__inst_mult_3_296 ;
wire Xd_0__inst_mult_3_297 ;
wire Xd_0__inst_mult_3_298 ;
wire Xd_0__inst_mult_6_384 ;
wire Xd_0__inst_mult_6_385 ;
wire Xd_0__inst_mult_6_386 ;
wire Xd_0__inst_mult_3_39_sumout ;
wire Xd_0__inst_mult_3_40 ;
wire Xd_0__inst_mult_3_41 ;
wire Xd_0__inst_mult_0_272 ;
wire Xd_0__inst_mult_0_273 ;
wire Xd_0__inst_mult_0_274 ;
wire Xd_0__inst_mult_0_276 ;
wire Xd_0__inst_mult_0_277 ;
wire Xd_0__inst_mult_0_278 ;
wire Xd_0__inst_mult_3_300 ;
wire Xd_0__inst_mult_3_301 ;
wire Xd_0__inst_mult_3_302 ;
wire Xd_0__inst_mult_7_388 ;
wire Xd_0__inst_mult_7_389 ;
wire Xd_0__inst_mult_7_390 ;
wire Xd_0__inst_mult_7_392 ;
wire Xd_0__inst_mult_4_261 ;
wire Xd_0__inst_mult_4_262 ;
wire Xd_0__inst_mult_5_261 ;
wire Xd_0__inst_mult_5_262 ;
wire Xd_0__inst_mult_2_261 ;
wire Xd_0__inst_mult_2_262 ;
wire Xd_0__inst_mult_3_305 ;
wire Xd_0__inst_mult_3_306 ;
wire Xd_0__inst_mult_0_281 ;
wire Xd_0__inst_mult_0_282 ;
wire Xd_0__inst_mult_1_265 ;
wire Xd_0__inst_mult_1_266 ;
wire Xd_0__inst_mult_6_388 ;
wire Xd_0__inst_mult_6_389 ;
wire Xd_0__inst_mult_6_390 ;
wire Xd_0__inst_mult_6_393 ;
wire Xd_0__inst_mult_6_394 ;
wire Xd_0__inst_mult_7_396 ;
wire Xd_0__inst_mult_7_397 ;
wire Xd_0__inst_mult_7_398 ;
wire Xd_0__inst_mult_7_401 ;
wire Xd_0__inst_mult_7_402 ;
wire Xd_0__inst_mult_4_264 ;
wire Xd_0__inst_mult_4_265 ;
wire Xd_0__inst_mult_4_266 ;
wire Xd_0__inst_mult_4_268 ;
wire Xd_0__inst_mult_4_269 ;
wire Xd_0__inst_mult_4_270 ;
wire Xd_0__inst_mult_5_264 ;
wire Xd_0__inst_mult_5_265 ;
wire Xd_0__inst_mult_5_266 ;
wire Xd_0__inst_mult_5_268 ;
wire Xd_0__inst_mult_5_269 ;
wire Xd_0__inst_mult_5_270 ;
wire Xd_0__inst_mult_2_264 ;
wire Xd_0__inst_mult_2_265 ;
wire Xd_0__inst_mult_2_266 ;
wire Xd_0__inst_mult_2_268 ;
wire Xd_0__inst_mult_2_269 ;
wire Xd_0__inst_mult_2_270 ;
wire Xd_0__inst_mult_3_308 ;
wire Xd_0__inst_mult_3_309 ;
wire Xd_0__inst_mult_3_310 ;
wire Xd_0__inst_mult_3_312 ;
wire Xd_0__inst_mult_3_313 ;
wire Xd_0__inst_mult_3_314 ;
wire Xd_0__inst_mult_0_284 ;
wire Xd_0__inst_mult_0_285 ;
wire Xd_0__inst_mult_0_286 ;
wire Xd_0__inst_mult_0_288 ;
wire Xd_0__inst_mult_0_289 ;
wire Xd_0__inst_mult_0_290 ;
wire Xd_0__inst_mult_1_268 ;
wire Xd_0__inst_mult_1_269 ;
wire Xd_0__inst_mult_1_270 ;
wire Xd_0__inst_mult_1_272 ;
wire Xd_0__inst_mult_1_273 ;
wire Xd_0__inst_mult_1_274 ;
wire Xd_0__inst_mult_6_397 ;
wire Xd_0__inst_mult_6_398 ;
wire Xd_0__inst_mult_7_405 ;
wire Xd_0__inst_mult_7_406 ;
wire Xd_0__inst_mult_4_272 ;
wire Xd_0__inst_mult_4_273 ;
wire Xd_0__inst_mult_4_274 ;
wire Xd_0__inst_mult_4_276 ;
wire Xd_0__inst_mult_4_277 ;
wire Xd_0__inst_mult_4_278 ;
wire Xd_0__inst_mult_5_35_sumout ;
wire Xd_0__inst_mult_5_36 ;
wire Xd_0__inst_mult_5_37 ;
wire Xd_0__inst_mult_5_272 ;
wire Xd_0__inst_mult_5_273 ;
wire Xd_0__inst_mult_5_274 ;
wire Xd_0__inst_mult_5_276 ;
wire Xd_0__inst_mult_5_277 ;
wire Xd_0__inst_mult_5_278 ;
wire Xd_0__inst_mult_1_47_sumout ;
wire Xd_0__inst_mult_1_48 ;
wire Xd_0__inst_mult_1_49 ;
wire Xd_0__inst_mult_2_272 ;
wire Xd_0__inst_mult_2_273 ;
wire Xd_0__inst_mult_2_274 ;
wire Xd_0__inst_mult_2_276 ;
wire Xd_0__inst_mult_2_277 ;
wire Xd_0__inst_mult_2_278 ;
wire Xd_0__inst_mult_5_39_sumout ;
wire Xd_0__inst_mult_5_40 ;
wire Xd_0__inst_mult_5_41 ;
wire Xd_0__inst_mult_3_316 ;
wire Xd_0__inst_mult_3_317 ;
wire Xd_0__inst_mult_3_318 ;
wire Xd_0__inst_mult_3_320 ;
wire Xd_0__inst_mult_3_321 ;
wire Xd_0__inst_mult_3_322 ;
wire Xd_0__inst_mult_0_39_sumout ;
wire Xd_0__inst_mult_0_40 ;
wire Xd_0__inst_mult_0_41 ;
wire Xd_0__inst_mult_0_292 ;
wire Xd_0__inst_mult_0_293 ;
wire Xd_0__inst_mult_0_294 ;
wire Xd_0__inst_mult_0_296 ;
wire Xd_0__inst_mult_0_297 ;
wire Xd_0__inst_mult_0_298 ;
wire Xd_0__inst_mult_5_43_sumout ;
wire Xd_0__inst_mult_5_44 ;
wire Xd_0__inst_mult_5_45 ;
wire Xd_0__inst_mult_1_276 ;
wire Xd_0__inst_mult_1_277 ;
wire Xd_0__inst_mult_1_278 ;
wire Xd_0__inst_mult_1_280 ;
wire Xd_0__inst_mult_1_281 ;
wire Xd_0__inst_mult_1_282 ;
wire Xd_0__inst_mult_0_43_sumout ;
wire Xd_0__inst_mult_0_44 ;
wire Xd_0__inst_mult_0_45 ;
wire Xd_0__inst_mult_6_400 ;
wire Xd_0__inst_mult_6_401 ;
wire Xd_0__inst_mult_6_402 ;
wire Xd_0__inst_mult_6_404 ;
wire Xd_0__inst_mult_6_405 ;
wire Xd_0__inst_mult_6_406 ;
wire Xd_0__inst_mult_0_47_sumout ;
wire Xd_0__inst_mult_0_48 ;
wire Xd_0__inst_mult_0_49 ;
wire Xd_0__inst_mult_7_408 ;
wire Xd_0__inst_mult_7_409 ;
wire Xd_0__inst_mult_7_410 ;
wire Xd_0__inst_mult_7_412 ;
wire Xd_0__inst_mult_7_413 ;
wire Xd_0__inst_mult_7_414 ;
wire Xd_0__inst_mult_5_47_sumout ;
wire Xd_0__inst_mult_5_48 ;
wire Xd_0__inst_mult_5_49 ;
wire Xd_0__inst_mult_4_280 ;
wire Xd_0__inst_mult_4_281 ;
wire Xd_0__inst_mult_4_282 ;
wire Xd_0__inst_mult_4_284 ;
wire Xd_0__inst_mult_4_285 ;
wire Xd_0__inst_mult_4_286 ;
wire Xd_0__inst_mult_5_280 ;
wire Xd_0__inst_mult_5_281 ;
wire Xd_0__inst_mult_5_282 ;
wire Xd_0__inst_mult_5_284 ;
wire Xd_0__inst_mult_5_285 ;
wire Xd_0__inst_mult_5_286 ;
wire Xd_0__inst_mult_2_280 ;
wire Xd_0__inst_mult_2_281 ;
wire Xd_0__inst_mult_2_282 ;
wire Xd_0__inst_mult_2_284 ;
wire Xd_0__inst_mult_2_285 ;
wire Xd_0__inst_mult_2_286 ;
wire Xd_0__inst_mult_3_324 ;
wire Xd_0__inst_mult_3_325 ;
wire Xd_0__inst_mult_3_326 ;
wire Xd_0__inst_mult_3_328 ;
wire Xd_0__inst_mult_3_329 ;
wire Xd_0__inst_mult_3_330 ;
wire Xd_0__inst_mult_0_300 ;
wire Xd_0__inst_mult_0_301 ;
wire Xd_0__inst_mult_0_302 ;
wire Xd_0__inst_mult_0_304 ;
wire Xd_0__inst_mult_0_305 ;
wire Xd_0__inst_mult_0_306 ;
wire Xd_0__inst_mult_1_284 ;
wire Xd_0__inst_mult_1_285 ;
wire Xd_0__inst_mult_1_286 ;
wire Xd_0__inst_mult_1_288 ;
wire Xd_0__inst_mult_1_289 ;
wire Xd_0__inst_mult_1_290 ;
wire Xd_0__inst_mult_6_408 ;
wire Xd_0__inst_mult_6_409 ;
wire Xd_0__inst_mult_6_410 ;
wire Xd_0__inst_mult_6_412 ;
wire Xd_0__inst_mult_6_413 ;
wire Xd_0__inst_mult_6_414 ;
wire Xd_0__inst_mult_7_416 ;
wire Xd_0__inst_mult_7_417 ;
wire Xd_0__inst_mult_7_418 ;
wire Xd_0__inst_mult_7_420 ;
wire Xd_0__inst_mult_7_421 ;
wire Xd_0__inst_mult_7_422 ;
wire Xd_0__inst_mult_4_288 ;
wire Xd_0__inst_mult_4_289 ;
wire Xd_0__inst_mult_4_290 ;
wire Xd_0__inst_mult_4_292 ;
wire Xd_0__inst_mult_4_293 ;
wire Xd_0__inst_mult_4_294 ;
wire Xd_0__inst_mult_5_288 ;
wire Xd_0__inst_mult_5_289 ;
wire Xd_0__inst_mult_5_290 ;
wire Xd_0__inst_mult_5_292 ;
wire Xd_0__inst_mult_5_293 ;
wire Xd_0__inst_mult_5_294 ;
wire Xd_0__inst_mult_2_288 ;
wire Xd_0__inst_mult_2_289 ;
wire Xd_0__inst_mult_2_290 ;
wire Xd_0__inst_mult_2_292 ;
wire Xd_0__inst_mult_2_293 ;
wire Xd_0__inst_mult_2_294 ;
wire Xd_0__inst_mult_3_332 ;
wire Xd_0__inst_mult_3_333 ;
wire Xd_0__inst_mult_3_334 ;
wire Xd_0__inst_mult_3_336 ;
wire Xd_0__inst_mult_3_337 ;
wire Xd_0__inst_mult_3_338 ;
wire Xd_0__inst_mult_0_308 ;
wire Xd_0__inst_mult_0_309 ;
wire Xd_0__inst_mult_0_310 ;
wire Xd_0__inst_mult_0_312 ;
wire Xd_0__inst_mult_0_313 ;
wire Xd_0__inst_mult_0_314 ;
wire Xd_0__inst_mult_1_292 ;
wire Xd_0__inst_mult_1_293 ;
wire Xd_0__inst_mult_1_294 ;
wire Xd_0__inst_mult_1_296 ;
wire Xd_0__inst_mult_1_297 ;
wire Xd_0__inst_mult_1_298 ;
wire Xd_0__inst_mult_6_416 ;
wire Xd_0__inst_mult_6_417 ;
wire Xd_0__inst_mult_6_418 ;
wire Xd_0__inst_mult_6_420 ;
wire Xd_0__inst_mult_6_421 ;
wire Xd_0__inst_mult_6_422 ;
wire Xd_0__inst_mult_6_55_sumout ;
wire Xd_0__inst_mult_6_56 ;
wire Xd_0__inst_mult_6_57 ;
wire Xd_0__inst_mult_7_424 ;
wire Xd_0__inst_mult_7_425 ;
wire Xd_0__inst_mult_7_426 ;
wire Xd_0__inst_mult_7_428 ;
wire Xd_0__inst_mult_7_429 ;
wire Xd_0__inst_mult_7_430 ;
wire Xd_0__inst_mult_7_55_sumout ;
wire Xd_0__inst_mult_7_56 ;
wire Xd_0__inst_mult_7_57 ;
wire Xd_0__inst_mult_4_296 ;
wire Xd_0__inst_mult_4_297 ;
wire Xd_0__inst_mult_4_298 ;
wire Xd_0__inst_mult_4_300 ;
wire Xd_0__inst_mult_4_301 ;
wire Xd_0__inst_mult_4_302 ;
wire Xd_0__inst_mult_5_296 ;
wire Xd_0__inst_mult_5_297 ;
wire Xd_0__inst_mult_5_298 ;
wire Xd_0__inst_mult_5_300 ;
wire Xd_0__inst_mult_5_301 ;
wire Xd_0__inst_mult_5_302 ;
wire Xd_0__inst_mult_2_296 ;
wire Xd_0__inst_mult_2_297 ;
wire Xd_0__inst_mult_2_298 ;
wire Xd_0__inst_mult_2_300 ;
wire Xd_0__inst_mult_2_301 ;
wire Xd_0__inst_mult_2_302 ;
wire Xd_0__inst_mult_3_340 ;
wire Xd_0__inst_mult_3_341 ;
wire Xd_0__inst_mult_3_342 ;
wire Xd_0__inst_mult_3_344 ;
wire Xd_0__inst_mult_3_345 ;
wire Xd_0__inst_mult_3_346 ;
wire Xd_0__inst_mult_0_316 ;
wire Xd_0__inst_mult_0_317 ;
wire Xd_0__inst_mult_0_318 ;
wire Xd_0__inst_mult_0_320 ;
wire Xd_0__inst_mult_0_321 ;
wire Xd_0__inst_mult_0_322 ;
wire Xd_0__inst_mult_1_300 ;
wire Xd_0__inst_mult_1_301 ;
wire Xd_0__inst_mult_1_302 ;
wire Xd_0__inst_mult_1_304 ;
wire Xd_0__inst_mult_1_305 ;
wire Xd_0__inst_mult_1_306 ;
wire Xd_0__inst_mult_6_424 ;
wire Xd_0__inst_mult_6_425 ;
wire Xd_0__inst_mult_6_426 ;
wire Xd_0__inst_mult_6_428 ;
wire Xd_0__inst_mult_6_429 ;
wire Xd_0__inst_mult_6_430 ;
wire Xd_0__inst_mult_6_59_sumout ;
wire Xd_0__inst_mult_6_60 ;
wire Xd_0__inst_mult_6_61 ;
wire Xd_0__inst_mult_6_432 ;
wire Xd_0__inst_mult_6_433 ;
wire Xd_0__inst_mult_6_434 ;
wire Xd_0__inst_mult_6_437 ;
wire Xd_0__inst_mult_6_438 ;
wire Xd_0__inst_mult_7_432 ;
wire Xd_0__inst_mult_7_433 ;
wire Xd_0__inst_mult_7_434 ;
wire Xd_0__inst_mult_7_436 ;
wire Xd_0__inst_mult_7_437 ;
wire Xd_0__inst_mult_7_438 ;
wire Xd_0__inst_mult_7_59_sumout ;
wire Xd_0__inst_mult_7_60 ;
wire Xd_0__inst_mult_7_61 ;
wire Xd_0__inst_mult_7_440 ;
wire Xd_0__inst_mult_7_441 ;
wire Xd_0__inst_mult_7_442 ;
wire Xd_0__inst_mult_7_445 ;
wire Xd_0__inst_mult_7_446 ;
wire Xd_0__inst_mult_4_304 ;
wire Xd_0__inst_mult_4_305 ;
wire Xd_0__inst_mult_4_306 ;
wire Xd_0__inst_mult_4_308 ;
wire Xd_0__inst_mult_4_309 ;
wire Xd_0__inst_mult_4_310 ;
wire Xd_0__inst_mult_5_304 ;
wire Xd_0__inst_mult_5_305 ;
wire Xd_0__inst_mult_5_306 ;
wire Xd_0__inst_mult_5_308 ;
wire Xd_0__inst_mult_5_309 ;
wire Xd_0__inst_mult_5_310 ;
wire Xd_0__inst_mult_2_304 ;
wire Xd_0__inst_mult_2_305 ;
wire Xd_0__inst_mult_2_306 ;
wire Xd_0__inst_mult_2_308 ;
wire Xd_0__inst_mult_2_309 ;
wire Xd_0__inst_mult_2_310 ;
wire Xd_0__inst_mult_3_348 ;
wire Xd_0__inst_mult_3_349 ;
wire Xd_0__inst_mult_3_350 ;
wire Xd_0__inst_mult_3_352 ;
wire Xd_0__inst_mult_3_353 ;
wire Xd_0__inst_mult_3_354 ;
wire Xd_0__inst_mult_0_324 ;
wire Xd_0__inst_mult_0_325 ;
wire Xd_0__inst_mult_0_326 ;
wire Xd_0__inst_mult_0_328 ;
wire Xd_0__inst_mult_0_329 ;
wire Xd_0__inst_mult_0_330 ;
wire Xd_0__inst_mult_1_308 ;
wire Xd_0__inst_mult_1_309 ;
wire Xd_0__inst_mult_1_310 ;
wire Xd_0__inst_mult_1_312 ;
wire Xd_0__inst_mult_1_313 ;
wire Xd_0__inst_mult_1_314 ;
wire Xd_0__inst_mult_6_440 ;
wire Xd_0__inst_mult_6_441 ;
wire Xd_0__inst_mult_6_442 ;
wire Xd_0__inst_mult_6_444 ;
wire Xd_0__inst_mult_6_445 ;
wire Xd_0__inst_mult_6_446 ;
wire Xd_0__inst_mult_6_63_sumout ;
wire Xd_0__inst_mult_6_64 ;
wire Xd_0__inst_mult_6_65 ;
wire Xd_0__inst_mult_6_448 ;
wire Xd_0__inst_mult_6_449 ;
wire Xd_0__inst_mult_6_450 ;
wire Xd_0__inst_mult_6_452 ;
wire Xd_0__inst_mult_6_453 ;
wire Xd_0__inst_mult_6_454 ;
wire Xd_0__inst_mult_7_448 ;
wire Xd_0__inst_mult_7_449 ;
wire Xd_0__inst_mult_7_450 ;
wire Xd_0__inst_mult_7_452 ;
wire Xd_0__inst_mult_7_453 ;
wire Xd_0__inst_mult_7_454 ;
wire Xd_0__inst_mult_7_63_sumout ;
wire Xd_0__inst_mult_7_64 ;
wire Xd_0__inst_mult_7_65 ;
wire Xd_0__inst_mult_7_456 ;
wire Xd_0__inst_mult_7_457 ;
wire Xd_0__inst_mult_7_458 ;
wire Xd_0__inst_mult_7_460 ;
wire Xd_0__inst_mult_7_461 ;
wire Xd_0__inst_mult_7_462 ;
wire Xd_0__inst_mult_4_312 ;
wire Xd_0__inst_mult_4_313 ;
wire Xd_0__inst_mult_4_314 ;
wire Xd_0__inst_mult_4_316 ;
wire Xd_0__inst_mult_4_317 ;
wire Xd_0__inst_mult_4_318 ;
wire Xd_0__inst_mult_5_312 ;
wire Xd_0__inst_mult_5_313 ;
wire Xd_0__inst_mult_5_314 ;
wire Xd_0__inst_mult_5_316 ;
wire Xd_0__inst_mult_5_317 ;
wire Xd_0__inst_mult_5_318 ;
wire Xd_0__inst_mult_2_312 ;
wire Xd_0__inst_mult_2_313 ;
wire Xd_0__inst_mult_2_314 ;
wire Xd_0__inst_mult_2_316 ;
wire Xd_0__inst_mult_2_317 ;
wire Xd_0__inst_mult_2_318 ;
wire Xd_0__inst_mult_3_356 ;
wire Xd_0__inst_mult_3_357 ;
wire Xd_0__inst_mult_3_358 ;
wire Xd_0__inst_mult_3_360 ;
wire Xd_0__inst_mult_3_361 ;
wire Xd_0__inst_mult_3_362 ;
wire Xd_0__inst_mult_0_332 ;
wire Xd_0__inst_mult_0_333 ;
wire Xd_0__inst_mult_0_334 ;
wire Xd_0__inst_mult_0_336 ;
wire Xd_0__inst_mult_0_337 ;
wire Xd_0__inst_mult_0_338 ;
wire Xd_0__inst_mult_1_316 ;
wire Xd_0__inst_mult_1_317 ;
wire Xd_0__inst_mult_1_318 ;
wire Xd_0__inst_mult_1_320 ;
wire Xd_0__inst_mult_1_321 ;
wire Xd_0__inst_mult_1_322 ;
wire Xd_0__inst_mult_6_456 ;
wire Xd_0__inst_mult_6_457 ;
wire Xd_0__inst_mult_6_458 ;
wire Xd_0__inst_mult_6_460 ;
wire Xd_0__inst_mult_6_461 ;
wire Xd_0__inst_mult_6_462 ;
wire Xd_0__inst_mult_6_67_sumout ;
wire Xd_0__inst_mult_6_68 ;
wire Xd_0__inst_mult_6_69 ;
wire Xd_0__inst_mult_6_464 ;
wire Xd_0__inst_mult_6_465 ;
wire Xd_0__inst_mult_6_466 ;
wire Xd_0__inst_mult_6_468 ;
wire Xd_0__inst_mult_6_469 ;
wire Xd_0__inst_mult_6_470 ;
wire Xd_0__inst_mult_6_472 ;
wire Xd_0__inst_mult_6_473 ;
wire Xd_0__inst_mult_6_474 ;
wire Xd_0__inst_mult_7_464 ;
wire Xd_0__inst_mult_7_465 ;
wire Xd_0__inst_mult_7_466 ;
wire Xd_0__inst_mult_7_468 ;
wire Xd_0__inst_mult_7_469 ;
wire Xd_0__inst_mult_7_470 ;
wire Xd_0__inst_mult_7_67_sumout ;
wire Xd_0__inst_mult_7_68 ;
wire Xd_0__inst_mult_7_69 ;
wire Xd_0__inst_mult_7_472 ;
wire Xd_0__inst_mult_7_473 ;
wire Xd_0__inst_mult_7_474 ;
wire Xd_0__inst_mult_7_476 ;
wire Xd_0__inst_mult_7_477 ;
wire Xd_0__inst_mult_7_478 ;
wire Xd_0__inst_mult_7_480 ;
wire Xd_0__inst_mult_7_481 ;
wire Xd_0__inst_mult_7_482 ;
wire Xd_0__inst_mult_4_320 ;
wire Xd_0__inst_mult_4_321 ;
wire Xd_0__inst_mult_4_322 ;
wire Xd_0__inst_mult_4_324 ;
wire Xd_0__inst_mult_4_325 ;
wire Xd_0__inst_mult_4_326 ;
wire Xd_0__inst_mult_5_320 ;
wire Xd_0__inst_mult_5_321 ;
wire Xd_0__inst_mult_5_322 ;
wire Xd_0__inst_mult_5_324 ;
wire Xd_0__inst_mult_5_325 ;
wire Xd_0__inst_mult_5_326 ;
wire Xd_0__inst_mult_2_320 ;
wire Xd_0__inst_mult_2_321 ;
wire Xd_0__inst_mult_2_322 ;
wire Xd_0__inst_mult_2_324 ;
wire Xd_0__inst_mult_2_325 ;
wire Xd_0__inst_mult_2_326 ;
wire Xd_0__inst_mult_3_364 ;
wire Xd_0__inst_mult_3_365 ;
wire Xd_0__inst_mult_3_366 ;
wire Xd_0__inst_mult_3_368 ;
wire Xd_0__inst_mult_3_369 ;
wire Xd_0__inst_mult_3_370 ;
wire Xd_0__inst_mult_0_340 ;
wire Xd_0__inst_mult_0_341 ;
wire Xd_0__inst_mult_0_342 ;
wire Xd_0__inst_mult_0_344 ;
wire Xd_0__inst_mult_0_345 ;
wire Xd_0__inst_mult_0_346 ;
wire Xd_0__inst_mult_1_324 ;
wire Xd_0__inst_mult_1_325 ;
wire Xd_0__inst_mult_1_326 ;
wire Xd_0__inst_mult_1_328 ;
wire Xd_0__inst_mult_1_329 ;
wire Xd_0__inst_mult_1_330 ;
wire Xd_0__inst_mult_6_476 ;
wire Xd_0__inst_mult_6_477 ;
wire Xd_0__inst_mult_6_478 ;
wire Xd_0__inst_mult_6_480 ;
wire Xd_0__inst_mult_6_481 ;
wire Xd_0__inst_mult_6_482 ;
wire Xd_0__inst_mult_6_484 ;
wire Xd_0__inst_mult_6_485 ;
wire Xd_0__inst_mult_6_486 ;
wire Xd_0__inst_mult_6_488 ;
wire Xd_0__inst_mult_6_489 ;
wire Xd_0__inst_mult_6_490 ;
wire Xd_0__inst_mult_6_492 ;
wire Xd_0__inst_mult_6_493 ;
wire Xd_0__inst_mult_6_494 ;
wire Xd_0__inst_mult_7_484 ;
wire Xd_0__inst_mult_7_485 ;
wire Xd_0__inst_mult_7_486 ;
wire Xd_0__inst_mult_7_488 ;
wire Xd_0__inst_mult_7_489 ;
wire Xd_0__inst_mult_7_490 ;
wire Xd_0__inst_mult_7_492 ;
wire Xd_0__inst_mult_7_493 ;
wire Xd_0__inst_mult_7_494 ;
wire Xd_0__inst_mult_7_496 ;
wire Xd_0__inst_mult_7_497 ;
wire Xd_0__inst_mult_7_498 ;
wire Xd_0__inst_mult_7_500 ;
wire Xd_0__inst_mult_7_501 ;
wire Xd_0__inst_mult_7_502 ;
wire Xd_0__inst_mult_4_328 ;
wire Xd_0__inst_mult_4_329 ;
wire Xd_0__inst_mult_4_330 ;
wire Xd_0__inst_mult_4_332 ;
wire Xd_0__inst_mult_4_333 ;
wire Xd_0__inst_mult_4_334 ;
wire Xd_0__inst_mult_5_328 ;
wire Xd_0__inst_mult_5_329 ;
wire Xd_0__inst_mult_5_330 ;
wire Xd_0__inst_mult_5_332 ;
wire Xd_0__inst_mult_5_333 ;
wire Xd_0__inst_mult_5_334 ;
wire Xd_0__inst_mult_2_328 ;
wire Xd_0__inst_mult_2_329 ;
wire Xd_0__inst_mult_2_330 ;
wire Xd_0__inst_mult_2_332 ;
wire Xd_0__inst_mult_2_333 ;
wire Xd_0__inst_mult_2_334 ;
wire Xd_0__inst_mult_3_372 ;
wire Xd_0__inst_mult_3_373 ;
wire Xd_0__inst_mult_3_374 ;
wire Xd_0__inst_mult_0_348 ;
wire Xd_0__inst_mult_0_349 ;
wire Xd_0__inst_mult_0_350 ;
wire Xd_0__inst_mult_1_332 ;
wire Xd_0__inst_mult_1_333 ;
wire Xd_0__inst_mult_1_334 ;
wire Xd_0__inst_mult_1_336 ;
wire Xd_0__inst_mult_1_337 ;
wire Xd_0__inst_mult_1_338 ;
wire Xd_0__inst_mult_6_496 ;
wire Xd_0__inst_mult_6_500 ;
wire Xd_0__inst_mult_6_501 ;
wire Xd_0__inst_mult_6_502 ;
wire Xd_0__inst_mult_6_504 ;
wire Xd_0__inst_mult_6_505 ;
wire Xd_0__inst_mult_6_506 ;
wire Xd_0__inst_mult_6_508 ;
wire Xd_0__inst_mult_6_509 ;
wire Xd_0__inst_mult_6_510 ;
wire Xd_0__inst_mult_6_512 ;
wire Xd_0__inst_mult_6_513 ;
wire Xd_0__inst_mult_6_514 ;
wire Xd_0__inst_mult_7_504 ;
wire Xd_0__inst_mult_7_505 ;
wire Xd_0__inst_mult_7_506 ;
wire Xd_0__inst_mult_7_508 ;
wire Xd_0__inst_mult_7_509 ;
wire Xd_0__inst_mult_7_510 ;
wire Xd_0__inst_mult_7_512 ;
wire Xd_0__inst_mult_7_513 ;
wire Xd_0__inst_mult_7_514 ;
wire Xd_0__inst_mult_4_336 ;
wire Xd_0__inst_mult_4_337 ;
wire Xd_0__inst_mult_4_338 ;
wire Xd_0__inst_mult_4_340 ;
wire Xd_0__inst_mult_4_341 ;
wire Xd_0__inst_mult_4_342 ;
wire Xd_0__inst_mult_5_336 ;
wire Xd_0__inst_mult_5_337 ;
wire Xd_0__inst_mult_5_338 ;
wire Xd_0__inst_mult_5_340 ;
wire Xd_0__inst_mult_5_341 ;
wire Xd_0__inst_mult_5_342 ;
wire Xd_0__inst_mult_2_336 ;
wire Xd_0__inst_mult_2_337 ;
wire Xd_0__inst_mult_2_338 ;
wire Xd_0__inst_mult_2_340 ;
wire Xd_0__inst_mult_2_341 ;
wire Xd_0__inst_mult_2_342 ;
wire Xd_0__inst_mult_3_376 ;
wire Xd_0__inst_mult_3_377 ;
wire Xd_0__inst_mult_3_378 ;
wire Xd_0__inst_mult_0_352 ;
wire Xd_0__inst_mult_0_353 ;
wire Xd_0__inst_mult_0_354 ;
wire Xd_0__inst_mult_1_340 ;
wire Xd_0__inst_mult_1_341 ;
wire Xd_0__inst_mult_1_342 ;
wire Xd_0__inst_mult_1_344 ;
wire Xd_0__inst_mult_1_345 ;
wire Xd_0__inst_mult_1_346 ;
wire Xd_0__inst_mult_6_516 ;
wire Xd_0__inst_mult_6_517 ;
wire Xd_0__inst_mult_6_518 ;
wire Xd_0__inst_mult_6_520 ;
wire Xd_0__inst_mult_6_521 ;
wire Xd_0__inst_mult_6_522 ;
wire Xd_0__inst_mult_6_524 ;
wire Xd_0__inst_mult_6_525 ;
wire Xd_0__inst_mult_6_526 ;
wire Xd_0__inst_mult_7_516 ;
wire Xd_0__inst_mult_7_517 ;
wire Xd_0__inst_mult_7_518 ;
wire Xd_0__inst_mult_7_520 ;
wire Xd_0__inst_mult_7_521 ;
wire Xd_0__inst_mult_7_522 ;
wire Xd_0__inst_mult_7_524 ;
wire Xd_0__inst_mult_7_525 ;
wire Xd_0__inst_mult_7_526 ;
wire Xd_0__inst_mult_4_344 ;
wire Xd_0__inst_mult_4_345 ;
wire Xd_0__inst_mult_4_346 ;
wire Xd_0__inst_mult_4_348 ;
wire Xd_0__inst_mult_4_349 ;
wire Xd_0__inst_mult_4_350 ;
wire Xd_0__inst_mult_5_344 ;
wire Xd_0__inst_mult_5_345 ;
wire Xd_0__inst_mult_5_346 ;
wire Xd_0__inst_mult_5_348 ;
wire Xd_0__inst_mult_5_349 ;
wire Xd_0__inst_mult_5_350 ;
wire Xd_0__inst_mult_2_344 ;
wire Xd_0__inst_mult_2_345 ;
wire Xd_0__inst_mult_2_346 ;
wire Xd_0__inst_mult_2_348 ;
wire Xd_0__inst_mult_2_349 ;
wire Xd_0__inst_mult_2_350 ;
wire Xd_0__inst_mult_3_380 ;
wire Xd_0__inst_mult_3_381 ;
wire Xd_0__inst_mult_3_382 ;
wire Xd_0__inst_mult_0_356 ;
wire Xd_0__inst_mult_0_357 ;
wire Xd_0__inst_mult_0_358 ;
wire Xd_0__inst_mult_1_348 ;
wire Xd_0__inst_mult_1_349 ;
wire Xd_0__inst_mult_1_350 ;
wire Xd_0__inst_mult_1_352 ;
wire Xd_0__inst_mult_1_353 ;
wire Xd_0__inst_mult_1_354 ;
wire Xd_0__inst_mult_6_528 ;
wire Xd_0__inst_mult_6_529 ;
wire Xd_0__inst_mult_6_530 ;
wire Xd_0__inst_mult_6_532 ;
wire Xd_0__inst_mult_6_533 ;
wire Xd_0__inst_mult_6_534 ;
wire Xd_0__inst_mult_6_536 ;
wire Xd_0__inst_mult_6_537 ;
wire Xd_0__inst_mult_6_538 ;
wire Xd_0__inst_mult_7_528 ;
wire Xd_0__inst_mult_7_529 ;
wire Xd_0__inst_mult_7_530 ;
wire Xd_0__inst_mult_7_532 ;
wire Xd_0__inst_mult_7_533 ;
wire Xd_0__inst_mult_7_534 ;
wire Xd_0__inst_mult_7_536 ;
wire Xd_0__inst_mult_7_537 ;
wire Xd_0__inst_mult_7_538 ;
wire Xd_0__inst_mult_4_352 ;
wire Xd_0__inst_mult_4_356 ;
wire Xd_0__inst_mult_4_357 ;
wire Xd_0__inst_mult_4_358 ;
wire Xd_0__inst_mult_5_352 ;
wire Xd_0__inst_mult_5_356 ;
wire Xd_0__inst_mult_5_357 ;
wire Xd_0__inst_mult_5_358 ;
wire Xd_0__inst_mult_2_352 ;
wire Xd_0__inst_mult_2_356 ;
wire Xd_0__inst_mult_2_357 ;
wire Xd_0__inst_mult_2_358 ;
wire Xd_0__inst_mult_3_384 ;
wire Xd_0__inst_mult_3_385 ;
wire Xd_0__inst_mult_3_386 ;
wire Xd_0__inst_mult_0_360 ;
wire Xd_0__inst_mult_0_361 ;
wire Xd_0__inst_mult_0_362 ;
wire Xd_0__inst_mult_1_356 ;
wire Xd_0__inst_mult_1_360 ;
wire Xd_0__inst_mult_1_361 ;
wire Xd_0__inst_mult_1_362 ;
wire Xd_0__inst_mult_6_540 ;
wire Xd_0__inst_mult_6_541 ;
wire Xd_0__inst_mult_6_542 ;
wire Xd_0__inst_mult_6_544 ;
wire Xd_0__inst_mult_6_545 ;
wire Xd_0__inst_mult_6_546 ;
wire Xd_0__inst_mult_6_548 ;
wire Xd_0__inst_mult_6_549 ;
wire Xd_0__inst_mult_6_550 ;
wire Xd_0__inst_mult_7_540 ;
wire Xd_0__inst_mult_7_541 ;
wire Xd_0__inst_mult_7_542 ;
wire Xd_0__inst_mult_7_544 ;
wire Xd_0__inst_mult_7_545 ;
wire Xd_0__inst_mult_7_546 ;
wire Xd_0__inst_mult_4_360 ;
wire Xd_0__inst_mult_4_361 ;
wire Xd_0__inst_mult_4_362 ;
wire Xd_0__inst_mult_4_364 ;
wire Xd_0__inst_mult_4_365 ;
wire Xd_0__inst_mult_4_366 ;
wire Xd_0__inst_mult_4_39_sumout ;
wire Xd_0__inst_mult_4_40 ;
wire Xd_0__inst_mult_4_41 ;
wire Xd_0__inst_mult_5_360 ;
wire Xd_0__inst_mult_5_361 ;
wire Xd_0__inst_mult_5_362 ;
wire Xd_0__inst_mult_5_51_sumout ;
wire Xd_0__inst_mult_5_52 ;
wire Xd_0__inst_mult_5_53 ;
wire Xd_0__inst_mult_2_360 ;
wire Xd_0__inst_mult_2_361 ;
wire Xd_0__inst_mult_2_362 ;
wire Xd_0__inst_mult_2_51_sumout ;
wire Xd_0__inst_mult_2_52 ;
wire Xd_0__inst_mult_2_53 ;
wire Xd_0__inst_mult_3_388 ;
wire Xd_0__inst_mult_3_389 ;
wire Xd_0__inst_mult_3_390 ;
wire Xd_0__inst_mult_0_364 ;
wire Xd_0__inst_mult_0_365 ;
wire Xd_0__inst_mult_0_366 ;
wire Xd_0__inst_mult_0_51_sumout ;
wire Xd_0__inst_mult_0_52 ;
wire Xd_0__inst_mult_0_53 ;
wire Xd_0__inst_mult_1_364 ;
wire Xd_0__inst_mult_1_365 ;
wire Xd_0__inst_mult_1_366 ;
wire Xd_0__inst_mult_1_51_sumout ;
wire Xd_0__inst_mult_1_52 ;
wire Xd_0__inst_mult_1_53 ;
wire Xd_0__inst_mult_6_552 ;
wire Xd_0__inst_mult_6_553 ;
wire Xd_0__inst_mult_6_554 ;
wire Xd_0__inst_mult_6_556 ;
wire Xd_0__inst_mult_6_557 ;
wire Xd_0__inst_mult_6_558 ;
wire Xd_0__inst_mult_7_548 ;
wire Xd_0__inst_mult_7_549 ;
wire Xd_0__inst_mult_7_550 ;
wire Xd_0__inst_mult_7_552 ;
wire Xd_0__inst_mult_7_553 ;
wire Xd_0__inst_mult_7_554 ;
wire Xd_0__inst_mult_4_368 ;
wire Xd_0__inst_mult_4_369 ;
wire Xd_0__inst_mult_4_370 ;
wire Xd_0__inst_mult_4_43_sumout ;
wire Xd_0__inst_mult_4_44 ;
wire Xd_0__inst_mult_4_45 ;
wire Xd_0__inst_mult_5_364 ;
wire Xd_0__inst_mult_5_365 ;
wire Xd_0__inst_mult_5_366 ;
wire Xd_0__inst_mult_5_55_sumout ;
wire Xd_0__inst_mult_5_56 ;
wire Xd_0__inst_mult_5_57 ;
wire Xd_0__inst_mult_2_364 ;
wire Xd_0__inst_mult_2_365 ;
wire Xd_0__inst_mult_2_366 ;
wire Xd_0__inst_mult_2_55_sumout ;
wire Xd_0__inst_mult_2_56 ;
wire Xd_0__inst_mult_2_57 ;
wire Xd_0__inst_mult_3_392 ;
wire Xd_0__inst_mult_3_393 ;
wire Xd_0__inst_mult_3_394 ;
wire Xd_0__inst_mult_3_43_sumout ;
wire Xd_0__inst_mult_3_44 ;
wire Xd_0__inst_mult_3_45 ;
wire Xd_0__inst_mult_0_368 ;
wire Xd_0__inst_mult_0_369 ;
wire Xd_0__inst_mult_0_370 ;
wire Xd_0__inst_mult_0_55_sumout ;
wire Xd_0__inst_mult_0_56 ;
wire Xd_0__inst_mult_0_57 ;
wire Xd_0__inst_mult_1_368 ;
wire Xd_0__inst_mult_1_369 ;
wire Xd_0__inst_mult_1_370 ;
wire Xd_0__inst_mult_1_55_sumout ;
wire Xd_0__inst_mult_1_56 ;
wire Xd_0__inst_mult_1_57 ;
wire Xd_0__inst_mult_6_560 ;
wire Xd_0__inst_mult_6_564 ;
wire Xd_0__inst_mult_6_565 ;
wire Xd_0__inst_mult_6_566 ;
wire Xd_0__inst_mult_7_556 ;
wire Xd_0__inst_mult_7_560 ;
wire Xd_0__inst_mult_7_561 ;
wire Xd_0__inst_mult_7_562 ;
wire Xd_0__inst_mult_4_372 ;
wire Xd_0__inst_mult_4_373 ;
wire Xd_0__inst_mult_4_374 ;
wire Xd_0__inst_mult_4_47_sumout ;
wire Xd_0__inst_mult_4_48 ;
wire Xd_0__inst_mult_4_49 ;
wire Xd_0__inst_mult_5_368 ;
wire Xd_0__inst_mult_5_369 ;
wire Xd_0__inst_mult_5_370 ;
wire Xd_0__inst_mult_5_59_sumout ;
wire Xd_0__inst_mult_5_60 ;
wire Xd_0__inst_mult_5_61 ;
wire Xd_0__inst_mult_2_368 ;
wire Xd_0__inst_mult_2_369 ;
wire Xd_0__inst_mult_2_370 ;
wire Xd_0__inst_mult_3_396 ;
wire Xd_0__inst_mult_3_397 ;
wire Xd_0__inst_mult_3_398 ;
wire Xd_0__inst_mult_3_47_sumout ;
wire Xd_0__inst_mult_3_48 ;
wire Xd_0__inst_mult_3_49 ;
wire Xd_0__inst_mult_0_372 ;
wire Xd_0__inst_mult_0_373 ;
wire Xd_0__inst_mult_0_374 ;
wire Xd_0__inst_mult_1_372 ;
wire Xd_0__inst_mult_1_373 ;
wire Xd_0__inst_mult_1_374 ;
wire Xd_0__inst_mult_6_568 ;
wire Xd_0__inst_mult_6_569 ;
wire Xd_0__inst_mult_6_570 ;
wire Xd_0__inst_mult_7_564 ;
wire Xd_0__inst_mult_7_565 ;
wire Xd_0__inst_mult_7_566 ;
wire Xd_0__inst_mult_4_376 ;
wire Xd_0__inst_mult_4_377 ;
wire Xd_0__inst_mult_4_378 ;
wire Xd_0__inst_mult_4_51_sumout ;
wire Xd_0__inst_mult_4_52 ;
wire Xd_0__inst_mult_4_53 ;
wire Xd_0__inst_mult_5_372 ;
wire Xd_0__inst_mult_5_373 ;
wire Xd_0__inst_mult_5_374 ;
wire Xd_0__inst_mult_2_372 ;
wire Xd_0__inst_mult_2_373 ;
wire Xd_0__inst_mult_2_374 ;
wire Xd_0__inst_mult_3_400 ;
wire Xd_0__inst_mult_3_401 ;
wire Xd_0__inst_mult_3_402 ;
wire Xd_0__inst_mult_3_51_sumout ;
wire Xd_0__inst_mult_3_52 ;
wire Xd_0__inst_mult_3_53 ;
wire Xd_0__inst_mult_0_376 ;
wire Xd_0__inst_mult_0_377 ;
wire Xd_0__inst_mult_0_378 ;
wire Xd_0__inst_mult_1_376 ;
wire Xd_0__inst_mult_1_377 ;
wire Xd_0__inst_mult_1_378 ;
wire Xd_0__inst_mult_6_572 ;
wire Xd_0__inst_mult_7_568 ;
wire Xd_0__inst_mult_4_380 ;
wire Xd_0__inst_mult_4_55_sumout ;
wire Xd_0__inst_mult_4_56 ;
wire Xd_0__inst_mult_4_57 ;
wire Xd_0__inst_mult_5_376 ;
wire Xd_0__inst_mult_2_376 ;
wire Xd_0__inst_mult_3_404 ;
wire Xd_0__inst_mult_3_55_sumout ;
wire Xd_0__inst_mult_3_56 ;
wire Xd_0__inst_mult_3_57 ;
wire Xd_0__inst_mult_0_380 ;
wire Xd_0__inst_mult_1_380 ;
wire Xd_0__inst_mult_3_408 ;
wire Xd_0__inst_mult_3_409 ;
wire Xd_0__inst_mult_3_410 ;
wire Xd_0__inst_mult_3_412 ;
wire Xd_0__inst_mult_0_384 ;
wire Xd_0__inst_mult_0_385 ;
wire Xd_0__inst_mult_0_386 ;
wire Xd_0__inst_mult_0_388 ;
wire Xd_0__inst_mult_3_416 ;
wire Xd_0__inst_mult_3_417 ;
wire Xd_0__inst_mult_3_418 ;
wire Xd_0__inst_mult_4_384 ;
wire Xd_0__inst_mult_4_385 ;
wire Xd_0__inst_mult_4_386 ;
wire Xd_0__inst_mult_4_388 ;
wire Xd_0__inst_mult_4_389 ;
wire Xd_0__inst_mult_4_390 ;
wire Xd_0__inst_mult_5_380 ;
wire Xd_0__inst_mult_5_381 ;
wire Xd_0__inst_mult_5_382 ;
wire Xd_0__inst_mult_5_384 ;
wire Xd_0__inst_mult_5_385 ;
wire Xd_0__inst_mult_5_386 ;
wire Xd_0__inst_mult_2_380 ;
wire Xd_0__inst_mult_2_381 ;
wire Xd_0__inst_mult_2_382 ;
wire Xd_0__inst_mult_2_384 ;
wire Xd_0__inst_mult_2_385 ;
wire Xd_0__inst_mult_2_386 ;
wire Xd_0__inst_mult_3_420 ;
wire Xd_0__inst_mult_3_421 ;
wire Xd_0__inst_mult_3_422 ;
wire Xd_0__inst_mult_3_425 ;
wire Xd_0__inst_mult_3_426 ;
wire Xd_0__inst_mult_0_392 ;
wire Xd_0__inst_mult_0_393 ;
wire Xd_0__inst_mult_0_394 ;
wire Xd_0__inst_mult_0_397 ;
wire Xd_0__inst_mult_0_398 ;
wire Xd_0__inst_mult_5_63_sumout ;
wire Xd_0__inst_mult_5_64 ;
wire Xd_0__inst_mult_5_65 ;
wire Xd_0__inst_mult_4_393 ;
wire Xd_0__inst_mult_4_394 ;
wire Xd_0__inst_mult_5_389 ;
wire Xd_0__inst_mult_5_390 ;
wire Xd_0__inst_mult_2_389 ;
wire Xd_0__inst_mult_2_390 ;
wire Xd_0__inst_mult_3_429 ;
wire Xd_0__inst_mult_3_430 ;
wire Xd_0__inst_mult_0_401 ;
wire Xd_0__inst_mult_0_402 ;
wire Xd_0__inst_mult_1_385 ;
wire Xd_0__inst_mult_1_386 ;
wire Xd_0__inst_mult_7_572 ;
wire Xd_0__inst_mult_7_573 ;
wire Xd_0__inst_mult_7_574 ;
wire Xd_0__inst_mult_4_396 ;
wire Xd_0__inst_mult_4_397 ;
wire Xd_0__inst_mult_4_398 ;
wire Xd_0__inst_mult_4_400 ;
wire Xd_0__inst_mult_4_401 ;
wire Xd_0__inst_mult_4_402 ;
wire Xd_0__inst_mult_0_59_sumout ;
wire Xd_0__inst_mult_0_60 ;
wire Xd_0__inst_mult_0_61 ;
wire Xd_0__inst_mult_5_392 ;
wire Xd_0__inst_mult_5_393 ;
wire Xd_0__inst_mult_5_394 ;
wire Xd_0__inst_mult_5_396 ;
wire Xd_0__inst_mult_5_397 ;
wire Xd_0__inst_mult_5_398 ;
wire Xd_0__inst_mult_2_392 ;
wire Xd_0__inst_mult_2_393 ;
wire Xd_0__inst_mult_2_394 ;
wire Xd_0__inst_mult_2_396 ;
wire Xd_0__inst_mult_2_397 ;
wire Xd_0__inst_mult_2_398 ;
wire Xd_0__inst_mult_3_432 ;
wire Xd_0__inst_mult_3_433 ;
wire Xd_0__inst_mult_3_434 ;
wire Xd_0__inst_mult_3_436 ;
wire Xd_0__inst_mult_3_437 ;
wire Xd_0__inst_mult_3_438 ;
wire Xd_0__inst_mult_1_59_sumout ;
wire Xd_0__inst_mult_1_60 ;
wire Xd_0__inst_mult_1_61 ;
wire Xd_0__inst_mult_0_404 ;
wire Xd_0__inst_mult_0_405 ;
wire Xd_0__inst_mult_0_406 ;
wire Xd_0__inst_mult_0_408 ;
wire Xd_0__inst_mult_0_409 ;
wire Xd_0__inst_mult_0_410 ;
wire Xd_0__inst_mult_1_388 ;
wire Xd_0__inst_mult_1_389 ;
wire Xd_0__inst_mult_1_390 ;
wire Xd_0__inst_mult_1_392 ;
wire Xd_0__inst_mult_1_393 ;
wire Xd_0__inst_mult_1_394 ;
wire Xd_0__inst_mult_4_404 ;
wire Xd_0__inst_mult_4_405 ;
wire Xd_0__inst_mult_4_406 ;
wire Xd_0__inst_mult_4_408 ;
wire Xd_0__inst_mult_4_409 ;
wire Xd_0__inst_mult_4_410 ;
wire Xd_0__inst_mult_5_400 ;
wire Xd_0__inst_mult_5_401 ;
wire Xd_0__inst_mult_5_402 ;
wire Xd_0__inst_mult_5_404 ;
wire Xd_0__inst_mult_5_405 ;
wire Xd_0__inst_mult_5_406 ;
wire Xd_0__inst_mult_2_400 ;
wire Xd_0__inst_mult_2_401 ;
wire Xd_0__inst_mult_2_402 ;
wire Xd_0__inst_mult_2_404 ;
wire Xd_0__inst_mult_2_405 ;
wire Xd_0__inst_mult_2_406 ;
wire Xd_0__inst_mult_3_440 ;
wire Xd_0__inst_mult_3_441 ;
wire Xd_0__inst_mult_3_442 ;
wire Xd_0__inst_mult_3_444 ;
wire Xd_0__inst_mult_3_445 ;
wire Xd_0__inst_mult_3_446 ;
wire Xd_0__inst_mult_0_412 ;
wire Xd_0__inst_mult_0_413 ;
wire Xd_0__inst_mult_0_414 ;
wire Xd_0__inst_mult_0_416 ;
wire Xd_0__inst_mult_0_417 ;
wire Xd_0__inst_mult_0_418 ;
wire Xd_0__inst_mult_1_396 ;
wire Xd_0__inst_mult_1_397 ;
wire Xd_0__inst_mult_1_398 ;
wire Xd_0__inst_mult_1_400 ;
wire Xd_0__inst_mult_1_401 ;
wire Xd_0__inst_mult_1_402 ;
wire Xd_0__inst_mult_4_412 ;
wire Xd_0__inst_mult_4_413 ;
wire Xd_0__inst_mult_4_414 ;
wire Xd_0__inst_mult_4_416 ;
wire Xd_0__inst_mult_4_417 ;
wire Xd_0__inst_mult_4_418 ;
wire Xd_0__inst_mult_4_59_sumout ;
wire Xd_0__inst_mult_4_60 ;
wire Xd_0__inst_mult_4_61 ;
wire Xd_0__inst_mult_5_408 ;
wire Xd_0__inst_mult_5_409 ;
wire Xd_0__inst_mult_5_410 ;
wire Xd_0__inst_mult_5_412 ;
wire Xd_0__inst_mult_5_413 ;
wire Xd_0__inst_mult_5_414 ;
wire Xd_0__inst_mult_2_408 ;
wire Xd_0__inst_mult_2_409 ;
wire Xd_0__inst_mult_2_410 ;
wire Xd_0__inst_mult_2_412 ;
wire Xd_0__inst_mult_2_413 ;
wire Xd_0__inst_mult_2_414 ;
wire Xd_0__inst_mult_2_59_sumout ;
wire Xd_0__inst_mult_2_60 ;
wire Xd_0__inst_mult_2_61 ;
wire Xd_0__inst_mult_3_448 ;
wire Xd_0__inst_mult_3_449 ;
wire Xd_0__inst_mult_3_450 ;
wire Xd_0__inst_mult_3_452 ;
wire Xd_0__inst_mult_3_453 ;
wire Xd_0__inst_mult_3_454 ;
wire Xd_0__inst_mult_3_59_sumout ;
wire Xd_0__inst_mult_3_60 ;
wire Xd_0__inst_mult_3_61 ;
wire Xd_0__inst_mult_0_420 ;
wire Xd_0__inst_mult_0_421 ;
wire Xd_0__inst_mult_0_422 ;
wire Xd_0__inst_mult_0_424 ;
wire Xd_0__inst_mult_0_425 ;
wire Xd_0__inst_mult_0_426 ;
wire Xd_0__inst_mult_0_63_sumout ;
wire Xd_0__inst_mult_0_64 ;
wire Xd_0__inst_mult_0_65 ;
wire Xd_0__inst_mult_1_404 ;
wire Xd_0__inst_mult_1_405 ;
wire Xd_0__inst_mult_1_406 ;
wire Xd_0__inst_mult_1_408 ;
wire Xd_0__inst_mult_1_409 ;
wire Xd_0__inst_mult_1_410 ;
wire Xd_0__inst_mult_4_420 ;
wire Xd_0__inst_mult_4_421 ;
wire Xd_0__inst_mult_4_422 ;
wire Xd_0__inst_mult_4_424 ;
wire Xd_0__inst_mult_4_425 ;
wire Xd_0__inst_mult_4_426 ;
wire Xd_0__inst_mult_4_63_sumout ;
wire Xd_0__inst_mult_4_64 ;
wire Xd_0__inst_mult_4_65 ;
wire Xd_0__inst_mult_4_428 ;
wire Xd_0__inst_mult_4_429 ;
wire Xd_0__inst_mult_4_430 ;
wire Xd_0__inst_mult_4_433 ;
wire Xd_0__inst_mult_4_434 ;
wire Xd_0__inst_mult_5_416 ;
wire Xd_0__inst_mult_5_417 ;
wire Xd_0__inst_mult_5_418 ;
wire Xd_0__inst_mult_5_420 ;
wire Xd_0__inst_mult_5_421 ;
wire Xd_0__inst_mult_5_422 ;
wire Xd_0__inst_mult_5_67_sumout ;
wire Xd_0__inst_mult_5_68 ;
wire Xd_0__inst_mult_5_69 ;
wire Xd_0__inst_mult_5_424 ;
wire Xd_0__inst_mult_5_425 ;
wire Xd_0__inst_mult_5_426 ;
wire Xd_0__inst_mult_5_429 ;
wire Xd_0__inst_mult_5_430 ;
wire Xd_0__inst_mult_2_416 ;
wire Xd_0__inst_mult_2_417 ;
wire Xd_0__inst_mult_2_418 ;
wire Xd_0__inst_mult_2_420 ;
wire Xd_0__inst_mult_2_421 ;
wire Xd_0__inst_mult_2_422 ;
wire Xd_0__inst_mult_2_63_sumout ;
wire Xd_0__inst_mult_2_64 ;
wire Xd_0__inst_mult_2_65 ;
wire Xd_0__inst_mult_2_424 ;
wire Xd_0__inst_mult_2_425 ;
wire Xd_0__inst_mult_2_426 ;
wire Xd_0__inst_mult_2_429 ;
wire Xd_0__inst_mult_2_430 ;
wire Xd_0__inst_mult_3_456 ;
wire Xd_0__inst_mult_3_457 ;
wire Xd_0__inst_mult_3_458 ;
wire Xd_0__inst_mult_3_460 ;
wire Xd_0__inst_mult_3_461 ;
wire Xd_0__inst_mult_3_462 ;
wire Xd_0__inst_mult_3_63_sumout ;
wire Xd_0__inst_mult_3_64 ;
wire Xd_0__inst_mult_3_65 ;
wire Xd_0__inst_mult_3_464 ;
wire Xd_0__inst_mult_3_465 ;
wire Xd_0__inst_mult_3_466 ;
wire Xd_0__inst_mult_3_469 ;
wire Xd_0__inst_mult_3_470 ;
wire Xd_0__inst_mult_0_428 ;
wire Xd_0__inst_mult_0_429 ;
wire Xd_0__inst_mult_0_430 ;
wire Xd_0__inst_mult_0_432 ;
wire Xd_0__inst_mult_0_433 ;
wire Xd_0__inst_mult_0_434 ;
wire Xd_0__inst_mult_0_436 ;
wire Xd_0__inst_mult_0_437 ;
wire Xd_0__inst_mult_0_438 ;
wire Xd_0__inst_mult_0_441 ;
wire Xd_0__inst_mult_0_442 ;
wire Xd_0__inst_mult_1_412 ;
wire Xd_0__inst_mult_1_413 ;
wire Xd_0__inst_mult_1_414 ;
wire Xd_0__inst_mult_1_416 ;
wire Xd_0__inst_mult_1_417 ;
wire Xd_0__inst_mult_1_418 ;
wire Xd_0__inst_mult_1_63_sumout ;
wire Xd_0__inst_mult_1_64 ;
wire Xd_0__inst_mult_1_65 ;
wire Xd_0__inst_mult_1_420 ;
wire Xd_0__inst_mult_1_421 ;
wire Xd_0__inst_mult_1_422 ;
wire Xd_0__inst_mult_1_425 ;
wire Xd_0__inst_mult_1_426 ;
wire Xd_0__inst_mult_4_436 ;
wire Xd_0__inst_mult_4_437 ;
wire Xd_0__inst_mult_4_438 ;
wire Xd_0__inst_mult_4_440 ;
wire Xd_0__inst_mult_4_441 ;
wire Xd_0__inst_mult_4_442 ;
wire Xd_0__inst_mult_4_67_sumout ;
wire Xd_0__inst_mult_4_68 ;
wire Xd_0__inst_mult_4_69 ;
wire Xd_0__inst_mult_4_444 ;
wire Xd_0__inst_mult_4_445 ;
wire Xd_0__inst_mult_4_446 ;
wire Xd_0__inst_mult_4_448 ;
wire Xd_0__inst_mult_4_449 ;
wire Xd_0__inst_mult_4_450 ;
wire Xd_0__inst_mult_5_432 ;
wire Xd_0__inst_mult_5_433 ;
wire Xd_0__inst_mult_5_434 ;
wire Xd_0__inst_mult_5_436 ;
wire Xd_0__inst_mult_5_437 ;
wire Xd_0__inst_mult_5_438 ;
wire Xd_0__inst_mult_5_440 ;
wire Xd_0__inst_mult_5_441 ;
wire Xd_0__inst_mult_5_442 ;
wire Xd_0__inst_mult_5_444 ;
wire Xd_0__inst_mult_5_445 ;
wire Xd_0__inst_mult_5_446 ;
wire Xd_0__inst_mult_2_432 ;
wire Xd_0__inst_mult_2_433 ;
wire Xd_0__inst_mult_2_434 ;
wire Xd_0__inst_mult_2_436 ;
wire Xd_0__inst_mult_2_437 ;
wire Xd_0__inst_mult_2_438 ;
wire Xd_0__inst_mult_2_67_sumout ;
wire Xd_0__inst_mult_2_68 ;
wire Xd_0__inst_mult_2_69 ;
wire Xd_0__inst_mult_2_440 ;
wire Xd_0__inst_mult_2_441 ;
wire Xd_0__inst_mult_2_442 ;
wire Xd_0__inst_mult_2_444 ;
wire Xd_0__inst_mult_2_445 ;
wire Xd_0__inst_mult_2_446 ;
wire Xd_0__inst_mult_3_472 ;
wire Xd_0__inst_mult_3_473 ;
wire Xd_0__inst_mult_3_474 ;
wire Xd_0__inst_mult_3_476 ;
wire Xd_0__inst_mult_3_477 ;
wire Xd_0__inst_mult_3_478 ;
wire Xd_0__inst_mult_3_480 ;
wire Xd_0__inst_mult_3_481 ;
wire Xd_0__inst_mult_3_482 ;
wire Xd_0__inst_mult_3_484 ;
wire Xd_0__inst_mult_3_485 ;
wire Xd_0__inst_mult_3_486 ;
wire Xd_0__inst_mult_0_444 ;
wire Xd_0__inst_mult_0_445 ;
wire Xd_0__inst_mult_0_446 ;
wire Xd_0__inst_mult_0_448 ;
wire Xd_0__inst_mult_0_449 ;
wire Xd_0__inst_mult_0_450 ;
wire Xd_0__inst_mult_0_452 ;
wire Xd_0__inst_mult_0_453 ;
wire Xd_0__inst_mult_0_454 ;
wire Xd_0__inst_mult_0_456 ;
wire Xd_0__inst_mult_0_457 ;
wire Xd_0__inst_mult_0_458 ;
wire Xd_0__inst_mult_1_428 ;
wire Xd_0__inst_mult_1_429 ;
wire Xd_0__inst_mult_1_430 ;
wire Xd_0__inst_mult_1_432 ;
wire Xd_0__inst_mult_1_433 ;
wire Xd_0__inst_mult_1_434 ;
wire Xd_0__inst_mult_1_436 ;
wire Xd_0__inst_mult_1_437 ;
wire Xd_0__inst_mult_1_438 ;
wire Xd_0__inst_mult_1_440 ;
wire Xd_0__inst_mult_1_441 ;
wire Xd_0__inst_mult_1_442 ;
wire Xd_0__inst_mult_6_577 ;
wire Xd_0__inst_mult_6_578 ;
wire Xd_0__inst_mult_7_577 ;
wire Xd_0__inst_mult_7_578 ;
wire Xd_0__inst_mult_4_452 ;
wire Xd_0__inst_mult_4_453 ;
wire Xd_0__inst_mult_4_454 ;
wire Xd_0__inst_mult_4_456 ;
wire Xd_0__inst_mult_4_457 ;
wire Xd_0__inst_mult_4_458 ;
wire Xd_0__inst_mult_4_460 ;
wire Xd_0__inst_mult_4_461 ;
wire Xd_0__inst_mult_4_462 ;
wire Xd_0__inst_mult_4_464 ;
wire Xd_0__inst_mult_4_465 ;
wire Xd_0__inst_mult_4_466 ;
wire Xd_0__inst_mult_4_468 ;
wire Xd_0__inst_mult_4_469 ;
wire Xd_0__inst_mult_4_470 ;
wire Xd_0__inst_mult_5_448 ;
wire Xd_0__inst_mult_5_449 ;
wire Xd_0__inst_mult_5_450 ;
wire Xd_0__inst_mult_5_452 ;
wire Xd_0__inst_mult_5_453 ;
wire Xd_0__inst_mult_5_454 ;
wire Xd_0__inst_mult_5_456 ;
wire Xd_0__inst_mult_5_457 ;
wire Xd_0__inst_mult_5_458 ;
wire Xd_0__inst_mult_5_460 ;
wire Xd_0__inst_mult_5_461 ;
wire Xd_0__inst_mult_5_462 ;
wire Xd_0__inst_mult_5_464 ;
wire Xd_0__inst_mult_5_465 ;
wire Xd_0__inst_mult_5_466 ;
wire Xd_0__inst_mult_2_448 ;
wire Xd_0__inst_mult_2_449 ;
wire Xd_0__inst_mult_2_450 ;
wire Xd_0__inst_mult_2_452 ;
wire Xd_0__inst_mult_2_453 ;
wire Xd_0__inst_mult_2_454 ;
wire Xd_0__inst_mult_2_456 ;
wire Xd_0__inst_mult_2_457 ;
wire Xd_0__inst_mult_2_458 ;
wire Xd_0__inst_mult_2_460 ;
wire Xd_0__inst_mult_2_461 ;
wire Xd_0__inst_mult_2_462 ;
wire Xd_0__inst_mult_2_464 ;
wire Xd_0__inst_mult_2_465 ;
wire Xd_0__inst_mult_2_466 ;
wire Xd_0__inst_mult_3_488 ;
wire Xd_0__inst_mult_3_489 ;
wire Xd_0__inst_mult_3_490 ;
wire Xd_0__inst_mult_3_492 ;
wire Xd_0__inst_mult_3_493 ;
wire Xd_0__inst_mult_3_494 ;
wire Xd_0__inst_mult_3_496 ;
wire Xd_0__inst_mult_3_497 ;
wire Xd_0__inst_mult_3_498 ;
wire Xd_0__inst_mult_3_500 ;
wire Xd_0__inst_mult_3_501 ;
wire Xd_0__inst_mult_3_502 ;
wire Xd_0__inst_mult_3_504 ;
wire Xd_0__inst_mult_3_505 ;
wire Xd_0__inst_mult_3_506 ;
wire Xd_0__inst_mult_0_460 ;
wire Xd_0__inst_mult_0_461 ;
wire Xd_0__inst_mult_0_462 ;
wire Xd_0__inst_mult_0_464 ;
wire Xd_0__inst_mult_0_465 ;
wire Xd_0__inst_mult_0_466 ;
wire Xd_0__inst_mult_0_468 ;
wire Xd_0__inst_mult_0_469 ;
wire Xd_0__inst_mult_0_470 ;
wire Xd_0__inst_mult_0_472 ;
wire Xd_0__inst_mult_0_473 ;
wire Xd_0__inst_mult_0_474 ;
wire Xd_0__inst_mult_0_476 ;
wire Xd_0__inst_mult_0_477 ;
wire Xd_0__inst_mult_0_478 ;
wire Xd_0__inst_mult_1_444 ;
wire Xd_0__inst_mult_1_445 ;
wire Xd_0__inst_mult_1_446 ;
wire Xd_0__inst_mult_1_448 ;
wire Xd_0__inst_mult_1_449 ;
wire Xd_0__inst_mult_1_450 ;
wire Xd_0__inst_mult_1_452 ;
wire Xd_0__inst_mult_1_453 ;
wire Xd_0__inst_mult_1_454 ;
wire Xd_0__inst_mult_1_456 ;
wire Xd_0__inst_mult_1_457 ;
wire Xd_0__inst_mult_1_458 ;
wire Xd_0__inst_mult_1_460 ;
wire Xd_0__inst_mult_1_461 ;
wire Xd_0__inst_mult_1_462 ;
wire Xd_0__inst_mult_6_581 ;
wire Xd_0__inst_mult_6_582 ;
wire Xd_0__inst_mult_7_581 ;
wire Xd_0__inst_mult_7_582 ;
wire Xd_0__inst_mult_4_472 ;
wire Xd_0__inst_mult_4_473 ;
wire Xd_0__inst_mult_4_474 ;
wire Xd_0__inst_mult_4_476 ;
wire Xd_0__inst_mult_4_477 ;
wire Xd_0__inst_mult_4_478 ;
wire Xd_0__inst_mult_4_480 ;
wire Xd_0__inst_mult_4_481 ;
wire Xd_0__inst_mult_4_482 ;
wire Xd_0__inst_mult_4_484 ;
wire Xd_0__inst_mult_4_485 ;
wire Xd_0__inst_mult_4_486 ;
wire Xd_0__inst_mult_4_488 ;
wire Xd_0__inst_mult_4_489 ;
wire Xd_0__inst_mult_4_490 ;
wire Xd_0__inst_mult_5_468 ;
wire Xd_0__inst_mult_5_469 ;
wire Xd_0__inst_mult_5_470 ;
wire Xd_0__inst_mult_5_472 ;
wire Xd_0__inst_mult_5_473 ;
wire Xd_0__inst_mult_5_474 ;
wire Xd_0__inst_mult_5_476 ;
wire Xd_0__inst_mult_5_477 ;
wire Xd_0__inst_mult_5_478 ;
wire Xd_0__inst_mult_5_480 ;
wire Xd_0__inst_mult_5_481 ;
wire Xd_0__inst_mult_5_482 ;
wire Xd_0__inst_mult_5_484 ;
wire Xd_0__inst_mult_5_485 ;
wire Xd_0__inst_mult_5_486 ;
wire Xd_0__inst_mult_2_468 ;
wire Xd_0__inst_mult_2_469 ;
wire Xd_0__inst_mult_2_470 ;
wire Xd_0__inst_mult_2_472 ;
wire Xd_0__inst_mult_2_473 ;
wire Xd_0__inst_mult_2_474 ;
wire Xd_0__inst_mult_2_476 ;
wire Xd_0__inst_mult_2_477 ;
wire Xd_0__inst_mult_2_478 ;
wire Xd_0__inst_mult_2_480 ;
wire Xd_0__inst_mult_2_481 ;
wire Xd_0__inst_mult_2_482 ;
wire Xd_0__inst_mult_2_484 ;
wire Xd_0__inst_mult_2_485 ;
wire Xd_0__inst_mult_2_486 ;
wire Xd_0__inst_mult_3_508 ;
wire Xd_0__inst_mult_3_509 ;
wire Xd_0__inst_mult_3_510 ;
wire Xd_0__inst_mult_3_512 ;
wire Xd_0__inst_mult_3_513 ;
wire Xd_0__inst_mult_3_514 ;
wire Xd_0__inst_mult_3_516 ;
wire Xd_0__inst_mult_3_517 ;
wire Xd_0__inst_mult_3_518 ;
wire Xd_0__inst_mult_3_520 ;
wire Xd_0__inst_mult_3_521 ;
wire Xd_0__inst_mult_3_522 ;
wire Xd_0__inst_mult_3_524 ;
wire Xd_0__inst_mult_3_525 ;
wire Xd_0__inst_mult_3_526 ;
wire Xd_0__inst_mult_0_480 ;
wire Xd_0__inst_mult_0_481 ;
wire Xd_0__inst_mult_0_482 ;
wire Xd_0__inst_mult_0_484 ;
wire Xd_0__inst_mult_0_485 ;
wire Xd_0__inst_mult_0_486 ;
wire Xd_0__inst_mult_0_488 ;
wire Xd_0__inst_mult_0_489 ;
wire Xd_0__inst_mult_0_490 ;
wire Xd_0__inst_mult_0_492 ;
wire Xd_0__inst_mult_0_493 ;
wire Xd_0__inst_mult_0_494 ;
wire Xd_0__inst_mult_0_496 ;
wire Xd_0__inst_mult_0_497 ;
wire Xd_0__inst_mult_0_498 ;
wire Xd_0__inst_mult_1_464 ;
wire Xd_0__inst_mult_1_465 ;
wire Xd_0__inst_mult_1_466 ;
wire Xd_0__inst_mult_1_468 ;
wire Xd_0__inst_mult_1_469 ;
wire Xd_0__inst_mult_1_470 ;
wire Xd_0__inst_mult_1_472 ;
wire Xd_0__inst_mult_1_473 ;
wire Xd_0__inst_mult_1_474 ;
wire Xd_0__inst_mult_1_476 ;
wire Xd_0__inst_mult_1_477 ;
wire Xd_0__inst_mult_1_478 ;
wire Xd_0__inst_mult_1_480 ;
wire Xd_0__inst_mult_1_481 ;
wire Xd_0__inst_mult_1_482 ;
wire Xd_0__inst_mult_4_492 ;
wire Xd_0__inst_mult_4_496 ;
wire Xd_0__inst_mult_4_497 ;
wire Xd_0__inst_mult_4_498 ;
wire Xd_0__inst_mult_4_500 ;
wire Xd_0__inst_mult_4_501 ;
wire Xd_0__inst_mult_4_502 ;
wire Xd_0__inst_mult_4_504 ;
wire Xd_0__inst_mult_4_505 ;
wire Xd_0__inst_mult_4_506 ;
wire Xd_0__inst_mult_4_508 ;
wire Xd_0__inst_mult_4_509 ;
wire Xd_0__inst_mult_4_510 ;
wire Xd_0__inst_mult_5_488 ;
wire Xd_0__inst_mult_5_492 ;
wire Xd_0__inst_mult_5_493 ;
wire Xd_0__inst_mult_5_494 ;
wire Xd_0__inst_mult_5_496 ;
wire Xd_0__inst_mult_5_497 ;
wire Xd_0__inst_mult_5_498 ;
wire Xd_0__inst_mult_5_500 ;
wire Xd_0__inst_mult_5_501 ;
wire Xd_0__inst_mult_5_502 ;
wire Xd_0__inst_mult_5_504 ;
wire Xd_0__inst_mult_5_505 ;
wire Xd_0__inst_mult_5_506 ;
wire Xd_0__inst_mult_2_488 ;
wire Xd_0__inst_mult_2_492 ;
wire Xd_0__inst_mult_2_493 ;
wire Xd_0__inst_mult_2_494 ;
wire Xd_0__inst_mult_2_496 ;
wire Xd_0__inst_mult_2_497 ;
wire Xd_0__inst_mult_2_498 ;
wire Xd_0__inst_mult_2_500 ;
wire Xd_0__inst_mult_2_501 ;
wire Xd_0__inst_mult_2_502 ;
wire Xd_0__inst_mult_2_504 ;
wire Xd_0__inst_mult_2_505 ;
wire Xd_0__inst_mult_2_506 ;
wire Xd_0__inst_mult_3_528 ;
wire Xd_0__inst_mult_3_529 ;
wire Xd_0__inst_mult_3_530 ;
wire Xd_0__inst_mult_3_532 ;
wire Xd_0__inst_mult_3_533 ;
wire Xd_0__inst_mult_3_534 ;
wire Xd_0__inst_mult_3_536 ;
wire Xd_0__inst_mult_3_537 ;
wire Xd_0__inst_mult_3_538 ;
wire Xd_0__inst_mult_0_500 ;
wire Xd_0__inst_mult_0_501 ;
wire Xd_0__inst_mult_0_502 ;
wire Xd_0__inst_mult_0_504 ;
wire Xd_0__inst_mult_0_505 ;
wire Xd_0__inst_mult_0_506 ;
wire Xd_0__inst_mult_0_508 ;
wire Xd_0__inst_mult_0_509 ;
wire Xd_0__inst_mult_0_510 ;
wire Xd_0__inst_mult_1_484 ;
wire Xd_0__inst_mult_1_488 ;
wire Xd_0__inst_mult_1_489 ;
wire Xd_0__inst_mult_1_490 ;
wire Xd_0__inst_mult_1_492 ;
wire Xd_0__inst_mult_1_493 ;
wire Xd_0__inst_mult_1_494 ;
wire Xd_0__inst_mult_1_496 ;
wire Xd_0__inst_mult_1_497 ;
wire Xd_0__inst_mult_1_498 ;
wire Xd_0__inst_mult_1_500 ;
wire Xd_0__inst_mult_1_501 ;
wire Xd_0__inst_mult_1_502 ;
wire Xd_0__inst_mult_4_512 ;
wire Xd_0__inst_mult_4_513 ;
wire Xd_0__inst_mult_4_514 ;
wire Xd_0__inst_mult_4_516 ;
wire Xd_0__inst_mult_4_517 ;
wire Xd_0__inst_mult_4_518 ;
wire Xd_0__inst_mult_4_520 ;
wire Xd_0__inst_mult_4_521 ;
wire Xd_0__inst_mult_4_522 ;
wire Xd_0__inst_mult_4_524 ;
wire Xd_0__inst_mult_4_525 ;
wire Xd_0__inst_mult_4_526 ;
wire Xd_0__inst_mult_5_508 ;
wire Xd_0__inst_mult_5_509 ;
wire Xd_0__inst_mult_5_510 ;
wire Xd_0__inst_mult_5_512 ;
wire Xd_0__inst_mult_5_513 ;
wire Xd_0__inst_mult_5_514 ;
wire Xd_0__inst_mult_5_516 ;
wire Xd_0__inst_mult_5_517 ;
wire Xd_0__inst_mult_5_518 ;
wire Xd_0__inst_mult_5_520 ;
wire Xd_0__inst_mult_5_521 ;
wire Xd_0__inst_mult_5_522 ;
wire Xd_0__inst_mult_2_508 ;
wire Xd_0__inst_mult_2_509 ;
wire Xd_0__inst_mult_2_510 ;
wire Xd_0__inst_mult_2_512 ;
wire Xd_0__inst_mult_2_513 ;
wire Xd_0__inst_mult_2_514 ;
wire Xd_0__inst_mult_2_516 ;
wire Xd_0__inst_mult_2_517 ;
wire Xd_0__inst_mult_2_518 ;
wire Xd_0__inst_mult_2_520 ;
wire Xd_0__inst_mult_2_521 ;
wire Xd_0__inst_mult_2_522 ;
wire Xd_0__inst_mult_3_540 ;
wire Xd_0__inst_mult_3_541 ;
wire Xd_0__inst_mult_3_542 ;
wire Xd_0__inst_mult_3_544 ;
wire Xd_0__inst_mult_3_545 ;
wire Xd_0__inst_mult_3_546 ;
wire Xd_0__inst_mult_0_512 ;
wire Xd_0__inst_mult_0_513 ;
wire Xd_0__inst_mult_0_514 ;
wire Xd_0__inst_mult_0_516 ;
wire Xd_0__inst_mult_0_517 ;
wire Xd_0__inst_mult_0_518 ;
wire Xd_0__inst_mult_0_520 ;
wire Xd_0__inst_mult_0_521 ;
wire Xd_0__inst_mult_0_522 ;
wire Xd_0__inst_mult_1_504 ;
wire Xd_0__inst_mult_1_505 ;
wire Xd_0__inst_mult_1_506 ;
wire Xd_0__inst_mult_1_508 ;
wire Xd_0__inst_mult_1_509 ;
wire Xd_0__inst_mult_1_510 ;
wire Xd_0__inst_mult_1_512 ;
wire Xd_0__inst_mult_1_513 ;
wire Xd_0__inst_mult_1_514 ;
wire Xd_0__inst_mult_1_516 ;
wire Xd_0__inst_mult_1_517 ;
wire Xd_0__inst_mult_1_518 ;
wire Xd_0__inst_mult_4_528 ;
wire Xd_0__inst_mult_4_532 ;
wire Xd_0__inst_mult_4_533 ;
wire Xd_0__inst_mult_4_534 ;
wire Xd_0__inst_mult_4_536 ;
wire Xd_0__inst_mult_4_537 ;
wire Xd_0__inst_mult_4_538 ;
wire Xd_0__inst_mult_4_540 ;
wire Xd_0__inst_mult_4_541 ;
wire Xd_0__inst_mult_4_542 ;
wire Xd_0__inst_mult_5_524 ;
wire Xd_0__inst_mult_5_528 ;
wire Xd_0__inst_mult_5_529 ;
wire Xd_0__inst_mult_5_530 ;
wire Xd_0__inst_mult_5_532 ;
wire Xd_0__inst_mult_5_533 ;
wire Xd_0__inst_mult_5_534 ;
wire Xd_0__inst_mult_5_536 ;
wire Xd_0__inst_mult_5_537 ;
wire Xd_0__inst_mult_5_538 ;
wire Xd_0__inst_mult_2_524 ;
wire Xd_0__inst_mult_2_528 ;
wire Xd_0__inst_mult_2_529 ;
wire Xd_0__inst_mult_2_530 ;
wire Xd_0__inst_mult_2_532 ;
wire Xd_0__inst_mult_2_533 ;
wire Xd_0__inst_mult_2_534 ;
wire Xd_0__inst_mult_2_536 ;
wire Xd_0__inst_mult_2_537 ;
wire Xd_0__inst_mult_2_538 ;
wire Xd_0__inst_mult_3_548 ;
wire Xd_0__inst_mult_3_549 ;
wire Xd_0__inst_mult_3_550 ;
wire Xd_0__inst_mult_3_552 ;
wire Xd_0__inst_mult_3_553 ;
wire Xd_0__inst_mult_3_554 ;
wire Xd_0__inst_mult_0_524 ;
wire Xd_0__inst_mult_0_525 ;
wire Xd_0__inst_mult_0_526 ;
wire Xd_0__inst_mult_0_528 ;
wire Xd_0__inst_mult_0_529 ;
wire Xd_0__inst_mult_0_530 ;
wire Xd_0__inst_mult_0_532 ;
wire Xd_0__inst_mult_0_533 ;
wire Xd_0__inst_mult_0_534 ;
wire Xd_0__inst_mult_1_520 ;
wire Xd_0__inst_mult_1_524 ;
wire Xd_0__inst_mult_1_525 ;
wire Xd_0__inst_mult_1_526 ;
wire Xd_0__inst_mult_1_528 ;
wire Xd_0__inst_mult_1_529 ;
wire Xd_0__inst_mult_1_530 ;
wire Xd_0__inst_mult_1_532 ;
wire Xd_0__inst_mult_1_533 ;
wire Xd_0__inst_mult_1_534 ;
wire Xd_0__inst_mult_4_544 ;
wire Xd_0__inst_mult_4_545 ;
wire Xd_0__inst_mult_4_546 ;
wire Xd_0__inst_mult_4_548 ;
wire Xd_0__inst_mult_4_549 ;
wire Xd_0__inst_mult_4_550 ;
wire Xd_0__inst_mult_5_540 ;
wire Xd_0__inst_mult_5_541 ;
wire Xd_0__inst_mult_5_542 ;
wire Xd_0__inst_mult_5_544 ;
wire Xd_0__inst_mult_5_545 ;
wire Xd_0__inst_mult_5_546 ;
wire Xd_0__inst_mult_5_548 ;
wire Xd_0__inst_mult_5_549 ;
wire Xd_0__inst_mult_5_550 ;
wire Xd_0__inst_mult_2_540 ;
wire Xd_0__inst_mult_2_541 ;
wire Xd_0__inst_mult_2_542 ;
wire Xd_0__inst_mult_2_544 ;
wire Xd_0__inst_mult_2_545 ;
wire Xd_0__inst_mult_2_546 ;
wire Xd_0__inst_mult_1_536 ;
wire Xd_0__inst_mult_1_537 ;
wire Xd_0__inst_mult_1_538 ;
wire Xd_0__inst_mult_3_556 ;
wire Xd_0__inst_mult_3_557 ;
wire Xd_0__inst_mult_3_558 ;
wire Xd_0__inst_mult_2_548 ;
wire Xd_0__inst_mult_2_549 ;
wire Xd_0__inst_mult_2_550 ;
wire Xd_0__inst_mult_0_536 ;
wire Xd_0__inst_mult_0_537 ;
wire Xd_0__inst_mult_0_538 ;
wire Xd_0__inst_mult_0_540 ;
wire Xd_0__inst_mult_0_541 ;
wire Xd_0__inst_mult_0_542 ;
wire Xd_0__inst_mult_0_544 ;
wire Xd_0__inst_mult_0_545 ;
wire Xd_0__inst_mult_0_546 ;
wire Xd_0__inst_mult_1_540 ;
wire Xd_0__inst_mult_1_541 ;
wire Xd_0__inst_mult_1_542 ;
wire Xd_0__inst_mult_1_544 ;
wire Xd_0__inst_mult_1_545 ;
wire Xd_0__inst_mult_1_546 ;
wire Xd_0__inst_mult_1_548 ;
wire Xd_0__inst_mult_1_549 ;
wire Xd_0__inst_mult_1_550 ;
wire Xd_0__inst_mult_4_552 ;
wire Xd_0__inst_mult_4_553 ;
wire Xd_0__inst_mult_4_554 ;
wire Xd_0__inst_mult_4_556 ;
wire Xd_0__inst_mult_4_557 ;
wire Xd_0__inst_mult_4_558 ;
wire Xd_0__inst_mult_5_552 ;
wire Xd_0__inst_mult_5_553 ;
wire Xd_0__inst_mult_5_554 ;
wire Xd_0__inst_mult_5_556 ;
wire Xd_0__inst_mult_5_557 ;
wire Xd_0__inst_mult_5_558 ;
wire Xd_0__inst_mult_2_552 ;
wire Xd_0__inst_mult_2_553 ;
wire Xd_0__inst_mult_2_554 ;
wire Xd_0__inst_mult_2_556 ;
wire Xd_0__inst_mult_2_557 ;
wire Xd_0__inst_mult_2_558 ;
wire Xd_0__inst_mult_3_560 ;
wire Xd_0__inst_mult_3_561 ;
wire Xd_0__inst_mult_3_562 ;
wire Xd_0__inst_mult_0_548 ;
wire Xd_0__inst_mult_0_549 ;
wire Xd_0__inst_mult_0_550 ;
wire Xd_0__inst_mult_0_552 ;
wire Xd_0__inst_mult_0_553 ;
wire Xd_0__inst_mult_0_554 ;
wire Xd_0__inst_mult_1_552 ;
wire Xd_0__inst_mult_1_553 ;
wire Xd_0__inst_mult_1_554 ;
wire Xd_0__inst_mult_1_556 ;
wire Xd_0__inst_mult_1_557 ;
wire Xd_0__inst_mult_1_558 ;
wire Xd_0__inst_mult_4_560 ;
wire Xd_0__inst_mult_4_564 ;
wire Xd_0__inst_mult_4_565 ;
wire Xd_0__inst_mult_4_566 ;
wire Xd_0__inst_mult_5_560 ;
wire Xd_0__inst_mult_5_564 ;
wire Xd_0__inst_mult_5_565 ;
wire Xd_0__inst_mult_5_566 ;
wire Xd_0__inst_mult_2_560 ;
wire Xd_0__inst_mult_2_564 ;
wire Xd_0__inst_mult_2_565 ;
wire Xd_0__inst_mult_2_566 ;
wire Xd_0__inst_mult_3_564 ;
wire Xd_0__inst_mult_0_556 ;
wire Xd_0__inst_mult_0_560 ;
wire Xd_0__inst_mult_0_561 ;
wire Xd_0__inst_mult_0_562 ;
wire Xd_0__inst_mult_1_560 ;
wire Xd_0__inst_mult_1_564 ;
wire Xd_0__inst_mult_1_565 ;
wire Xd_0__inst_mult_1_566 ;
wire Xd_0__inst_mult_4_568 ;
wire Xd_0__inst_mult_4_569 ;
wire Xd_0__inst_mult_4_570 ;
wire Xd_0__inst_mult_5_568 ;
wire Xd_0__inst_mult_5_569 ;
wire Xd_0__inst_mult_5_570 ;
wire Xd_0__inst_mult_2_568 ;
wire Xd_0__inst_mult_2_569 ;
wire Xd_0__inst_mult_2_570 ;
wire Xd_0__inst_mult_0_564 ;
wire Xd_0__inst_mult_0_565 ;
wire Xd_0__inst_mult_0_566 ;
wire Xd_0__inst_mult_1_568 ;
wire Xd_0__inst_mult_1_569 ;
wire Xd_0__inst_mult_1_570 ;
wire Xd_0__inst_mult_4_572 ;
wire Xd_0__inst_mult_5_572 ;
wire Xd_0__inst_mult_2_572 ;
wire Xd_0__inst_mult_0_568 ;
wire Xd_0__inst_mult_1_572 ;
wire Xd_0__inst_mult_4_577 ;
wire Xd_0__inst_mult_4_578 ;
wire Xd_0__inst_mult_5_577 ;
wire Xd_0__inst_mult_5_578 ;
wire Xd_0__inst_mult_2_577 ;
wire Xd_0__inst_mult_2_578 ;
wire Xd_0__inst_mult_3_569 ;
wire Xd_0__inst_mult_3_570 ;
wire Xd_0__inst_mult_0_573 ;
wire Xd_0__inst_mult_0_574 ;
wire Xd_0__inst_mult_4_581 ;
wire Xd_0__inst_mult_4_582 ;
wire Xd_0__inst_mult_5_581 ;
wire Xd_0__inst_mult_5_582 ;
wire Xd_0__inst_mult_2_581 ;
wire Xd_0__inst_mult_2_582 ;
wire Xd_0__inst_mult_3_573 ;
wire Xd_0__inst_mult_3_574 ;
wire Xd_0__inst_mult_0_577 ;
wire Xd_0__inst_mult_0_578 ;
wire Xd_0__inst_mult_1_577 ;
wire Xd_0__inst_mult_1_578 ;
wire Xd_0__inst_mult_6_585 ;
wire Xd_0__inst_mult_6_586 ;
wire Xd_0__inst_mult_7_585 ;
wire Xd_0__inst_mult_7_586 ;
wire Xd_0__inst_mult_4_585 ;
wire Xd_0__inst_mult_4_586 ;
wire Xd_0__inst_mult_5_585 ;
wire Xd_0__inst_mult_5_586 ;
wire Xd_0__inst_mult_2_585 ;
wire Xd_0__inst_mult_2_586 ;
wire Xd_0__inst_mult_3_577 ;
wire Xd_0__inst_mult_3_578 ;
wire Xd_0__inst_mult_0_581 ;
wire Xd_0__inst_mult_0_582 ;
wire Xd_0__inst_mult_1_581 ;
wire Xd_0__inst_mult_1_582 ;
wire Xd_0__inst_mult_3_581 ;
wire Xd_0__inst_mult_3_582 ;
wire Xd_0__inst_inst_first_level_0__0__q ;
wire Xd_0__inst_inst_first_level_1__0__q ;
wire Xd_0__inst_inst_first_level_0__1__q ;
wire Xd_0__inst_inst_first_level_1__1__q ;
wire Xd_0__inst_inst_first_level_0__2__q ;
wire Xd_0__inst_inst_first_level_1__2__q ;
wire Xd_0__inst_inst_first_level_0__3__q ;
wire Xd_0__inst_inst_first_level_1__3__q ;
wire Xd_0__inst_inst_first_level_0__4__q ;
wire Xd_0__inst_inst_first_level_1__4__q ;
wire Xd_0__inst_inst_first_level_0__5__q ;
wire Xd_0__inst_inst_first_level_1__5__q ;
wire Xd_0__inst_inst_first_level_0__6__q ;
wire Xd_0__inst_inst_first_level_1__6__q ;
wire Xd_0__inst_inst_first_level_0__7__q ;
wire Xd_0__inst_inst_first_level_1__7__q ;
wire Xd_0__inst_inst_first_level_0__8__q ;
wire Xd_0__inst_inst_first_level_1__8__q ;
wire Xd_0__inst_inst_first_level_0__9__q ;
wire Xd_0__inst_inst_first_level_1__9__q ;
wire Xd_0__inst_inst_first_level_0__10__q ;
wire Xd_0__inst_inst_first_level_1__10__q ;
wire Xd_0__inst_inst_first_level_0__11__q ;
wire Xd_0__inst_inst_first_level_1__11__q ;
wire Xd_0__inst_inst_first_level_0__12__q ;
wire Xd_0__inst_inst_first_level_1__12__q ;
wire Xd_0__inst_inst_first_level_0__13__q ;
wire Xd_0__inst_inst_first_level_1__13__q ;
wire Xd_0__inst_inst_first_level_0__14__q ;
wire Xd_0__inst_inst_first_level_1__14__q ;
wire Xd_0__inst_inst_first_level_0__15__q ;
wire Xd_0__inst_inst_first_level_1__15__q ;
wire Xd_0__inst_inst_first_level_0__16__q ;
wire Xd_0__inst_inst_first_level_1__16__q ;
wire Xd_0__inst_inst_first_level_0__17__q ;
wire Xd_0__inst_inst_first_level_1__17__q ;
wire Xd_0__inst_inst_first_level_0__18__q ;
wire Xd_0__inst_inst_first_level_1__18__q ;
wire Xd_0__inst_inst_first_level_0__19__q ;
wire Xd_0__inst_inst_first_level_1__19__q ;
wire Xd_0__inst_inst_first_level_0__20__q ;
wire Xd_0__inst_inst_first_level_1__20__q ;
wire Xd_0__inst_inst_first_level_0__21__q ;
wire Xd_0__inst_inst_first_level_1__21__q ;
wire Xd_0__inst_inst_first_level_0__22__q ;
wire Xd_0__inst_inst_first_level_1__22__q ;
wire Xd_0__inst_inst_first_level_0__23__q ;
wire Xd_0__inst_inst_first_level_1__25__q ;
wire Xd_0__inst_inst_first_level_0__24__q ;
wire Xd_0__inst_inst_first_level_0__25__q ;
wire Xd_0__inst_r_sum1_3__0__q ;
wire Xd_0__inst_r_sum1_3__1__q ;
wire Xd_0__inst_r_sum1_3__2__q ;
wire Xd_0__inst_r_sum1_3__3__q ;
wire Xd_0__inst_r_sum1_3__4__q ;
wire Xd_0__inst_r_sum1_3__5__q ;
wire Xd_0__inst_r_sum1_3__6__q ;
wire Xd_0__inst_r_sum1_3__7__q ;
wire Xd_0__inst_r_sum1_3__8__q ;
wire Xd_0__inst_r_sum1_3__9__q ;
wire Xd_0__inst_r_sum1_3__10__q ;
wire Xd_0__inst_r_sum1_3__11__q ;
wire Xd_0__inst_r_sum1_3__12__q ;
wire Xd_0__inst_r_sum1_3__13__q ;
wire Xd_0__inst_r_sum1_3__14__q ;
wire Xd_0__inst_r_sum1_3__15__q ;
wire Xd_0__inst_r_sum1_3__16__q ;
wire Xd_0__inst_r_sum1_3__17__q ;
wire Xd_0__inst_r_sum1_3__18__q ;
wire Xd_0__inst_r_sum1_3__19__q ;
wire Xd_0__inst_r_sum1_3__20__q ;
wire Xd_0__inst_r_sum1_3__21__q ;
wire Xd_0__inst_r_sum1_3__22__q ;
wire Xd_0__inst_r_sum1_3__23__q ;
wire Xd_0__inst_r_sum1_2__0__q ;
wire Xd_0__inst_r_sum1_1__0__q ;
wire Xd_0__inst_r_sum1_0__0__q ;
wire Xd_0__inst_r_sum1_2__1__q ;
wire Xd_0__inst_r_sum1_1__1__q ;
wire Xd_0__inst_r_sum1_0__1__q ;
wire Xd_0__inst_r_sum1_2__2__q ;
wire Xd_0__inst_r_sum1_1__2__q ;
wire Xd_0__inst_r_sum1_0__2__q ;
wire Xd_0__inst_r_sum1_2__3__q ;
wire Xd_0__inst_r_sum1_1__3__q ;
wire Xd_0__inst_r_sum1_0__3__q ;
wire Xd_0__inst_r_sum1_2__4__q ;
wire Xd_0__inst_r_sum1_1__4__q ;
wire Xd_0__inst_r_sum1_0__4__q ;
wire Xd_0__inst_r_sum1_2__5__q ;
wire Xd_0__inst_r_sum1_1__5__q ;
wire Xd_0__inst_r_sum1_0__5__q ;
wire Xd_0__inst_r_sum1_2__6__q ;
wire Xd_0__inst_r_sum1_1__6__q ;
wire Xd_0__inst_r_sum1_0__6__q ;
wire Xd_0__inst_r_sum1_2__7__q ;
wire Xd_0__inst_r_sum1_1__7__q ;
wire Xd_0__inst_r_sum1_0__7__q ;
wire Xd_0__inst_r_sum1_2__8__q ;
wire Xd_0__inst_r_sum1_1__8__q ;
wire Xd_0__inst_r_sum1_0__8__q ;
wire Xd_0__inst_r_sum1_2__9__q ;
wire Xd_0__inst_r_sum1_1__9__q ;
wire Xd_0__inst_r_sum1_0__9__q ;
wire Xd_0__inst_r_sum1_2__10__q ;
wire Xd_0__inst_r_sum1_1__10__q ;
wire Xd_0__inst_r_sum1_0__10__q ;
wire Xd_0__inst_r_sum1_2__11__q ;
wire Xd_0__inst_r_sum1_1__11__q ;
wire Xd_0__inst_r_sum1_0__11__q ;
wire Xd_0__inst_r_sum1_2__12__q ;
wire Xd_0__inst_r_sum1_1__12__q ;
wire Xd_0__inst_r_sum1_0__12__q ;
wire Xd_0__inst_r_sum1_2__13__q ;
wire Xd_0__inst_r_sum1_1__13__q ;
wire Xd_0__inst_r_sum1_0__13__q ;
wire Xd_0__inst_r_sum1_2__14__q ;
wire Xd_0__inst_r_sum1_1__14__q ;
wire Xd_0__inst_r_sum1_0__14__q ;
wire Xd_0__inst_r_sum1_2__15__q ;
wire Xd_0__inst_r_sum1_1__15__q ;
wire Xd_0__inst_r_sum1_0__15__q ;
wire Xd_0__inst_r_sum1_2__16__q ;
wire Xd_0__inst_r_sum1_1__16__q ;
wire Xd_0__inst_r_sum1_0__16__q ;
wire Xd_0__inst_r_sum1_2__17__q ;
wire Xd_0__inst_r_sum1_1__17__q ;
wire Xd_0__inst_r_sum1_0__17__q ;
wire Xd_0__inst_r_sum1_2__18__q ;
wire Xd_0__inst_r_sum1_1__18__q ;
wire Xd_0__inst_r_sum1_0__18__q ;
wire Xd_0__inst_r_sum1_2__19__q ;
wire Xd_0__inst_r_sum1_1__19__q ;
wire Xd_0__inst_r_sum1_0__19__q ;
wire Xd_0__inst_r_sum1_2__20__q ;
wire Xd_0__inst_r_sum1_1__20__q ;
wire Xd_0__inst_r_sum1_0__20__q ;
wire Xd_0__inst_r_sum1_2__21__q ;
wire Xd_0__inst_r_sum1_1__21__q ;
wire Xd_0__inst_r_sum1_0__21__q ;
wire Xd_0__inst_r_sum1_2__22__q ;
wire Xd_0__inst_r_sum1_1__22__q ;
wire Xd_0__inst_r_sum1_0__22__q ;
wire Xd_0__inst_r_sum1_2__23__q ;
wire Xd_0__inst_r_sum1_1__23__q ;
wire Xd_0__inst_r_sum1_0__23__q ;
wire Xd_0__inst_product_6__0__q ;
wire Xd_0__inst_product_7__0__q ;
wire Xd_0__inst_product_6__1__q ;
wire Xd_0__inst_product_7__1__q ;
wire Xd_0__inst_product_6__2__q ;
wire Xd_0__inst_product_7__2__q ;
wire Xd_0__inst_product_6__3__q ;
wire Xd_0__inst_product_7__3__q ;
wire Xd_0__inst_product_6__4__q ;
wire Xd_0__inst_product_7__4__q ;
wire Xd_0__inst_product_6__5__q ;
wire Xd_0__inst_product_7__5__q ;
wire Xd_0__inst_product_6__6__q ;
wire Xd_0__inst_product_7__6__q ;
wire Xd_0__inst_product_6__7__q ;
wire Xd_0__inst_product_7__7__q ;
wire Xd_0__inst_product_6__8__q ;
wire Xd_0__inst_product_7__8__q ;
wire Xd_0__inst_product_6__9__q ;
wire Xd_0__inst_product_7__9__q ;
wire Xd_0__inst_product_6__10__q ;
wire Xd_0__inst_product_7__10__q ;
wire Xd_0__inst_product_6__11__q ;
wire Xd_0__inst_product_7__11__q ;
wire Xd_0__inst_product_6__12__q ;
wire Xd_0__inst_product_7__12__q ;
wire Xd_0__inst_product_6__13__q ;
wire Xd_0__inst_product_7__13__q ;
wire Xd_0__inst_product_6__14__q ;
wire Xd_0__inst_product_7__14__q ;
wire Xd_0__inst_product_6__15__q ;
wire Xd_0__inst_product_7__15__q ;
wire Xd_0__inst_product_6__16__q ;
wire Xd_0__inst_product_7__16__q ;
wire Xd_0__inst_product_6__17__q ;
wire Xd_0__inst_product_7__17__q ;
wire Xd_0__inst_product_6__18__q ;
wire Xd_0__inst_product_7__18__q ;
wire Xd_0__inst_product_6__19__q ;
wire Xd_0__inst_product_7__19__q ;
wire Xd_0__inst_product_6__20__q ;
wire Xd_0__inst_product_7__20__q ;
wire Xd_0__inst_product_6__21__q ;
wire Xd_0__inst_product_7__21__q ;
wire Xd_0__inst_product_4__0__q ;
wire Xd_0__inst_product_5__0__q ;
wire Xd_0__inst_product_2__0__q ;
wire Xd_0__inst_product_3__0__q ;
wire Xd_0__inst_product_0__0__q ;
wire Xd_0__inst_product_1__0__q ;
wire Xd_0__inst_product1_6__0__q ;
wire Xd_0__inst_product1_7__0__q ;
wire Xd_0__inst_product_4__1__q ;
wire Xd_0__inst_product_5__1__q ;
wire Xd_0__inst_product_2__1__q ;
wire Xd_0__inst_product_3__1__q ;
wire Xd_0__inst_product_0__1__q ;
wire Xd_0__inst_product_1__1__q ;
wire Xd_0__inst_product1_6__1__q ;
wire Xd_0__inst_product1_7__1__q ;
wire Xd_0__inst_product_4__2__q ;
wire Xd_0__inst_product_5__2__q ;
wire Xd_0__inst_product_2__2__q ;
wire Xd_0__inst_product_3__2__q ;
wire Xd_0__inst_product_0__2__q ;
wire Xd_0__inst_product_1__2__q ;
wire Xd_0__inst_product1_6__2__q ;
wire Xd_0__inst_product1_7__2__q ;
wire Xd_0__inst_product_4__3__q ;
wire Xd_0__inst_product_5__3__q ;
wire Xd_0__inst_product_2__3__q ;
wire Xd_0__inst_product_3__3__q ;
wire Xd_0__inst_product_0__3__q ;
wire Xd_0__inst_product_1__3__q ;
wire Xd_0__inst_product1_6__3__q ;
wire Xd_0__inst_product1_7__3__q ;
wire Xd_0__inst_product_4__4__q ;
wire Xd_0__inst_product_5__4__q ;
wire Xd_0__inst_product_2__4__q ;
wire Xd_0__inst_product_3__4__q ;
wire Xd_0__inst_product_0__4__q ;
wire Xd_0__inst_product_1__4__q ;
wire Xd_0__inst_product1_6__4__q ;
wire Xd_0__inst_product1_7__4__q ;
wire Xd_0__inst_product_4__5__q ;
wire Xd_0__inst_product_5__5__q ;
wire Xd_0__inst_product_2__5__q ;
wire Xd_0__inst_product_3__5__q ;
wire Xd_0__inst_product_0__5__q ;
wire Xd_0__inst_product_1__5__q ;
wire Xd_0__inst_product_4__6__q ;
wire Xd_0__inst_product_5__6__q ;
wire Xd_0__inst_product_2__6__q ;
wire Xd_0__inst_product_3__6__q ;
wire Xd_0__inst_product_0__6__q ;
wire Xd_0__inst_product_1__6__q ;
wire Xd_0__inst_product_4__7__q ;
wire Xd_0__inst_product_5__7__q ;
wire Xd_0__inst_product_2__7__q ;
wire Xd_0__inst_product_3__7__q ;
wire Xd_0__inst_product_0__7__q ;
wire Xd_0__inst_product_1__7__q ;
wire Xd_0__inst_product_4__8__q ;
wire Xd_0__inst_product_5__8__q ;
wire Xd_0__inst_product_2__8__q ;
wire Xd_0__inst_product_3__8__q ;
wire Xd_0__inst_product_0__8__q ;
wire Xd_0__inst_product_1__8__q ;
wire Xd_0__inst_product_4__9__q ;
wire Xd_0__inst_product_5__9__q ;
wire Xd_0__inst_product_2__9__q ;
wire Xd_0__inst_product_3__9__q ;
wire Xd_0__inst_product_0__9__q ;
wire Xd_0__inst_product_1__9__q ;
wire Xd_0__inst_product_4__10__q ;
wire Xd_0__inst_product_5__10__q ;
wire Xd_0__inst_product_2__10__q ;
wire Xd_0__inst_product_3__10__q ;
wire Xd_0__inst_product_0__10__q ;
wire Xd_0__inst_product_1__10__q ;
wire Xd_0__inst_product_4__11__q ;
wire Xd_0__inst_product_5__11__q ;
wire Xd_0__inst_product_2__11__q ;
wire Xd_0__inst_product_3__11__q ;
wire Xd_0__inst_product_0__11__q ;
wire Xd_0__inst_product_1__11__q ;
wire Xd_0__inst_product_4__12__q ;
wire Xd_0__inst_product_5__12__q ;
wire Xd_0__inst_product_2__12__q ;
wire Xd_0__inst_product_3__12__q ;
wire Xd_0__inst_product_0__12__q ;
wire Xd_0__inst_product_1__12__q ;
wire Xd_0__inst_product_4__13__q ;
wire Xd_0__inst_product_5__13__q ;
wire Xd_0__inst_product_2__13__q ;
wire Xd_0__inst_product_3__13__q ;
wire Xd_0__inst_product_0__13__q ;
wire Xd_0__inst_product_1__13__q ;
wire Xd_0__inst_product_4__14__q ;
wire Xd_0__inst_product_5__14__q ;
wire Xd_0__inst_product_2__14__q ;
wire Xd_0__inst_product_3__14__q ;
wire Xd_0__inst_product_0__14__q ;
wire Xd_0__inst_product_1__14__q ;
wire Xd_0__inst_product_4__15__q ;
wire Xd_0__inst_product_5__15__q ;
wire Xd_0__inst_product_2__15__q ;
wire Xd_0__inst_product_3__15__q ;
wire Xd_0__inst_product_0__15__q ;
wire Xd_0__inst_product_1__15__q ;
wire Xd_0__inst_product_4__16__q ;
wire Xd_0__inst_product_5__16__q ;
wire Xd_0__inst_product_2__16__q ;
wire Xd_0__inst_product_3__16__q ;
wire Xd_0__inst_product_0__16__q ;
wire Xd_0__inst_product_1__16__q ;
wire Xd_0__inst_product_4__17__q ;
wire Xd_0__inst_product_5__17__q ;
wire Xd_0__inst_product_2__17__q ;
wire Xd_0__inst_product_3__17__q ;
wire Xd_0__inst_product_0__17__q ;
wire Xd_0__inst_product_1__17__q ;
wire Xd_0__inst_product_4__18__q ;
wire Xd_0__inst_product_5__18__q ;
wire Xd_0__inst_product_2__18__q ;
wire Xd_0__inst_product_3__18__q ;
wire Xd_0__inst_product_0__18__q ;
wire Xd_0__inst_product_1__18__q ;
wire Xd_0__inst_product_4__19__q ;
wire Xd_0__inst_product_5__19__q ;
wire Xd_0__inst_product_2__19__q ;
wire Xd_0__inst_product_3__19__q ;
wire Xd_0__inst_product_0__19__q ;
wire Xd_0__inst_product_1__19__q ;
wire Xd_0__inst_product_4__20__q ;
wire Xd_0__inst_product_5__20__q ;
wire Xd_0__inst_product_2__20__q ;
wire Xd_0__inst_product_3__20__q ;
wire Xd_0__inst_product_0__20__q ;
wire Xd_0__inst_product_1__20__q ;
wire Xd_0__inst_product_4__21__q ;
wire Xd_0__inst_product_5__21__q ;
wire Xd_0__inst_product_2__21__q ;
wire Xd_0__inst_product_3__21__q ;
wire Xd_0__inst_product_0__21__q ;
wire Xd_0__inst_product_1__21__q ;
wire Xd_0__inst_product1_4__0__q ;
wire Xd_0__inst_product1_5__0__q ;
wire Xd_0__inst_product1_2__0__q ;
wire Xd_0__inst_product1_3__0__q ;
wire Xd_0__inst_product1_0__0__q ;
wire Xd_0__inst_product1_1__0__q ;
wire Xd_0__inst_product1_4__1__q ;
wire Xd_0__inst_product1_5__1__q ;
wire Xd_0__inst_product1_2__1__q ;
wire Xd_0__inst_product1_3__1__q ;
wire Xd_0__inst_product1_0__1__q ;
wire Xd_0__inst_product1_1__1__q ;
wire Xd_0__inst_product1_4__2__q ;
wire Xd_0__inst_product1_5__2__q ;
wire Xd_0__inst_product1_2__2__q ;
wire Xd_0__inst_product1_3__2__q ;
wire Xd_0__inst_product1_0__2__q ;
wire Xd_0__inst_product1_1__2__q ;
wire Xd_0__inst_product1_4__3__q ;
wire Xd_0__inst_product1_5__3__q ;
wire Xd_0__inst_product1_2__3__q ;
wire Xd_0__inst_product1_3__3__q ;
wire Xd_0__inst_product1_0__3__q ;
wire Xd_0__inst_product1_1__3__q ;
wire Xd_0__inst_product1_4__4__q ;
wire Xd_0__inst_product1_5__4__q ;
wire Xd_0__inst_product1_2__4__q ;
wire Xd_0__inst_product1_3__4__q ;
wire Xd_0__inst_product1_0__4__q ;
wire Xd_0__inst_product1_1__4__q ;
wire Xd_0__inst_mult_6_0_q ;
wire Xd_0__inst_mult_6_1_q ;
wire Xd_0__inst_mult_7_0_q ;
wire Xd_0__inst_mult_7_1_q ;
wire Xd_0__inst_mult_6_2_q ;
wire Xd_0__inst_mult_6_3_q ;
wire Xd_0__inst_mult_7_2_q ;
wire Xd_0__inst_mult_7_3_q ;
wire Xd_0__inst_mult_6_4_q ;
wire Xd_0__inst_mult_6_5_q ;
wire Xd_0__inst_mult_7_4_q ;
wire Xd_0__inst_mult_7_5_q ;
wire Xd_0__inst_mult_6_6_q ;
wire Xd_0__inst_mult_6_7_q ;
wire Xd_0__inst_mult_7_6_q ;
wire Xd_0__inst_mult_7_7_q ;
wire Xd_0__inst_mult_6_8_q ;
wire Xd_0__inst_mult_6_9_q ;
wire Xd_0__inst_mult_7_8_q ;
wire Xd_0__inst_mult_7_9_q ;
wire Xd_0__inst_mult_6_10_q ;
wire Xd_0__inst_mult_6_11_q ;
wire Xd_0__inst_mult_7_10_q ;
wire Xd_0__inst_mult_7_11_q ;
wire Xd_0__inst_mult_6_12_q ;
wire Xd_0__inst_mult_6_13_q ;
wire Xd_0__inst_mult_7_12_q ;
wire Xd_0__inst_mult_7_13_q ;
wire Xd_0__inst_mult_6_14_q ;
wire Xd_0__inst_mult_6_15_q ;
wire Xd_0__inst_mult_7_14_q ;
wire Xd_0__inst_mult_7_15_q ;
wire Xd_0__inst_mult_6_16_q ;
wire Xd_0__inst_mult_6_17_q ;
wire Xd_0__inst_mult_7_16_q ;
wire Xd_0__inst_mult_7_17_q ;
wire Xd_0__inst_mult_6_18_q ;
wire Xd_0__inst_mult_6_19_q ;
wire Xd_0__inst_mult_7_18_q ;
wire Xd_0__inst_mult_7_19_q ;
wire Xd_0__inst_mult_6_20_q ;
wire Xd_0__inst_mult_6_21_q ;
wire Xd_0__inst_mult_6_22_q ;
wire Xd_0__inst_mult_6_23_q ;
wire Xd_0__inst_mult_7_20_q ;
wire Xd_0__inst_mult_7_21_q ;
wire Xd_0__inst_mult_7_22_q ;
wire Xd_0__inst_mult_7_23_q ;
wire Xd_0__inst_mult_6_24_q ;
wire Xd_0__inst_mult_6_25_q ;
wire Xd_0__inst_mult_7_24_q ;
wire Xd_0__inst_mult_7_25_q ;
wire Xd_0__inst_mult_6_26_q ;
wire Xd_0__inst_mult_6_27_q ;
wire Xd_0__inst_mult_7_26_q ;
wire Xd_0__inst_mult_7_27_q ;
wire Xd_0__inst_mult_6_28_q ;
wire Xd_0__inst_mult_6_29_q ;
wire Xd_0__inst_mult_7_28_q ;
wire Xd_0__inst_mult_7_29_q ;
wire Xd_0__inst_mult_6_30_q ;
wire Xd_0__inst_mult_6_31_q ;
wire Xd_0__inst_mult_7_30_q ;
wire Xd_0__inst_mult_7_31_q ;
wire Xd_0__inst_mult_6_32_q ;
wire Xd_0__inst_mult_6_33_q ;
wire Xd_0__inst_mult_7_32_q ;
wire Xd_0__inst_mult_7_33_q ;
wire Xd_0__inst_mult_4_0_q ;
wire Xd_0__inst_mult_4_1_q ;
wire Xd_0__inst_mult_5_0_q ;
wire Xd_0__inst_mult_5_1_q ;
wire Xd_0__inst_mult_2_0_q ;
wire Xd_0__inst_mult_2_1_q ;
wire Xd_0__inst_mult_3_0_q ;
wire Xd_0__inst_mult_3_1_q ;
wire Xd_0__inst_mult_0_0_q ;
wire Xd_0__inst_mult_0_1_q ;
wire Xd_0__inst_mult_1_0_q ;
wire Xd_0__inst_mult_1_1_q ;
wire Xd_0__inst_mult_4_2_q ;
wire Xd_0__inst_mult_4_3_q ;
wire Xd_0__inst_mult_5_2_q ;
wire Xd_0__inst_mult_5_3_q ;
wire Xd_0__inst_mult_2_2_q ;
wire Xd_0__inst_mult_2_3_q ;
wire Xd_0__inst_mult_3_2_q ;
wire Xd_0__inst_mult_3_3_q ;
wire Xd_0__inst_mult_0_2_q ;
wire Xd_0__inst_mult_0_3_q ;
wire Xd_0__inst_mult_1_2_q ;
wire Xd_0__inst_mult_1_3_q ;
wire Xd_0__inst_mult_4_4_q ;
wire Xd_0__inst_mult_4_5_q ;
wire Xd_0__inst_mult_5_4_q ;
wire Xd_0__inst_mult_5_5_q ;
wire Xd_0__inst_mult_2_4_q ;
wire Xd_0__inst_mult_2_5_q ;
wire Xd_0__inst_mult_3_4_q ;
wire Xd_0__inst_mult_3_5_q ;
wire Xd_0__inst_mult_0_4_q ;
wire Xd_0__inst_mult_0_5_q ;
wire Xd_0__inst_mult_1_4_q ;
wire Xd_0__inst_mult_1_5_q ;
wire Xd_0__inst_mult_4_6_q ;
wire Xd_0__inst_mult_4_7_q ;
wire Xd_0__inst_mult_5_6_q ;
wire Xd_0__inst_mult_5_7_q ;
wire Xd_0__inst_mult_2_6_q ;
wire Xd_0__inst_mult_2_7_q ;
wire Xd_0__inst_mult_3_6_q ;
wire Xd_0__inst_mult_3_7_q ;
wire Xd_0__inst_mult_0_6_q ;
wire Xd_0__inst_mult_0_7_q ;
wire Xd_0__inst_mult_1_6_q ;
wire Xd_0__inst_mult_1_7_q ;
wire Xd_0__inst_mult_4_8_q ;
wire Xd_0__inst_mult_4_9_q ;
wire Xd_0__inst_mult_5_8_q ;
wire Xd_0__inst_mult_5_9_q ;
wire Xd_0__inst_mult_2_8_q ;
wire Xd_0__inst_mult_2_9_q ;
wire Xd_0__inst_mult_3_8_q ;
wire Xd_0__inst_mult_3_9_q ;
wire Xd_0__inst_mult_0_8_q ;
wire Xd_0__inst_mult_0_9_q ;
wire Xd_0__inst_mult_1_8_q ;
wire Xd_0__inst_mult_1_9_q ;
wire Xd_0__inst_mult_4_10_q ;
wire Xd_0__inst_mult_4_11_q ;
wire Xd_0__inst_mult_5_10_q ;
wire Xd_0__inst_mult_5_11_q ;
wire Xd_0__inst_mult_2_10_q ;
wire Xd_0__inst_mult_2_11_q ;
wire Xd_0__inst_mult_3_10_q ;
wire Xd_0__inst_mult_3_11_q ;
wire Xd_0__inst_mult_0_10_q ;
wire Xd_0__inst_mult_0_11_q ;
wire Xd_0__inst_mult_1_10_q ;
wire Xd_0__inst_mult_1_11_q ;
wire Xd_0__inst_mult_4_12_q ;
wire Xd_0__inst_mult_4_13_q ;
wire Xd_0__inst_mult_5_12_q ;
wire Xd_0__inst_mult_5_13_q ;
wire Xd_0__inst_mult_2_12_q ;
wire Xd_0__inst_mult_2_13_q ;
wire Xd_0__inst_mult_3_12_q ;
wire Xd_0__inst_mult_3_13_q ;
wire Xd_0__inst_mult_0_12_q ;
wire Xd_0__inst_mult_0_13_q ;
wire Xd_0__inst_mult_1_12_q ;
wire Xd_0__inst_mult_1_13_q ;
wire Xd_0__inst_mult_4_14_q ;
wire Xd_0__inst_mult_4_15_q ;
wire Xd_0__inst_mult_5_14_q ;
wire Xd_0__inst_mult_5_15_q ;
wire Xd_0__inst_mult_2_14_q ;
wire Xd_0__inst_mult_2_15_q ;
wire Xd_0__inst_mult_3_14_q ;
wire Xd_0__inst_mult_3_15_q ;
wire Xd_0__inst_mult_0_14_q ;
wire Xd_0__inst_mult_0_15_q ;
wire Xd_0__inst_mult_1_14_q ;
wire Xd_0__inst_mult_1_15_q ;
wire Xd_0__inst_mult_4_16_q ;
wire Xd_0__inst_mult_4_17_q ;
wire Xd_0__inst_mult_5_16_q ;
wire Xd_0__inst_mult_5_17_q ;
wire Xd_0__inst_mult_2_16_q ;
wire Xd_0__inst_mult_2_17_q ;
wire Xd_0__inst_mult_3_16_q ;
wire Xd_0__inst_mult_3_17_q ;
wire Xd_0__inst_mult_0_16_q ;
wire Xd_0__inst_mult_0_17_q ;
wire Xd_0__inst_mult_1_16_q ;
wire Xd_0__inst_mult_1_17_q ;
wire Xd_0__inst_mult_4_18_q ;
wire Xd_0__inst_mult_4_19_q ;
wire Xd_0__inst_mult_5_18_q ;
wire Xd_0__inst_mult_5_19_q ;
wire Xd_0__inst_mult_2_18_q ;
wire Xd_0__inst_mult_2_19_q ;
wire Xd_0__inst_mult_3_18_q ;
wire Xd_0__inst_mult_3_19_q ;
wire Xd_0__inst_mult_0_18_q ;
wire Xd_0__inst_mult_0_19_q ;
wire Xd_0__inst_mult_1_18_q ;
wire Xd_0__inst_mult_1_19_q ;
wire Xd_0__inst_mult_4_20_q ;
wire Xd_0__inst_mult_4_21_q ;
wire Xd_0__inst_mult_4_22_q ;
wire Xd_0__inst_mult_4_23_q ;
wire Xd_0__inst_mult_5_20_q ;
wire Xd_0__inst_mult_5_21_q ;
wire Xd_0__inst_mult_5_22_q ;
wire Xd_0__inst_mult_5_23_q ;
wire Xd_0__inst_mult_2_20_q ;
wire Xd_0__inst_mult_2_21_q ;
wire Xd_0__inst_mult_2_22_q ;
wire Xd_0__inst_mult_2_23_q ;
wire Xd_0__inst_mult_3_20_q ;
wire Xd_0__inst_mult_3_21_q ;
wire Xd_0__inst_mult_3_22_q ;
wire Xd_0__inst_mult_3_23_q ;
wire Xd_0__inst_mult_0_20_q ;
wire Xd_0__inst_mult_0_21_q ;
wire Xd_0__inst_mult_0_22_q ;
wire Xd_0__inst_mult_0_23_q ;
wire Xd_0__inst_mult_1_20_q ;
wire Xd_0__inst_mult_1_21_q ;
wire Xd_0__inst_mult_1_22_q ;
wire Xd_0__inst_mult_1_23_q ;
wire Xd_0__inst_mult_4_24_q ;
wire Xd_0__inst_mult_4_25_q ;
wire Xd_0__inst_mult_5_24_q ;
wire Xd_0__inst_mult_5_25_q ;
wire Xd_0__inst_mult_2_24_q ;
wire Xd_0__inst_mult_2_25_q ;
wire Xd_0__inst_mult_3_24_q ;
wire Xd_0__inst_mult_3_25_q ;
wire Xd_0__inst_mult_0_24_q ;
wire Xd_0__inst_mult_0_25_q ;
wire Xd_0__inst_mult_1_24_q ;
wire Xd_0__inst_mult_1_25_q ;
wire Xd_0__inst_mult_4_26_q ;
wire Xd_0__inst_mult_4_27_q ;
wire Xd_0__inst_mult_5_26_q ;
wire Xd_0__inst_mult_5_27_q ;
wire Xd_0__inst_mult_2_26_q ;
wire Xd_0__inst_mult_2_27_q ;
wire Xd_0__inst_mult_3_26_q ;
wire Xd_0__inst_mult_3_27_q ;
wire Xd_0__inst_mult_0_26_q ;
wire Xd_0__inst_mult_0_27_q ;
wire Xd_0__inst_mult_1_26_q ;
wire Xd_0__inst_mult_1_27_q ;
wire Xd_0__inst_mult_4_28_q ;
wire Xd_0__inst_mult_4_29_q ;
wire Xd_0__inst_mult_5_28_q ;
wire Xd_0__inst_mult_5_29_q ;
wire Xd_0__inst_mult_2_28_q ;
wire Xd_0__inst_mult_2_29_q ;
wire Xd_0__inst_mult_3_28_q ;
wire Xd_0__inst_mult_3_29_q ;
wire Xd_0__inst_mult_0_28_q ;
wire Xd_0__inst_mult_0_29_q ;
wire Xd_0__inst_mult_1_28_q ;
wire Xd_0__inst_mult_1_29_q ;
wire Xd_0__inst_mult_4_30_q ;
wire Xd_0__inst_mult_4_31_q ;
wire Xd_0__inst_mult_5_30_q ;
wire Xd_0__inst_mult_5_31_q ;
wire Xd_0__inst_mult_2_30_q ;
wire Xd_0__inst_mult_2_31_q ;
wire Xd_0__inst_mult_3_30_q ;
wire Xd_0__inst_mult_3_31_q ;
wire Xd_0__inst_mult_0_30_q ;
wire Xd_0__inst_mult_0_31_q ;
wire Xd_0__inst_mult_1_30_q ;
wire Xd_0__inst_mult_1_31_q ;
wire Xd_0__inst_mult_4_32_q ;
wire Xd_0__inst_mult_4_33_q ;
wire Xd_0__inst_mult_5_32_q ;
wire Xd_0__inst_mult_5_33_q ;
wire Xd_0__inst_mult_2_32_q ;
wire Xd_0__inst_mult_2_33_q ;
wire Xd_0__inst_mult_3_32_q ;
wire Xd_0__inst_mult_3_33_q ;
wire Xd_0__inst_mult_0_32_q ;
wire Xd_0__inst_mult_0_33_q ;
wire Xd_0__inst_mult_1_32_q ;
wire Xd_0__inst_mult_1_33_q ;
wire [0:7] Xd_0__inst_sign1 ;
wire [0:7] Xd_0__inst_sign ;
wire [25:0] Xd_0__inst_inst_inst_dout ;
wire [23:0] Xd_0__inst_a1_3__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_2__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_1__adder1_inst_dout ;
wire [23:0] Xd_0__inst_a1_0__adder1_inst_dout ;


twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_inst_inst_add_0_2  = CARRY(( !Xd_0__inst_inst_first_level_0__0__q  $ (!Xd_0__inst_inst_first_level_1__0__q ) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_inst_inst_add_0_3  = SHARE((Xd_0__inst_inst_first_level_0__0__q  & Xd_0__inst_inst_first_level_1__0__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__0__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q ) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_6  = CARRY(( !Xd_0__inst_inst_first_level_0__1__q  $ (!Xd_0__inst_inst_first_level_1__1__q ) ) + ( Xd_0__inst_inst_inst_add_0_3  ) + ( Xd_0__inst_inst_inst_add_0_2  ))
// Xd_0__inst_inst_inst_add_0_7  = SHARE((Xd_0__inst_inst_first_level_0__1__q  & Xd_0__inst_inst_first_level_1__1__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__1__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q ) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_10  = CARRY(( !Xd_0__inst_inst_first_level_0__2__q  $ (!Xd_0__inst_inst_first_level_1__2__q ) ) + ( Xd_0__inst_inst_inst_add_0_7  ) + ( Xd_0__inst_inst_inst_add_0_6  ))
// Xd_0__inst_inst_inst_add_0_11  = SHARE((Xd_0__inst_inst_first_level_0__2__q  & Xd_0__inst_inst_first_level_1__2__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__2__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q ) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_14  = CARRY(( !Xd_0__inst_inst_first_level_0__3__q  $ (!Xd_0__inst_inst_first_level_1__3__q ) ) + ( Xd_0__inst_inst_inst_add_0_11  ) + ( Xd_0__inst_inst_inst_add_0_10  ))
// Xd_0__inst_inst_inst_add_0_15  = SHARE((Xd_0__inst_inst_first_level_0__3__q  & Xd_0__inst_inst_first_level_1__3__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__3__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q ) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_18  = CARRY(( !Xd_0__inst_inst_first_level_0__4__q  $ (!Xd_0__inst_inst_first_level_1__4__q ) ) + ( Xd_0__inst_inst_inst_add_0_15  ) + ( Xd_0__inst_inst_inst_add_0_14  ))
// Xd_0__inst_inst_inst_add_0_19  = SHARE((Xd_0__inst_inst_first_level_0__4__q  & Xd_0__inst_inst_first_level_1__4__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__4__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q ) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_22  = CARRY(( !Xd_0__inst_inst_first_level_0__5__q  $ (!Xd_0__inst_inst_first_level_1__5__q ) ) + ( Xd_0__inst_inst_inst_add_0_19  ) + ( Xd_0__inst_inst_inst_add_0_18  ))
// Xd_0__inst_inst_inst_add_0_23  = SHARE((Xd_0__inst_inst_first_level_0__5__q  & Xd_0__inst_inst_first_level_1__5__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__5__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q ) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_26  = CARRY(( !Xd_0__inst_inst_first_level_0__6__q  $ (!Xd_0__inst_inst_first_level_1__6__q ) ) + ( Xd_0__inst_inst_inst_add_0_23  ) + ( Xd_0__inst_inst_inst_add_0_22  ))
// Xd_0__inst_inst_inst_add_0_27  = SHARE((Xd_0__inst_inst_first_level_0__6__q  & Xd_0__inst_inst_first_level_1__6__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__6__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q ) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_30  = CARRY(( !Xd_0__inst_inst_first_level_0__7__q  $ (!Xd_0__inst_inst_first_level_1__7__q ) ) + ( Xd_0__inst_inst_inst_add_0_27  ) + ( Xd_0__inst_inst_inst_add_0_26  ))
// Xd_0__inst_inst_inst_add_0_31  = SHARE((Xd_0__inst_inst_first_level_0__7__q  & Xd_0__inst_inst_first_level_1__7__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__7__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q ) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_34  = CARRY(( !Xd_0__inst_inst_first_level_0__8__q  $ (!Xd_0__inst_inst_first_level_1__8__q ) ) + ( Xd_0__inst_inst_inst_add_0_31  ) + ( Xd_0__inst_inst_inst_add_0_30  ))
// Xd_0__inst_inst_inst_add_0_35  = SHARE((Xd_0__inst_inst_first_level_0__8__q  & Xd_0__inst_inst_first_level_1__8__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__8__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q ) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_38  = CARRY(( !Xd_0__inst_inst_first_level_0__9__q  $ (!Xd_0__inst_inst_first_level_1__9__q ) ) + ( Xd_0__inst_inst_inst_add_0_35  ) + ( Xd_0__inst_inst_inst_add_0_34  ))
// Xd_0__inst_inst_inst_add_0_39  = SHARE((Xd_0__inst_inst_first_level_0__9__q  & Xd_0__inst_inst_first_level_1__9__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__9__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q ) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_42  = CARRY(( !Xd_0__inst_inst_first_level_0__10__q  $ (!Xd_0__inst_inst_first_level_1__10__q ) ) + ( Xd_0__inst_inst_inst_add_0_39  ) + ( Xd_0__inst_inst_inst_add_0_38  ))
// Xd_0__inst_inst_inst_add_0_43  = SHARE((Xd_0__inst_inst_first_level_0__10__q  & Xd_0__inst_inst_first_level_1__10__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__10__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q ) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_46  = CARRY(( !Xd_0__inst_inst_first_level_0__11__q  $ (!Xd_0__inst_inst_first_level_1__11__q ) ) + ( Xd_0__inst_inst_inst_add_0_43  ) + ( Xd_0__inst_inst_inst_add_0_42  ))
// Xd_0__inst_inst_inst_add_0_47  = SHARE((Xd_0__inst_inst_first_level_0__11__q  & Xd_0__inst_inst_first_level_1__11__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__11__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q ) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_50  = CARRY(( !Xd_0__inst_inst_first_level_0__12__q  $ (!Xd_0__inst_inst_first_level_1__12__q ) ) + ( Xd_0__inst_inst_inst_add_0_47  ) + ( Xd_0__inst_inst_inst_add_0_46  ))
// Xd_0__inst_inst_inst_add_0_51  = SHARE((Xd_0__inst_inst_first_level_0__12__q  & Xd_0__inst_inst_first_level_1__12__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__12__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q ) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_54  = CARRY(( !Xd_0__inst_inst_first_level_0__13__q  $ (!Xd_0__inst_inst_first_level_1__13__q ) ) + ( Xd_0__inst_inst_inst_add_0_51  ) + ( Xd_0__inst_inst_inst_add_0_50  ))
// Xd_0__inst_inst_inst_add_0_55  = SHARE((Xd_0__inst_inst_first_level_0__13__q  & Xd_0__inst_inst_first_level_1__13__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__13__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q ) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_58  = CARRY(( !Xd_0__inst_inst_first_level_0__14__q  $ (!Xd_0__inst_inst_first_level_1__14__q ) ) + ( Xd_0__inst_inst_inst_add_0_55  ) + ( Xd_0__inst_inst_inst_add_0_54  ))
// Xd_0__inst_inst_inst_add_0_59  = SHARE((Xd_0__inst_inst_first_level_0__14__q  & Xd_0__inst_inst_first_level_1__14__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__14__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q ) ) + ( Xd_0__inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_add_0_58  ))
// Xd_0__inst_inst_inst_add_0_62  = CARRY(( !Xd_0__inst_inst_first_level_0__15__q  $ (!Xd_0__inst_inst_first_level_1__15__q ) ) + ( Xd_0__inst_inst_inst_add_0_59  ) + ( Xd_0__inst_inst_inst_add_0_58  ))
// Xd_0__inst_inst_inst_add_0_63  = SHARE((Xd_0__inst_inst_first_level_0__15__q  & Xd_0__inst_inst_first_level_1__15__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__15__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_62 ),
	.shareout(Xd_0__inst_inst_inst_add_0_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_65 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_65_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__16__q  $ (!Xd_0__inst_inst_first_level_1__16__q ) ) + ( Xd_0__inst_inst_inst_add_0_63  ) + ( Xd_0__inst_inst_inst_add_0_62  ))
// Xd_0__inst_inst_inst_add_0_66  = CARRY(( !Xd_0__inst_inst_first_level_0__16__q  $ (!Xd_0__inst_inst_first_level_1__16__q ) ) + ( Xd_0__inst_inst_inst_add_0_63  ) + ( Xd_0__inst_inst_inst_add_0_62  ))
// Xd_0__inst_inst_inst_add_0_67  = SHARE((Xd_0__inst_inst_first_level_0__16__q  & Xd_0__inst_inst_first_level_1__16__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__16__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_62 ),
	.sharein(Xd_0__inst_inst_inst_add_0_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_65_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_66 ),
	.shareout(Xd_0__inst_inst_inst_add_0_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_69 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_69_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__17__q  $ (!Xd_0__inst_inst_first_level_1__17__q ) ) + ( Xd_0__inst_inst_inst_add_0_67  ) + ( Xd_0__inst_inst_inst_add_0_66  ))
// Xd_0__inst_inst_inst_add_0_70  = CARRY(( !Xd_0__inst_inst_first_level_0__17__q  $ (!Xd_0__inst_inst_first_level_1__17__q ) ) + ( Xd_0__inst_inst_inst_add_0_67  ) + ( Xd_0__inst_inst_inst_add_0_66  ))
// Xd_0__inst_inst_inst_add_0_71  = SHARE((Xd_0__inst_inst_first_level_0__17__q  & Xd_0__inst_inst_first_level_1__17__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__17__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_66 ),
	.sharein(Xd_0__inst_inst_inst_add_0_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_69_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_70 ),
	.shareout(Xd_0__inst_inst_inst_add_0_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_73 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_73_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__18__q  $ (!Xd_0__inst_inst_first_level_1__18__q ) ) + ( Xd_0__inst_inst_inst_add_0_71  ) + ( Xd_0__inst_inst_inst_add_0_70  ))
// Xd_0__inst_inst_inst_add_0_74  = CARRY(( !Xd_0__inst_inst_first_level_0__18__q  $ (!Xd_0__inst_inst_first_level_1__18__q ) ) + ( Xd_0__inst_inst_inst_add_0_71  ) + ( Xd_0__inst_inst_inst_add_0_70  ))
// Xd_0__inst_inst_inst_add_0_75  = SHARE((Xd_0__inst_inst_first_level_0__18__q  & Xd_0__inst_inst_first_level_1__18__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__18__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_70 ),
	.sharein(Xd_0__inst_inst_inst_add_0_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_73_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_74 ),
	.shareout(Xd_0__inst_inst_inst_add_0_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_77 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_77_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__19__q  $ (!Xd_0__inst_inst_first_level_1__19__q ) ) + ( Xd_0__inst_inst_inst_add_0_75  ) + ( Xd_0__inst_inst_inst_add_0_74  ))
// Xd_0__inst_inst_inst_add_0_78  = CARRY(( !Xd_0__inst_inst_first_level_0__19__q  $ (!Xd_0__inst_inst_first_level_1__19__q ) ) + ( Xd_0__inst_inst_inst_add_0_75  ) + ( Xd_0__inst_inst_inst_add_0_74  ))
// Xd_0__inst_inst_inst_add_0_79  = SHARE((Xd_0__inst_inst_first_level_0__19__q  & Xd_0__inst_inst_first_level_1__19__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__19__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_74 ),
	.sharein(Xd_0__inst_inst_inst_add_0_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_77_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_78 ),
	.shareout(Xd_0__inst_inst_inst_add_0_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_81 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_81_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__20__q  $ (!Xd_0__inst_inst_first_level_1__20__q ) ) + ( Xd_0__inst_inst_inst_add_0_79  ) + ( Xd_0__inst_inst_inst_add_0_78  ))
// Xd_0__inst_inst_inst_add_0_82  = CARRY(( !Xd_0__inst_inst_first_level_0__20__q  $ (!Xd_0__inst_inst_first_level_1__20__q ) ) + ( Xd_0__inst_inst_inst_add_0_79  ) + ( Xd_0__inst_inst_inst_add_0_78  ))
// Xd_0__inst_inst_inst_add_0_83  = SHARE((Xd_0__inst_inst_first_level_0__20__q  & Xd_0__inst_inst_first_level_1__20__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__20__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_78 ),
	.sharein(Xd_0__inst_inst_inst_add_0_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_82 ),
	.shareout(Xd_0__inst_inst_inst_add_0_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_85 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_85_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__21__q  $ (!Xd_0__inst_inst_first_level_1__21__q ) ) + ( Xd_0__inst_inst_inst_add_0_83  ) + ( Xd_0__inst_inst_inst_add_0_82  ))
// Xd_0__inst_inst_inst_add_0_86  = CARRY(( !Xd_0__inst_inst_first_level_0__21__q  $ (!Xd_0__inst_inst_first_level_1__21__q ) ) + ( Xd_0__inst_inst_inst_add_0_83  ) + ( Xd_0__inst_inst_inst_add_0_82  ))
// Xd_0__inst_inst_inst_add_0_87  = SHARE((Xd_0__inst_inst_first_level_0__21__q  & Xd_0__inst_inst_first_level_1__21__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__21__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_82 ),
	.sharein(Xd_0__inst_inst_inst_add_0_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_85_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_86 ),
	.shareout(Xd_0__inst_inst_inst_add_0_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_89 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_89_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__22__q  $ (!Xd_0__inst_inst_first_level_1__22__q ) ) + ( Xd_0__inst_inst_inst_add_0_87  ) + ( Xd_0__inst_inst_inst_add_0_86  ))
// Xd_0__inst_inst_inst_add_0_90  = CARRY(( !Xd_0__inst_inst_first_level_0__22__q  $ (!Xd_0__inst_inst_first_level_1__22__q ) ) + ( Xd_0__inst_inst_inst_add_0_87  ) + ( Xd_0__inst_inst_inst_add_0_86  ))
// Xd_0__inst_inst_inst_add_0_91  = SHARE((Xd_0__inst_inst_first_level_0__22__q  & Xd_0__inst_inst_first_level_1__22__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__22__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_86 ),
	.sharein(Xd_0__inst_inst_inst_add_0_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_89_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_90 ),
	.shareout(Xd_0__inst_inst_inst_add_0_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_93 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_93_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__23__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_91  ) + ( Xd_0__inst_inst_inst_add_0_90  ))
// Xd_0__inst_inst_inst_add_0_94  = CARRY(( !Xd_0__inst_inst_first_level_0__23__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_91  ) + ( Xd_0__inst_inst_inst_add_0_90  ))
// Xd_0__inst_inst_inst_add_0_95  = SHARE((Xd_0__inst_inst_first_level_0__23__q  & Xd_0__inst_inst_first_level_1__25__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__23__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_90 ),
	.sharein(Xd_0__inst_inst_inst_add_0_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_93_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_94 ),
	.shareout(Xd_0__inst_inst_inst_add_0_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00000055000055AA),
	.shared_arith("on")
) Xd_0__inst_inst_inst_add_0_97 (
// Equation(s):
// Xd_0__inst_inst_inst_add_0_97_sumout  = SUM(( !Xd_0__inst_inst_first_level_0__24__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_95  ) + ( Xd_0__inst_inst_inst_add_0_94  ))
// Xd_0__inst_inst_inst_add_0_98  = CARRY(( !Xd_0__inst_inst_first_level_0__24__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_95  ) + ( Xd_0__inst_inst_inst_add_0_94  ))
// Xd_0__inst_inst_inst_add_0_99  = SHARE((Xd_0__inst_inst_first_level_0__24__q  & Xd_0__inst_inst_first_level_1__25__q ))

	.dataa(!Xd_0__inst_inst_first_level_0__24__q ),
	.datab(gnd),
	.datac(gnd),
	.datad(!Xd_0__inst_inst_first_level_1__25__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_94 ),
	.sharein(Xd_0__inst_inst_inst_add_0_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_inst_add_0_97_sumout ),
	.cout(Xd_0__inst_inst_inst_add_0_98 ),
	.shareout(Xd_0__inst_inst_inst_add_0_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_168 (
// Equation(s):
// Xd_0__inst_mult_1_169  = SUM(( !Xd_0__inst_inst_first_level_0__25__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_99  ) + ( Xd_0__inst_inst_inst_add_0_98  ))
// Xd_0__inst_mult_1_170  = CARRY(( !Xd_0__inst_inst_first_level_0__25__q  $ (!Xd_0__inst_inst_first_level_1__25__q ) ) + ( Xd_0__inst_inst_inst_add_0_99  ) + ( Xd_0__inst_inst_inst_add_0_98  ))
// Xd_0__inst_mult_1_171  = SHARE(Xd_0__inst_mult_1_173 )

	.dataa(!Xd_0__inst_inst_first_level_0__25__q ),
	.datab(!Xd_0__inst_inst_first_level_1__25__q ),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_1_173 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_inst_add_0_98 ),
	.sharein(Xd_0__inst_inst_inst_add_0_99 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_169 ),
	.cout(Xd_0__inst_mult_1_170 ),
	.shareout(Xd_0__inst_mult_1_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1 (
// Equation(s):
// Xd_0__inst_mult_1_173  = SUM(( (!din_a[14] & (((din_a[15] & din_b[12])))) # (din_a[14] & (!din_b[13] $ (((!din_a[15]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_178  ) + ( Xd_0__inst_mult_1_177  ))
// Xd_0__inst_mult_1_174  = CARRY(( (!din_a[14] & (((din_a[15] & din_b[12])))) # (din_a[14] & (!din_b[13] $ (((!din_a[15]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_178  ) + ( Xd_0__inst_mult_1_177  ))
// Xd_0__inst_mult_1_175  = SHARE((din_a[14] & (din_b[13] & (din_a[15] & din_b[12]))))

	.dataa(!din_a[14]),
	.datab(!din_b[13]),
	.datac(!din_a[15]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_177 ),
	.sharein(Xd_0__inst_mult_1_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_173 ),
	.cout(Xd_0__inst_mult_1_174 ),
	.shareout(Xd_0__inst_mult_1_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_1 (
// Equation(s):
// Xd_0__inst_inst_add_0_1_sumout  = SUM(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_3_171  ) + ( Xd_0__inst_mult_3_170  ))
// Xd_0__inst_inst_add_0_2  = CARRY(( !Xd_0__inst_r_sum1_2__0__q  $ (!Xd_0__inst_r_sum1_1__0__q  $ (Xd_0__inst_r_sum1_0__0__q )) ) + ( Xd_0__inst_mult_3_171  ) + ( Xd_0__inst_mult_3_170  ))
// Xd_0__inst_inst_add_0_3  = SHARE((!Xd_0__inst_r_sum1_2__0__q  & (Xd_0__inst_r_sum1_1__0__q  & Xd_0__inst_r_sum1_0__0__q )) # (Xd_0__inst_r_sum1_2__0__q  & ((Xd_0__inst_r_sum1_0__0__q ) # (Xd_0__inst_r_sum1_1__0__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__0__q ),
	.datac(!Xd_0__inst_r_sum1_1__0__q ),
	.datad(!Xd_0__inst_r_sum1_0__0__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_170 ),
	.sharein(Xd_0__inst_mult_3_171 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_1_sumout ),
	.cout(Xd_0__inst_inst_add_0_2 ),
	.shareout(Xd_0__inst_inst_add_0_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_5 (
// Equation(s):
// Xd_0__inst_inst_add_0_5_sumout  = SUM(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_6  = CARRY(( !Xd_0__inst_r_sum1_2__1__q  $ (!Xd_0__inst_r_sum1_1__1__q  $ (Xd_0__inst_r_sum1_0__1__q )) ) + ( Xd_0__inst_inst_add_0_3  ) + ( Xd_0__inst_inst_add_0_2  ))
// Xd_0__inst_inst_add_0_7  = SHARE((!Xd_0__inst_r_sum1_2__1__q  & (Xd_0__inst_r_sum1_1__1__q  & Xd_0__inst_r_sum1_0__1__q )) # (Xd_0__inst_r_sum1_2__1__q  & ((Xd_0__inst_r_sum1_0__1__q ) # (Xd_0__inst_r_sum1_1__1__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__1__q ),
	.datac(!Xd_0__inst_r_sum1_1__1__q ),
	.datad(!Xd_0__inst_r_sum1_0__1__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_2 ),
	.sharein(Xd_0__inst_inst_add_0_3 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_5_sumout ),
	.cout(Xd_0__inst_inst_add_0_6 ),
	.shareout(Xd_0__inst_inst_add_0_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_9 (
// Equation(s):
// Xd_0__inst_inst_add_0_9_sumout  = SUM(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_10  = CARRY(( !Xd_0__inst_r_sum1_2__2__q  $ (!Xd_0__inst_r_sum1_1__2__q  $ (Xd_0__inst_r_sum1_0__2__q )) ) + ( Xd_0__inst_inst_add_0_7  ) + ( Xd_0__inst_inst_add_0_6  ))
// Xd_0__inst_inst_add_0_11  = SHARE((!Xd_0__inst_r_sum1_2__2__q  & (Xd_0__inst_r_sum1_1__2__q  & Xd_0__inst_r_sum1_0__2__q )) # (Xd_0__inst_r_sum1_2__2__q  & ((Xd_0__inst_r_sum1_0__2__q ) # (Xd_0__inst_r_sum1_1__2__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__2__q ),
	.datac(!Xd_0__inst_r_sum1_1__2__q ),
	.datad(!Xd_0__inst_r_sum1_0__2__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_6 ),
	.sharein(Xd_0__inst_inst_add_0_7 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_9_sumout ),
	.cout(Xd_0__inst_inst_add_0_10 ),
	.shareout(Xd_0__inst_inst_add_0_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_13 (
// Equation(s):
// Xd_0__inst_inst_add_0_13_sumout  = SUM(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_14  = CARRY(( !Xd_0__inst_r_sum1_2__3__q  $ (!Xd_0__inst_r_sum1_1__3__q  $ (Xd_0__inst_r_sum1_0__3__q )) ) + ( Xd_0__inst_inst_add_0_11  ) + ( Xd_0__inst_inst_add_0_10  ))
// Xd_0__inst_inst_add_0_15  = SHARE((!Xd_0__inst_r_sum1_2__3__q  & (Xd_0__inst_r_sum1_1__3__q  & Xd_0__inst_r_sum1_0__3__q )) # (Xd_0__inst_r_sum1_2__3__q  & ((Xd_0__inst_r_sum1_0__3__q ) # (Xd_0__inst_r_sum1_1__3__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__3__q ),
	.datac(!Xd_0__inst_r_sum1_1__3__q ),
	.datad(!Xd_0__inst_r_sum1_0__3__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_10 ),
	.sharein(Xd_0__inst_inst_add_0_11 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_13_sumout ),
	.cout(Xd_0__inst_inst_add_0_14 ),
	.shareout(Xd_0__inst_inst_add_0_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_17 (
// Equation(s):
// Xd_0__inst_inst_add_0_17_sumout  = SUM(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_18  = CARRY(( !Xd_0__inst_r_sum1_2__4__q  $ (!Xd_0__inst_r_sum1_1__4__q  $ (Xd_0__inst_r_sum1_0__4__q )) ) + ( Xd_0__inst_inst_add_0_15  ) + ( Xd_0__inst_inst_add_0_14  ))
// Xd_0__inst_inst_add_0_19  = SHARE((!Xd_0__inst_r_sum1_2__4__q  & (Xd_0__inst_r_sum1_1__4__q  & Xd_0__inst_r_sum1_0__4__q )) # (Xd_0__inst_r_sum1_2__4__q  & ((Xd_0__inst_r_sum1_0__4__q ) # (Xd_0__inst_r_sum1_1__4__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__4__q ),
	.datac(!Xd_0__inst_r_sum1_1__4__q ),
	.datad(!Xd_0__inst_r_sum1_0__4__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_14 ),
	.sharein(Xd_0__inst_inst_add_0_15 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_17_sumout ),
	.cout(Xd_0__inst_inst_add_0_18 ),
	.shareout(Xd_0__inst_inst_add_0_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_21 (
// Equation(s):
// Xd_0__inst_inst_add_0_21_sumout  = SUM(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_22  = CARRY(( !Xd_0__inst_r_sum1_2__5__q  $ (!Xd_0__inst_r_sum1_1__5__q  $ (Xd_0__inst_r_sum1_0__5__q )) ) + ( Xd_0__inst_inst_add_0_19  ) + ( Xd_0__inst_inst_add_0_18  ))
// Xd_0__inst_inst_add_0_23  = SHARE((!Xd_0__inst_r_sum1_2__5__q  & (Xd_0__inst_r_sum1_1__5__q  & Xd_0__inst_r_sum1_0__5__q )) # (Xd_0__inst_r_sum1_2__5__q  & ((Xd_0__inst_r_sum1_0__5__q ) # (Xd_0__inst_r_sum1_1__5__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__5__q ),
	.datac(!Xd_0__inst_r_sum1_1__5__q ),
	.datad(!Xd_0__inst_r_sum1_0__5__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_18 ),
	.sharein(Xd_0__inst_inst_add_0_19 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_21_sumout ),
	.cout(Xd_0__inst_inst_add_0_22 ),
	.shareout(Xd_0__inst_inst_add_0_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_25 (
// Equation(s):
// Xd_0__inst_inst_add_0_25_sumout  = SUM(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_26  = CARRY(( !Xd_0__inst_r_sum1_2__6__q  $ (!Xd_0__inst_r_sum1_1__6__q  $ (Xd_0__inst_r_sum1_0__6__q )) ) + ( Xd_0__inst_inst_add_0_23  ) + ( Xd_0__inst_inst_add_0_22  ))
// Xd_0__inst_inst_add_0_27  = SHARE((!Xd_0__inst_r_sum1_2__6__q  & (Xd_0__inst_r_sum1_1__6__q  & Xd_0__inst_r_sum1_0__6__q )) # (Xd_0__inst_r_sum1_2__6__q  & ((Xd_0__inst_r_sum1_0__6__q ) # (Xd_0__inst_r_sum1_1__6__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__6__q ),
	.datac(!Xd_0__inst_r_sum1_1__6__q ),
	.datad(!Xd_0__inst_r_sum1_0__6__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_22 ),
	.sharein(Xd_0__inst_inst_add_0_23 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_25_sumout ),
	.cout(Xd_0__inst_inst_add_0_26 ),
	.shareout(Xd_0__inst_inst_add_0_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_29 (
// Equation(s):
// Xd_0__inst_inst_add_0_29_sumout  = SUM(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_30  = CARRY(( !Xd_0__inst_r_sum1_2__7__q  $ (!Xd_0__inst_r_sum1_1__7__q  $ (Xd_0__inst_r_sum1_0__7__q )) ) + ( Xd_0__inst_inst_add_0_27  ) + ( Xd_0__inst_inst_add_0_26  ))
// Xd_0__inst_inst_add_0_31  = SHARE((!Xd_0__inst_r_sum1_2__7__q  & (Xd_0__inst_r_sum1_1__7__q  & Xd_0__inst_r_sum1_0__7__q )) # (Xd_0__inst_r_sum1_2__7__q  & ((Xd_0__inst_r_sum1_0__7__q ) # (Xd_0__inst_r_sum1_1__7__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__7__q ),
	.datac(!Xd_0__inst_r_sum1_1__7__q ),
	.datad(!Xd_0__inst_r_sum1_0__7__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_26 ),
	.sharein(Xd_0__inst_inst_add_0_27 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_29_sumout ),
	.cout(Xd_0__inst_inst_add_0_30 ),
	.shareout(Xd_0__inst_inst_add_0_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_33 (
// Equation(s):
// Xd_0__inst_inst_add_0_33_sumout  = SUM(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_34  = CARRY(( !Xd_0__inst_r_sum1_2__8__q  $ (!Xd_0__inst_r_sum1_1__8__q  $ (Xd_0__inst_r_sum1_0__8__q )) ) + ( Xd_0__inst_inst_add_0_31  ) + ( Xd_0__inst_inst_add_0_30  ))
// Xd_0__inst_inst_add_0_35  = SHARE((!Xd_0__inst_r_sum1_2__8__q  & (Xd_0__inst_r_sum1_1__8__q  & Xd_0__inst_r_sum1_0__8__q )) # (Xd_0__inst_r_sum1_2__8__q  & ((Xd_0__inst_r_sum1_0__8__q ) # (Xd_0__inst_r_sum1_1__8__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__8__q ),
	.datac(!Xd_0__inst_r_sum1_1__8__q ),
	.datad(!Xd_0__inst_r_sum1_0__8__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_30 ),
	.sharein(Xd_0__inst_inst_add_0_31 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_33_sumout ),
	.cout(Xd_0__inst_inst_add_0_34 ),
	.shareout(Xd_0__inst_inst_add_0_35 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_37 (
// Equation(s):
// Xd_0__inst_inst_add_0_37_sumout  = SUM(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_38  = CARRY(( !Xd_0__inst_r_sum1_2__9__q  $ (!Xd_0__inst_r_sum1_1__9__q  $ (Xd_0__inst_r_sum1_0__9__q )) ) + ( Xd_0__inst_inst_add_0_35  ) + ( Xd_0__inst_inst_add_0_34  ))
// Xd_0__inst_inst_add_0_39  = SHARE((!Xd_0__inst_r_sum1_2__9__q  & (Xd_0__inst_r_sum1_1__9__q  & Xd_0__inst_r_sum1_0__9__q )) # (Xd_0__inst_r_sum1_2__9__q  & ((Xd_0__inst_r_sum1_0__9__q ) # (Xd_0__inst_r_sum1_1__9__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__9__q ),
	.datac(!Xd_0__inst_r_sum1_1__9__q ),
	.datad(!Xd_0__inst_r_sum1_0__9__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_34 ),
	.sharein(Xd_0__inst_inst_add_0_35 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_37_sumout ),
	.cout(Xd_0__inst_inst_add_0_38 ),
	.shareout(Xd_0__inst_inst_add_0_39 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_41 (
// Equation(s):
// Xd_0__inst_inst_add_0_41_sumout  = SUM(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_42  = CARRY(( !Xd_0__inst_r_sum1_2__10__q  $ (!Xd_0__inst_r_sum1_1__10__q  $ (Xd_0__inst_r_sum1_0__10__q )) ) + ( Xd_0__inst_inst_add_0_39  ) + ( Xd_0__inst_inst_add_0_38  ))
// Xd_0__inst_inst_add_0_43  = SHARE((!Xd_0__inst_r_sum1_2__10__q  & (Xd_0__inst_r_sum1_1__10__q  & Xd_0__inst_r_sum1_0__10__q )) # (Xd_0__inst_r_sum1_2__10__q  & ((Xd_0__inst_r_sum1_0__10__q ) # (Xd_0__inst_r_sum1_1__10__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__10__q ),
	.datac(!Xd_0__inst_r_sum1_1__10__q ),
	.datad(!Xd_0__inst_r_sum1_0__10__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_38 ),
	.sharein(Xd_0__inst_inst_add_0_39 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_41_sumout ),
	.cout(Xd_0__inst_inst_add_0_42 ),
	.shareout(Xd_0__inst_inst_add_0_43 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_45 (
// Equation(s):
// Xd_0__inst_inst_add_0_45_sumout  = SUM(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_46  = CARRY(( !Xd_0__inst_r_sum1_2__11__q  $ (!Xd_0__inst_r_sum1_1__11__q  $ (Xd_0__inst_r_sum1_0__11__q )) ) + ( Xd_0__inst_inst_add_0_43  ) + ( Xd_0__inst_inst_add_0_42  ))
// Xd_0__inst_inst_add_0_47  = SHARE((!Xd_0__inst_r_sum1_2__11__q  & (Xd_0__inst_r_sum1_1__11__q  & Xd_0__inst_r_sum1_0__11__q )) # (Xd_0__inst_r_sum1_2__11__q  & ((Xd_0__inst_r_sum1_0__11__q ) # (Xd_0__inst_r_sum1_1__11__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__11__q ),
	.datac(!Xd_0__inst_r_sum1_1__11__q ),
	.datad(!Xd_0__inst_r_sum1_0__11__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_42 ),
	.sharein(Xd_0__inst_inst_add_0_43 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_45_sumout ),
	.cout(Xd_0__inst_inst_add_0_46 ),
	.shareout(Xd_0__inst_inst_add_0_47 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_49 (
// Equation(s):
// Xd_0__inst_inst_add_0_49_sumout  = SUM(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_50  = CARRY(( !Xd_0__inst_r_sum1_2__12__q  $ (!Xd_0__inst_r_sum1_1__12__q  $ (Xd_0__inst_r_sum1_0__12__q )) ) + ( Xd_0__inst_inst_add_0_47  ) + ( Xd_0__inst_inst_add_0_46  ))
// Xd_0__inst_inst_add_0_51  = SHARE((!Xd_0__inst_r_sum1_2__12__q  & (Xd_0__inst_r_sum1_1__12__q  & Xd_0__inst_r_sum1_0__12__q )) # (Xd_0__inst_r_sum1_2__12__q  & ((Xd_0__inst_r_sum1_0__12__q ) # (Xd_0__inst_r_sum1_1__12__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__12__q ),
	.datac(!Xd_0__inst_r_sum1_1__12__q ),
	.datad(!Xd_0__inst_r_sum1_0__12__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_46 ),
	.sharein(Xd_0__inst_inst_add_0_47 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_49_sumout ),
	.cout(Xd_0__inst_inst_add_0_50 ),
	.shareout(Xd_0__inst_inst_add_0_51 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_53 (
// Equation(s):
// Xd_0__inst_inst_add_0_53_sumout  = SUM(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_54  = CARRY(( !Xd_0__inst_r_sum1_2__13__q  $ (!Xd_0__inst_r_sum1_1__13__q  $ (Xd_0__inst_r_sum1_0__13__q )) ) + ( Xd_0__inst_inst_add_0_51  ) + ( Xd_0__inst_inst_add_0_50  ))
// Xd_0__inst_inst_add_0_55  = SHARE((!Xd_0__inst_r_sum1_2__13__q  & (Xd_0__inst_r_sum1_1__13__q  & Xd_0__inst_r_sum1_0__13__q )) # (Xd_0__inst_r_sum1_2__13__q  & ((Xd_0__inst_r_sum1_0__13__q ) # (Xd_0__inst_r_sum1_1__13__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__13__q ),
	.datac(!Xd_0__inst_r_sum1_1__13__q ),
	.datad(!Xd_0__inst_r_sum1_0__13__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_50 ),
	.sharein(Xd_0__inst_inst_add_0_51 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_53_sumout ),
	.cout(Xd_0__inst_inst_add_0_54 ),
	.shareout(Xd_0__inst_inst_add_0_55 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_57 (
// Equation(s):
// Xd_0__inst_inst_add_0_57_sumout  = SUM(( !Xd_0__inst_r_sum1_2__14__q  $ (!Xd_0__inst_r_sum1_1__14__q  $ (Xd_0__inst_r_sum1_0__14__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_58  = CARRY(( !Xd_0__inst_r_sum1_2__14__q  $ (!Xd_0__inst_r_sum1_1__14__q  $ (Xd_0__inst_r_sum1_0__14__q )) ) + ( Xd_0__inst_inst_add_0_55  ) + ( Xd_0__inst_inst_add_0_54  ))
// Xd_0__inst_inst_add_0_59  = SHARE((!Xd_0__inst_r_sum1_2__14__q  & (Xd_0__inst_r_sum1_1__14__q  & Xd_0__inst_r_sum1_0__14__q )) # (Xd_0__inst_r_sum1_2__14__q  & ((Xd_0__inst_r_sum1_0__14__q ) # (Xd_0__inst_r_sum1_1__14__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__14__q ),
	.datac(!Xd_0__inst_r_sum1_1__14__q ),
	.datad(!Xd_0__inst_r_sum1_0__14__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_54 ),
	.sharein(Xd_0__inst_inst_add_0_55 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_57_sumout ),
	.cout(Xd_0__inst_inst_add_0_58 ),
	.shareout(Xd_0__inst_inst_add_0_59 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_61 (
// Equation(s):
// Xd_0__inst_inst_add_0_61_sumout  = SUM(( !Xd_0__inst_r_sum1_2__15__q  $ (!Xd_0__inst_r_sum1_1__15__q  $ (Xd_0__inst_r_sum1_0__15__q )) ) + ( Xd_0__inst_inst_add_0_59  ) + ( Xd_0__inst_inst_add_0_58  ))
// Xd_0__inst_inst_add_0_62  = CARRY(( !Xd_0__inst_r_sum1_2__15__q  $ (!Xd_0__inst_r_sum1_1__15__q  $ (Xd_0__inst_r_sum1_0__15__q )) ) + ( Xd_0__inst_inst_add_0_59  ) + ( Xd_0__inst_inst_add_0_58  ))
// Xd_0__inst_inst_add_0_63  = SHARE((!Xd_0__inst_r_sum1_2__15__q  & (Xd_0__inst_r_sum1_1__15__q  & Xd_0__inst_r_sum1_0__15__q )) # (Xd_0__inst_r_sum1_2__15__q  & ((Xd_0__inst_r_sum1_0__15__q ) # (Xd_0__inst_r_sum1_1__15__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__15__q ),
	.datac(!Xd_0__inst_r_sum1_1__15__q ),
	.datad(!Xd_0__inst_r_sum1_0__15__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_58 ),
	.sharein(Xd_0__inst_inst_add_0_59 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_61_sumout ),
	.cout(Xd_0__inst_inst_add_0_62 ),
	.shareout(Xd_0__inst_inst_add_0_63 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_65 (
// Equation(s):
// Xd_0__inst_inst_add_0_65_sumout  = SUM(( !Xd_0__inst_r_sum1_2__16__q  $ (!Xd_0__inst_r_sum1_1__16__q  $ (Xd_0__inst_r_sum1_0__16__q )) ) + ( Xd_0__inst_inst_add_0_63  ) + ( Xd_0__inst_inst_add_0_62  ))
// Xd_0__inst_inst_add_0_66  = CARRY(( !Xd_0__inst_r_sum1_2__16__q  $ (!Xd_0__inst_r_sum1_1__16__q  $ (Xd_0__inst_r_sum1_0__16__q )) ) + ( Xd_0__inst_inst_add_0_63  ) + ( Xd_0__inst_inst_add_0_62  ))
// Xd_0__inst_inst_add_0_67  = SHARE((!Xd_0__inst_r_sum1_2__16__q  & (Xd_0__inst_r_sum1_1__16__q  & Xd_0__inst_r_sum1_0__16__q )) # (Xd_0__inst_r_sum1_2__16__q  & ((Xd_0__inst_r_sum1_0__16__q ) # (Xd_0__inst_r_sum1_1__16__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__16__q ),
	.datac(!Xd_0__inst_r_sum1_1__16__q ),
	.datad(!Xd_0__inst_r_sum1_0__16__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_62 ),
	.sharein(Xd_0__inst_inst_add_0_63 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_65_sumout ),
	.cout(Xd_0__inst_inst_add_0_66 ),
	.shareout(Xd_0__inst_inst_add_0_67 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_69 (
// Equation(s):
// Xd_0__inst_inst_add_0_69_sumout  = SUM(( !Xd_0__inst_r_sum1_2__17__q  $ (!Xd_0__inst_r_sum1_1__17__q  $ (Xd_0__inst_r_sum1_0__17__q )) ) + ( Xd_0__inst_inst_add_0_67  ) + ( Xd_0__inst_inst_add_0_66  ))
// Xd_0__inst_inst_add_0_70  = CARRY(( !Xd_0__inst_r_sum1_2__17__q  $ (!Xd_0__inst_r_sum1_1__17__q  $ (Xd_0__inst_r_sum1_0__17__q )) ) + ( Xd_0__inst_inst_add_0_67  ) + ( Xd_0__inst_inst_add_0_66  ))
// Xd_0__inst_inst_add_0_71  = SHARE((!Xd_0__inst_r_sum1_2__17__q  & (Xd_0__inst_r_sum1_1__17__q  & Xd_0__inst_r_sum1_0__17__q )) # (Xd_0__inst_r_sum1_2__17__q  & ((Xd_0__inst_r_sum1_0__17__q ) # (Xd_0__inst_r_sum1_1__17__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__17__q ),
	.datac(!Xd_0__inst_r_sum1_1__17__q ),
	.datad(!Xd_0__inst_r_sum1_0__17__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_66 ),
	.sharein(Xd_0__inst_inst_add_0_67 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_69_sumout ),
	.cout(Xd_0__inst_inst_add_0_70 ),
	.shareout(Xd_0__inst_inst_add_0_71 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_73 (
// Equation(s):
// Xd_0__inst_inst_add_0_73_sumout  = SUM(( !Xd_0__inst_r_sum1_2__18__q  $ (!Xd_0__inst_r_sum1_1__18__q  $ (Xd_0__inst_r_sum1_0__18__q )) ) + ( Xd_0__inst_inst_add_0_71  ) + ( Xd_0__inst_inst_add_0_70  ))
// Xd_0__inst_inst_add_0_74  = CARRY(( !Xd_0__inst_r_sum1_2__18__q  $ (!Xd_0__inst_r_sum1_1__18__q  $ (Xd_0__inst_r_sum1_0__18__q )) ) + ( Xd_0__inst_inst_add_0_71  ) + ( Xd_0__inst_inst_add_0_70  ))
// Xd_0__inst_inst_add_0_75  = SHARE((!Xd_0__inst_r_sum1_2__18__q  & (Xd_0__inst_r_sum1_1__18__q  & Xd_0__inst_r_sum1_0__18__q )) # (Xd_0__inst_r_sum1_2__18__q  & ((Xd_0__inst_r_sum1_0__18__q ) # (Xd_0__inst_r_sum1_1__18__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__18__q ),
	.datac(!Xd_0__inst_r_sum1_1__18__q ),
	.datad(!Xd_0__inst_r_sum1_0__18__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_70 ),
	.sharein(Xd_0__inst_inst_add_0_71 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_73_sumout ),
	.cout(Xd_0__inst_inst_add_0_74 ),
	.shareout(Xd_0__inst_inst_add_0_75 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_77 (
// Equation(s):
// Xd_0__inst_inst_add_0_77_sumout  = SUM(( !Xd_0__inst_r_sum1_2__19__q  $ (!Xd_0__inst_r_sum1_1__19__q  $ (Xd_0__inst_r_sum1_0__19__q )) ) + ( Xd_0__inst_inst_add_0_75  ) + ( Xd_0__inst_inst_add_0_74  ))
// Xd_0__inst_inst_add_0_78  = CARRY(( !Xd_0__inst_r_sum1_2__19__q  $ (!Xd_0__inst_r_sum1_1__19__q  $ (Xd_0__inst_r_sum1_0__19__q )) ) + ( Xd_0__inst_inst_add_0_75  ) + ( Xd_0__inst_inst_add_0_74  ))
// Xd_0__inst_inst_add_0_79  = SHARE((!Xd_0__inst_r_sum1_2__19__q  & (Xd_0__inst_r_sum1_1__19__q  & Xd_0__inst_r_sum1_0__19__q )) # (Xd_0__inst_r_sum1_2__19__q  & ((Xd_0__inst_r_sum1_0__19__q ) # (Xd_0__inst_r_sum1_1__19__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__19__q ),
	.datac(!Xd_0__inst_r_sum1_1__19__q ),
	.datad(!Xd_0__inst_r_sum1_0__19__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_74 ),
	.sharein(Xd_0__inst_inst_add_0_75 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_77_sumout ),
	.cout(Xd_0__inst_inst_add_0_78 ),
	.shareout(Xd_0__inst_inst_add_0_79 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_81 (
// Equation(s):
// Xd_0__inst_inst_add_0_81_sumout  = SUM(( !Xd_0__inst_r_sum1_2__20__q  $ (!Xd_0__inst_r_sum1_1__20__q  $ (Xd_0__inst_r_sum1_0__20__q )) ) + ( Xd_0__inst_inst_add_0_79  ) + ( Xd_0__inst_inst_add_0_78  ))
// Xd_0__inst_inst_add_0_82  = CARRY(( !Xd_0__inst_r_sum1_2__20__q  $ (!Xd_0__inst_r_sum1_1__20__q  $ (Xd_0__inst_r_sum1_0__20__q )) ) + ( Xd_0__inst_inst_add_0_79  ) + ( Xd_0__inst_inst_add_0_78  ))
// Xd_0__inst_inst_add_0_83  = SHARE((!Xd_0__inst_r_sum1_2__20__q  & (Xd_0__inst_r_sum1_1__20__q  & Xd_0__inst_r_sum1_0__20__q )) # (Xd_0__inst_r_sum1_2__20__q  & ((Xd_0__inst_r_sum1_0__20__q ) # (Xd_0__inst_r_sum1_1__20__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__20__q ),
	.datac(!Xd_0__inst_r_sum1_1__20__q ),
	.datad(!Xd_0__inst_r_sum1_0__20__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_78 ),
	.sharein(Xd_0__inst_inst_add_0_79 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_81_sumout ),
	.cout(Xd_0__inst_inst_add_0_82 ),
	.shareout(Xd_0__inst_inst_add_0_83 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_85 (
// Equation(s):
// Xd_0__inst_inst_add_0_85_sumout  = SUM(( !Xd_0__inst_r_sum1_2__21__q  $ (!Xd_0__inst_r_sum1_1__21__q  $ (Xd_0__inst_r_sum1_0__21__q )) ) + ( Xd_0__inst_inst_add_0_83  ) + ( Xd_0__inst_inst_add_0_82  ))
// Xd_0__inst_inst_add_0_86  = CARRY(( !Xd_0__inst_r_sum1_2__21__q  $ (!Xd_0__inst_r_sum1_1__21__q  $ (Xd_0__inst_r_sum1_0__21__q )) ) + ( Xd_0__inst_inst_add_0_83  ) + ( Xd_0__inst_inst_add_0_82  ))
// Xd_0__inst_inst_add_0_87  = SHARE((!Xd_0__inst_r_sum1_2__21__q  & (Xd_0__inst_r_sum1_1__21__q  & Xd_0__inst_r_sum1_0__21__q )) # (Xd_0__inst_r_sum1_2__21__q  & ((Xd_0__inst_r_sum1_0__21__q ) # (Xd_0__inst_r_sum1_1__21__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__21__q ),
	.datac(!Xd_0__inst_r_sum1_1__21__q ),
	.datad(!Xd_0__inst_r_sum1_0__21__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_82 ),
	.sharein(Xd_0__inst_inst_add_0_83 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_85_sumout ),
	.cout(Xd_0__inst_inst_add_0_86 ),
	.shareout(Xd_0__inst_inst_add_0_87 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_89 (
// Equation(s):
// Xd_0__inst_inst_add_0_89_sumout  = SUM(( !Xd_0__inst_r_sum1_2__22__q  $ (!Xd_0__inst_r_sum1_1__22__q  $ (Xd_0__inst_r_sum1_0__22__q )) ) + ( Xd_0__inst_inst_add_0_87  ) + ( Xd_0__inst_inst_add_0_86  ))
// Xd_0__inst_inst_add_0_90  = CARRY(( !Xd_0__inst_r_sum1_2__22__q  $ (!Xd_0__inst_r_sum1_1__22__q  $ (Xd_0__inst_r_sum1_0__22__q )) ) + ( Xd_0__inst_inst_add_0_87  ) + ( Xd_0__inst_inst_add_0_86  ))
// Xd_0__inst_inst_add_0_91  = SHARE((!Xd_0__inst_r_sum1_2__22__q  & (Xd_0__inst_r_sum1_1__22__q  & Xd_0__inst_r_sum1_0__22__q )) # (Xd_0__inst_r_sum1_2__22__q  & ((Xd_0__inst_r_sum1_0__22__q ) # (Xd_0__inst_r_sum1_1__22__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__22__q ),
	.datac(!Xd_0__inst_r_sum1_1__22__q ),
	.datad(!Xd_0__inst_r_sum1_0__22__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_86 ),
	.sharein(Xd_0__inst_inst_add_0_87 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_89_sumout ),
	.cout(Xd_0__inst_inst_add_0_90 ),
	.shareout(Xd_0__inst_inst_add_0_91 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_93 (
// Equation(s):
// Xd_0__inst_inst_add_0_93_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_91  ) + ( Xd_0__inst_inst_add_0_90  ))
// Xd_0__inst_inst_add_0_94  = CARRY(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_91  ) + ( Xd_0__inst_inst_add_0_90  ))
// Xd_0__inst_inst_add_0_95  = SHARE((!Xd_0__inst_r_sum1_2__23__q  & (Xd_0__inst_r_sum1_1__23__q  & Xd_0__inst_r_sum1_0__23__q )) # (Xd_0__inst_r_sum1_2__23__q  & ((Xd_0__inst_r_sum1_0__23__q ) # (Xd_0__inst_r_sum1_1__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_90 ),
	.sharein(Xd_0__inst_inst_add_0_91 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_93_sumout ),
	.cout(Xd_0__inst_inst_add_0_94 ),
	.shareout(Xd_0__inst_inst_add_0_95 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000033F00003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_97 (
// Equation(s):
// Xd_0__inst_inst_add_0_97_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_95  ) + ( Xd_0__inst_inst_add_0_94  ))
// Xd_0__inst_inst_add_0_98  = CARRY(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_95  ) + ( Xd_0__inst_inst_add_0_94  ))
// Xd_0__inst_inst_add_0_99  = SHARE((!Xd_0__inst_r_sum1_2__23__q  & (Xd_0__inst_r_sum1_1__23__q  & Xd_0__inst_r_sum1_0__23__q )) # (Xd_0__inst_r_sum1_2__23__q  & ((Xd_0__inst_r_sum1_0__23__q ) # (Xd_0__inst_r_sum1_1__23__q ))))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_94 ),
	.sharein(Xd_0__inst_inst_add_0_95 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_97_sumout ),
	.cout(Xd_0__inst_inst_add_0_98 ),
	.shareout(Xd_0__inst_inst_add_0_99 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000003CC3),
	.shared_arith("on")
) Xd_0__inst_inst_add_0_101 (
// Equation(s):
// Xd_0__inst_inst_add_0_101_sumout  = SUM(( !Xd_0__inst_r_sum1_2__23__q  $ (!Xd_0__inst_r_sum1_1__23__q  $ (Xd_0__inst_r_sum1_0__23__q )) ) + ( Xd_0__inst_inst_add_0_99  ) + ( Xd_0__inst_inst_add_0_98  ))

	.dataa(gnd),
	.datab(!Xd_0__inst_r_sum1_2__23__q ),
	.datac(!Xd_0__inst_r_sum1_1__23__q ),
	.datad(!Xd_0__inst_r_sum1_0__23__q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_inst_add_0_98 ),
	.sharein(Xd_0__inst_inst_add_0_99 ),
	.combout(),
	.sumout(Xd_0__inst_inst_add_0_101_sumout ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_66 (
// Equation(s):
// Xd_0__inst_mult_1_176  = SUM(( (!din_a[13] & (((din_a[14] & din_b[12])))) # (din_a[13] & (!din_b[13] $ (((!din_a[14]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_182  ) + ( Xd_0__inst_mult_1_181  ))
// Xd_0__inst_mult_1_177  = CARRY(( (!din_a[13] & (((din_a[14] & din_b[12])))) # (din_a[13] & (!din_b[13] $ (((!din_a[14]) # (!din_b[12]))))) ) + ( Xd_0__inst_mult_1_182  ) + ( Xd_0__inst_mult_1_181  ))
// Xd_0__inst_mult_1_178  = SHARE((din_a[13] & (din_b[13] & (din_a[14] & din_b[12]))))

	.dataa(!din_a[13]),
	.datab(!din_b[13]),
	.datac(!din_a[14]),
	.datad(!din_b[12]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_181 ),
	.sharein(Xd_0__inst_mult_1_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_176 ),
	.cout(Xd_0__inst_mult_1_177 ),
	.shareout(Xd_0__inst_mult_1_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_168 (
// Equation(s):
// Xd_0__inst_mult_3_169  = SUM(( GND ) + ( Xd_0__inst_mult_3_175  ) + ( Xd_0__inst_mult_3_174  ))
// Xd_0__inst_mult_3_170  = CARRY(( GND ) + ( Xd_0__inst_mult_3_175  ) + ( Xd_0__inst_mult_3_174  ))
// Xd_0__inst_mult_3_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_174 ),
	.sharein(Xd_0__inst_mult_3_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_169 ),
	.cout(Xd_0__inst_mult_3_170 ),
	.shareout(Xd_0__inst_mult_3_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( Xd_0__inst_mult_7_175  ) + ( Xd_0__inst_mult_7_174  ))
// Xd_0__inst_a1_3__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_6__0__q  $ (!Xd_0__inst_product_7__0__q ) ) + ( Xd_0__inst_mult_7_175  ) + ( Xd_0__inst_mult_7_174  ))
// Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & ((Xd_0__inst_sign [6]))) # (Xd_0__inst_sign [7] & (!Xd_0__inst_product_7__0__q )))) # (Xd_0__inst_product_6__0__q  & ((!Xd_0__inst_sign [7] & 
// (Xd_0__inst_product_7__0__q )) # (Xd_0__inst_sign [7] & ((!Xd_0__inst_sign [6]))))))

	.dataa(!Xd_0__inst_product_6__0__q ),
	.datab(!Xd_0__inst_product_7__0__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_174 ),
	.sharein(Xd_0__inst_mult_7_175 ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_6__1__q  $ (!Xd_0__inst_product_7__1__q  $ (((Xd_0__inst_sign [7]) # (Xd_0__inst_sign [6])))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [6] & (Xd_0__inst_product_6__1__q  & (!Xd_0__inst_product_7__1__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_sign [6] & ((!Xd_0__inst_product_7__1__q  & ((Xd_0__inst_sign [7]))) # 
// (Xd_0__inst_product_7__1__q  & (!Xd_0__inst_product_6__1__q )))))

	.dataa(!Xd_0__inst_product_6__1__q ),
	.datab(!Xd_0__inst_product_7__1__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_6__2__q  $ (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__2__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__2__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__2__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__2__q ),
	.datab(!Xd_0__inst_product_7__2__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_6__3__q  $ (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__3__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__3__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__3__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__3__q ),
	.datab(!Xd_0__inst_product_7__3__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_6__4__q  $ (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__4__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__4__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__4__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__4__q ),
	.datab(!Xd_0__inst_product_7__4__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_6__5__q  $ (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__5__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__5__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__5__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__5__q ),
	.datab(!Xd_0__inst_product_7__5__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_6__6__q  $ (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__6__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__6__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__6__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__6__q ),
	.datab(!Xd_0__inst_product_7__6__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_6__7__q  $ (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__7__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__7__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__7__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__7__q ),
	.datab(!Xd_0__inst_product_7__7__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_6__8__q  $ (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__8__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__8__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__8__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__8__q ),
	.datab(!Xd_0__inst_product_7__8__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_6__9__q  $ (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__9__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__9__q  & (!Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__9__q 
//  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__9__q ),
	.datab(!Xd_0__inst_product_7__9__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_6__10__q  $ (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__10__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__10__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__10__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__10__q ),
	.datab(!Xd_0__inst_product_7__10__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_6__11__q  $ (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__11__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__11__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__11__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__11__q ),
	.datab(!Xd_0__inst_product_7__11__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_6__12__q  $ (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_6__12__q  $ (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__12__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__12__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__12__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__12__q ),
	.datab(!Xd_0__inst_product_7__12__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_6__13__q  $ (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_6__13__q  $ (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__13__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__13__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__13__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__13__q ),
	.datab(!Xd_0__inst_product_7__13__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_6__14__q  $ (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_6__14__q  $ (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__14__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__14__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__14__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__14__q ),
	.datab(!Xd_0__inst_product_7__14__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_6__15__q  $ (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_6__15__q  $ (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__15__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__15__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__15__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__15__q ),
	.datab(!Xd_0__inst_product_7__15__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_6__16__q  $ (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_6__16__q  $ (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__16__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__16__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__16__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__16__q ),
	.datab(!Xd_0__inst_product_7__16__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_6__17__q  $ (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_6__17__q  $ (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__17__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__17__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__17__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__17__q ),
	.datab(!Xd_0__inst_product_7__17__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_6__18__q  $ (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_6__18__q  $ (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__18__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__18__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__18__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__18__q ),
	.datab(!Xd_0__inst_product_7__18__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_6__19__q  $ (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_6__19__q  $ (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__19__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__19__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__19__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__19__q ),
	.datab(!Xd_0__inst_product_7__19__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_6__20__q  $ (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_6__20__q  $ (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__20__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__20__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__20__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__20__q ),
	.datab(!Xd_0__inst_product_7__20__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_6__21__q  $ (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_6__21__q  $ (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]))) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_6__21__q  & (Xd_0__inst_sign [6] & (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [7])))) # (Xd_0__inst_product_6__21__q  & (!Xd_0__inst_sign [6] & 
// (!Xd_0__inst_product_7__21__q  $ (!Xd_0__inst_sign [7])))))

	.dataa(!Xd_0__inst_product_6__21__q ),
	.datab(!Xd_0__inst_product_7__21__q ),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [6] & Xd_0__inst_sign [7]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_3__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_3__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [6] $ (!Xd_0__inst_sign [7]) ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_3__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [6]),
	.datad(!Xd_0__inst_sign [7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_3__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_3__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_3__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_67 (
// Equation(s):
// Xd_0__inst_mult_1_180  = SUM(( (din_a[13] & din_b[12]) ) + ( Xd_0__inst_mult_1_186  ) + ( Xd_0__inst_mult_1_185  ))
// Xd_0__inst_mult_1_181  = CARRY(( (din_a[13] & din_b[12]) ) + ( Xd_0__inst_mult_1_186  ) + ( Xd_0__inst_mult_1_185  ))
// Xd_0__inst_mult_1_182  = SHARE((din_a[12] & din_b[14]))

	.dataa(!din_a[13]),
	.datab(!din_b[12]),
	.datac(!din_a[12]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_185 ),
	.sharein(Xd_0__inst_mult_1_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_180 ),
	.cout(Xd_0__inst_mult_1_181 ),
	.shareout(Xd_0__inst_mult_1_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( Xd_0__inst_mult_3_178  ) + ( Xd_0__inst_mult_3_177  ))
// Xd_0__inst_a1_2__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_4__0__q  $ (!Xd_0__inst_product_5__0__q ) ) + ( Xd_0__inst_mult_3_178  ) + ( Xd_0__inst_mult_3_177  ))
// Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & ((Xd_0__inst_sign [4]))) # (Xd_0__inst_sign [5] & (!Xd_0__inst_product_5__0__q )))) # (Xd_0__inst_product_4__0__q  & ((!Xd_0__inst_sign [5] & 
// (Xd_0__inst_product_5__0__q )) # (Xd_0__inst_sign [5] & ((!Xd_0__inst_sign [4]))))))

	.dataa(!Xd_0__inst_product_4__0__q ),
	.datab(!Xd_0__inst_product_5__0__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_177 ),
	.sharein(Xd_0__inst_mult_3_178 ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_mult_6_175  ) + ( Xd_0__inst_mult_6_174  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_2__0__q  $ (!Xd_0__inst_product_3__0__q ) ) + ( Xd_0__inst_mult_6_175  ) + ( Xd_0__inst_mult_6_174  ))
// Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & ((Xd_0__inst_sign [2]))) # (Xd_0__inst_sign [3] & (!Xd_0__inst_product_3__0__q )))) # (Xd_0__inst_product_2__0__q  & ((!Xd_0__inst_sign [3] & 
// (Xd_0__inst_product_3__0__q )) # (Xd_0__inst_sign [3] & ((!Xd_0__inst_sign [2]))))))

	.dataa(!Xd_0__inst_product_2__0__q ),
	.datab(!Xd_0__inst_product_3__0__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_174 ),
	.sharein(Xd_0__inst_mult_6_175 ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h00001BD800006666),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc0 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [0] = SUM(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_mult_0_171  ) + ( Xd_0__inst_mult_0_170  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_COUT  = CARRY(( !Xd_0__inst_product_0__0__q  $ (!Xd_0__inst_product_1__0__q ) ) + ( Xd_0__inst_mult_0_171  ) + ( Xd_0__inst_mult_0_170  ))
// Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  = SHARE((!Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & ((Xd_0__inst_sign [0]))) # (Xd_0__inst_sign [1] & (!Xd_0__inst_product_1__0__q )))) # (Xd_0__inst_product_0__0__q  & ((!Xd_0__inst_sign [1] & 
// (Xd_0__inst_product_1__0__q )) # (Xd_0__inst_sign [1] & ((!Xd_0__inst_sign [0]))))))

	.dataa(!Xd_0__inst_product_0__0__q ),
	.datab(!Xd_0__inst_product_1__0__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_170 ),
	.sharein(Xd_0__inst_mult_0_171 ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3 (
// Equation(s):
// Xd_0__inst_mult_3_173  = SUM(( (din_a[44] & din_b[46]) ) + ( Xd_0__inst_mult_3_182  ) + ( Xd_0__inst_mult_3_181  ))
// Xd_0__inst_mult_3_174  = CARRY(( (din_a[44] & din_b[46]) ) + ( Xd_0__inst_mult_3_182  ) + ( Xd_0__inst_mult_3_181  ))
// Xd_0__inst_mult_3_175  = SHARE(GND)

	.dataa(!din_a[44]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_181 ),
	.sharein(Xd_0__inst_mult_3_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_173 ),
	.cout(Xd_0__inst_mult_3_174 ),
	.shareout(Xd_0__inst_mult_3_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_172 (
// Equation(s):
// Xd_0__inst_mult_7_173  = SUM(( GND ) + ( Xd_0__inst_mult_7_179  ) + ( Xd_0__inst_mult_7_178  ))
// Xd_0__inst_mult_7_174  = CARRY(( GND ) + ( Xd_0__inst_mult_7_179  ) + ( Xd_0__inst_mult_7_178  ))
// Xd_0__inst_mult_7_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_178 ),
	.sharein(Xd_0__inst_mult_7_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_173 ),
	.cout(Xd_0__inst_mult_7_174 ),
	.shareout(Xd_0__inst_mult_7_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_4__1__q  $ (!Xd_0__inst_product_5__1__q  $ (((Xd_0__inst_sign [5]) # (Xd_0__inst_sign [4])))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [4] & (Xd_0__inst_product_4__1__q  & (!Xd_0__inst_product_5__1__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_sign [4] & ((!Xd_0__inst_product_5__1__q  & ((Xd_0__inst_sign [5]))) # 
// (Xd_0__inst_product_5__1__q  & (!Xd_0__inst_product_4__1__q )))))

	.dataa(!Xd_0__inst_product_4__1__q ),
	.datab(!Xd_0__inst_product_5__1__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_2__1__q  $ (!Xd_0__inst_product_3__1__q  $ (((Xd_0__inst_sign [3]) # (Xd_0__inst_sign [2])))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [2] & (Xd_0__inst_product_2__1__q  & (!Xd_0__inst_product_3__1__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_sign [2] & ((!Xd_0__inst_product_3__1__q  & ((Xd_0__inst_sign [3]))) # 
// (Xd_0__inst_product_3__1__q  & (!Xd_0__inst_product_2__1__q )))))

	.dataa(!Xd_0__inst_product_2__1__q ),
	.datab(!Xd_0__inst_product_3__1__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124E00006999),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [1] = SUM(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT  
// ))
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  = CARRY(( !Xd_0__inst_product_0__1__q  $ (!Xd_0__inst_product_1__1__q  $ (((Xd_0__inst_sign [1]) # (Xd_0__inst_sign [0])))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc0_COUT 
//  ))
// Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  = SHARE((!Xd_0__inst_sign [0] & (Xd_0__inst_product_0__1__q  & (!Xd_0__inst_product_1__1__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_sign [0] & ((!Xd_0__inst_product_1__1__q  & ((Xd_0__inst_sign [1]))) # 
// (Xd_0__inst_product_1__1__q  & (!Xd_0__inst_product_0__1__q )))))

	.dataa(!Xd_0__inst_product_0__1__q ),
	.datab(!Xd_0__inst_product_1__1__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc0_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc0_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_4__2__q  $ (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__2__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__2__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__2__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__2__q ),
	.datab(!Xd_0__inst_product_5__2__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_2__2__q  $ (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__2__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__2__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__2__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__2__q ),
	.datab(!Xd_0__inst_product_3__2__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_2__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [2] = SUM(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  = CARRY(( !Xd_0__inst_product_0__2__q  $ (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_wc1_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__2__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__2__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__2__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__2__q ),
	.datab(!Xd_0__inst_product_1__2__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc1_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc1_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_4__3__q  $ (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__3__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__3__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__3__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__3__q ),
	.datab(!Xd_0__inst_product_5__3__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_2__3__q  $ (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__3__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__3__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__3__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__3__q ),
	.datab(!Xd_0__inst_product_3__3__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_3__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [3] = SUM(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  = CARRY(( !Xd_0__inst_product_0__3__q  $ (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__3__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__3__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__3__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__3__q ),
	.datab(!Xd_0__inst_product_1__3__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_2__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_4__4__q  $ (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__4__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__4__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__4__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__4__q ),
	.datab(!Xd_0__inst_product_5__4__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_2__4__q  $ (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__4__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__4__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__4__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__4__q ),
	.datab(!Xd_0__inst_product_3__4__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_4__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [4] = SUM(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  = CARRY(( !Xd_0__inst_product_0__4__q  $ (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__4__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__4__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__4__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__4__q ),
	.datab(!Xd_0__inst_product_1__4__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_3__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_4__5__q  $ (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__5__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__5__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__5__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__5__q ),
	.datab(!Xd_0__inst_product_5__5__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_2__5__q  $ (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__5__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__5__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__5__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__5__q ),
	.datab(!Xd_0__inst_product_3__5__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_5__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [5] = SUM(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  = CARRY(( !Xd_0__inst_product_0__5__q  $ (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__5__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__5__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__5__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__5__q ),
	.datab(!Xd_0__inst_product_1__5__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_4__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_4__6__q  $ (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__6__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__6__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__6__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__6__q ),
	.datab(!Xd_0__inst_product_5__6__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_2__6__q  $ (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__6__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__6__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__6__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__6__q ),
	.datab(!Xd_0__inst_product_3__6__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_6__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [6] = SUM(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  = CARRY(( !Xd_0__inst_product_0__6__q  $ (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__6__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__6__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__6__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__6__q ),
	.datab(!Xd_0__inst_product_1__6__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_5__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_4__7__q  $ (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__7__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__7__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__7__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__7__q ),
	.datab(!Xd_0__inst_product_5__7__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_2__7__q  $ (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__7__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__7__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__7__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__7__q ),
	.datab(!Xd_0__inst_product_3__7__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_7__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [7] = SUM(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  = CARRY(( !Xd_0__inst_product_0__7__q  $ (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__7__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__7__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__7__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__7__q ),
	.datab(!Xd_0__inst_product_1__7__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_6__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_4__8__q  $ (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__8__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__8__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__8__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__8__q ),
	.datab(!Xd_0__inst_product_5__8__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_2__8__q  $ (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__8__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__8__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__8__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__8__q ),
	.datab(!Xd_0__inst_product_3__8__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_8__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [8] = SUM(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  = CARRY(( !Xd_0__inst_product_0__8__q  $ (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__8__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__8__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__8__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__8__q ),
	.datab(!Xd_0__inst_product_1__8__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_7__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_4__9__q  $ (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__9__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__9__q  & (!Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__9__q 
//  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__9__q ),
	.datab(!Xd_0__inst_product_5__9__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_2__9__q  $ (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__9__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__9__q  & (!Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__9__q 
//  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__9__q ),
	.datab(!Xd_0__inst_product_3__9__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_9__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [9] = SUM(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  = CARRY(( !Xd_0__inst_product_0__9__q  $ (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__9__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__9__q  & (!Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__9__q 
//  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__9__q ),
	.datab(!Xd_0__inst_product_1__9__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_8__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_4__10__q  $ (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__10__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__10__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__10__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__10__q ),
	.datab(!Xd_0__inst_product_5__10__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_2__10__q  $ (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__10__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__10__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__10__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__10__q ),
	.datab(!Xd_0__inst_product_3__10__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_10__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [10] = SUM(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  = CARRY(( !Xd_0__inst_product_0__10__q  $ (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__10__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__10__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__10__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__10__q ),
	.datab(!Xd_0__inst_product_1__10__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_9__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_4__11__q  $ (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__11__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__11__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__11__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__11__q ),
	.datab(!Xd_0__inst_product_5__11__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_2__11__q  $ (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__11__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__11__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__11__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__11__q ),
	.datab(!Xd_0__inst_product_3__11__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_11__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [11] = SUM(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  = CARRY(( !Xd_0__inst_product_0__11__q  $ (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__11__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__11__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__11__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__11__q ),
	.datab(!Xd_0__inst_product_1__11__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_10__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_4__12__q  $ (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_4__12__q  $ (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__12__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__12__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__12__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__12__q ),
	.datab(!Xd_0__inst_product_5__12__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_2__12__q  $ (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_2__12__q  $ (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__12__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__12__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__12__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__12__q ),
	.datab(!Xd_0__inst_product_3__12__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_12__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [12] = SUM(( !Xd_0__inst_product_0__12__q  $ (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  = CARRY(( !Xd_0__inst_product_0__12__q  $ (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__12__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__12__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__12__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__12__q ),
	.datab(!Xd_0__inst_product_1__12__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_11__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_4__13__q  $ (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_4__13__q  $ (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__13__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__13__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__13__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__13__q ),
	.datab(!Xd_0__inst_product_5__13__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_2__13__q  $ (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_2__13__q  $ (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__13__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__13__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__13__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__13__q ),
	.datab(!Xd_0__inst_product_3__13__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_13__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [13] = SUM(( !Xd_0__inst_product_0__13__q  $ (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  = CARRY(( !Xd_0__inst_product_0__13__q  $ (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__13__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__13__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__13__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__13__q ),
	.datab(!Xd_0__inst_product_1__13__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_12__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_4__14__q  $ (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_4__14__q  $ (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__14__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__14__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__14__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__14__q ),
	.datab(!Xd_0__inst_product_5__14__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_2__14__q  $ (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_2__14__q  $ (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__14__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__14__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__14__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__14__q ),
	.datab(!Xd_0__inst_product_3__14__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_14__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [14] = SUM(( !Xd_0__inst_product_0__14__q  $ (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  = CARRY(( !Xd_0__inst_product_0__14__q  $ (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__14__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__14__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__14__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__14__q ),
	.datab(!Xd_0__inst_product_1__14__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_13__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [14]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_4__15__q  $ (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_4__15__q  $ (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__15__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__15__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__15__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__15__q ),
	.datab(!Xd_0__inst_product_5__15__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_2__15__q  $ (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_2__15__q  $ (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__15__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__15__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__15__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__15__q ),
	.datab(!Xd_0__inst_product_3__15__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_15__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [15] = SUM(( !Xd_0__inst_product_0__15__q  $ (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  = CARRY(( !Xd_0__inst_product_0__15__q  $ (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__15__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__15__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__15__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__15__q ),
	.datab(!Xd_0__inst_product_1__15__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_14__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [15]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_4__16__q  $ (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_4__16__q  $ (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__16__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__16__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__16__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__16__q ),
	.datab(!Xd_0__inst_product_5__16__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_2__16__q  $ (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_2__16__q  $ (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__16__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__16__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__16__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__16__q ),
	.datab(!Xd_0__inst_product_3__16__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_16__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [16] = SUM(( !Xd_0__inst_product_0__16__q  $ (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  = CARRY(( !Xd_0__inst_product_0__16__q  $ (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__16__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__16__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__16__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__16__q ),
	.datab(!Xd_0__inst_product_1__16__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_15__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [16]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_4__17__q  $ (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_4__17__q  $ (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__17__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__17__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__17__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__17__q ),
	.datab(!Xd_0__inst_product_5__17__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_2__17__q  $ (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_2__17__q  $ (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__17__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__17__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__17__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__17__q ),
	.datab(!Xd_0__inst_product_3__17__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_17__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [17] = SUM(( !Xd_0__inst_product_0__17__q  $ (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  = CARRY(( !Xd_0__inst_product_0__17__q  $ (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__17__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__17__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__17__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__17__q ),
	.datab(!Xd_0__inst_product_1__17__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_16__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [17]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_4__18__q  $ (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_4__18__q  $ (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__18__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__18__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__18__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__18__q ),
	.datab(!Xd_0__inst_product_5__18__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_2__18__q  $ (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_2__18__q  $ (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__18__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__18__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__18__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__18__q ),
	.datab(!Xd_0__inst_product_3__18__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_18__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [18] = SUM(( !Xd_0__inst_product_0__18__q  $ (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  = CARRY(( !Xd_0__inst_product_0__18__q  $ (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__18__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__18__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__18__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__18__q ),
	.datab(!Xd_0__inst_product_1__18__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_17__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [18]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_4__19__q  $ (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_4__19__q  $ (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__19__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__19__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__19__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__19__q ),
	.datab(!Xd_0__inst_product_5__19__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_2__19__q  $ (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_2__19__q  $ (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__19__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__19__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__19__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__19__q ),
	.datab(!Xd_0__inst_product_3__19__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_19__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [19] = SUM(( !Xd_0__inst_product_0__19__q  $ (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  = CARRY(( !Xd_0__inst_product_0__19__q  $ (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__19__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__19__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__19__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__19__q ),
	.datab(!Xd_0__inst_product_1__19__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_18__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [19]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_4__20__q  $ (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_4__20__q  $ (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__20__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__20__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__20__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__20__q ),
	.datab(!Xd_0__inst_product_5__20__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_2__20__q  $ (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_2__20__q  $ (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__20__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__20__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__20__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__20__q ),
	.datab(!Xd_0__inst_product_3__20__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_20__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [20] = SUM(( !Xd_0__inst_product_0__20__q  $ (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  = CARRY(( !Xd_0__inst_product_0__20__q  $ (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__20__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__20__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__20__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__20__q ),
	.datab(!Xd_0__inst_product_1__20__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_19__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [20]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_4__21__q  $ (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_4__21__q  $ (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]))) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_4__21__q  & (Xd_0__inst_sign [4] & (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [5])))) # (Xd_0__inst_product_4__21__q  & (!Xd_0__inst_sign [4] & 
// (!Xd_0__inst_product_5__21__q  $ (!Xd_0__inst_sign [5])))))

	.dataa(!Xd_0__inst_product_4__21__q ),
	.datab(!Xd_0__inst_product_5__21__q ),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_2__21__q  $ (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_2__21__q  $ (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]))) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_2__21__q  & (Xd_0__inst_sign [2] & (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [3])))) # (Xd_0__inst_product_2__21__q  & (!Xd_0__inst_sign [2] & 
// (!Xd_0__inst_product_3__21__q  $ (!Xd_0__inst_sign [3])))))

	.dataa(!Xd_0__inst_product_2__21__q ),
	.datab(!Xd_0__inst_product_3__21__q ),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000124800006996),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_gen_21__wc (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [21] = SUM(( !Xd_0__inst_product_0__21__q  $ (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  = CARRY(( !Xd_0__inst_product_0__21__q  $ (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]))) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT  ) + ( 
// Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  = SHARE((!Xd_0__inst_product_0__21__q  & (Xd_0__inst_sign [0] & (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [1])))) # (Xd_0__inst_product_0__21__q  & (!Xd_0__inst_sign [0] & 
// (!Xd_0__inst_product_1__21__q  $ (!Xd_0__inst_sign [1])))))

	.dataa(!Xd_0__inst_product_0__21__q ),
	.datab(!Xd_0__inst_product_1__21__q ),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_20__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [21]),
	.cout(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [4] & Xd_0__inst_sign [5]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [2] & Xd_0__inst_sign [3]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [22] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  = CARRY(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT  ))
// Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  = SHARE((Xd_0__inst_sign [0] & Xd_0__inst_sign [1]))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_gen_21__wc_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [22]),
	.cout(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.shareout(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_2__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_2__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [4] $ (!Xd_0__inst_sign [5]) ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_2__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [4]),
	.datad(!Xd_0__inst_sign [5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_2__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_2__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_2__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_1__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_1__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [2] $ (!Xd_0__inst_sign [3]) ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_1__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [2]),
	.datad(!Xd_0__inst_sign [3]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_1__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_1__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_1__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000FF0),
	.shared_arith("on")
) Xd_0__inst_a1_0__adder1_inst_wc_n_plus_1 (
// Equation(s):
// Xd_0__inst_a1_0__adder1_inst_dout [23] = SUM(( !Xd_0__inst_sign [0] $ (!Xd_0__inst_sign [1]) ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT  ) + ( Xd_0__inst_a1_0__adder1_inst_wc_n_COUT  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(!Xd_0__inst_sign [0]),
	.datad(!Xd_0__inst_sign [1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_a1_0__adder1_inst_wc_n_COUT ),
	.sharein(Xd_0__inst_a1_0__adder1_inst_wc_n_SHAREOUT ),
	.combout(),
	.sumout(Xd_0__inst_a1_0__adder1_inst_dout [23]),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_68 (
// Equation(s):
// Xd_0__inst_mult_1_184  = SUM(( (din_a[12] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_185  = CARRY(( (din_a[12] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_186  = SHARE((din_a[12] & din_b[13]))

	.dataa(!din_a[12]),
	.datab(!din_b[12]),
	.datac(!din_b[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_184 ),
	.cout(Xd_0__inst_mult_1_185 ),
	.shareout(Xd_0__inst_mult_1_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_66 (
// Equation(s):
// Xd_0__inst_mult_3_176  = SUM(( GND ) + ( Xd_0__inst_mult_3_186  ) + ( Xd_0__inst_mult_3_185  ))
// Xd_0__inst_mult_3_177  = CARRY(( GND ) + ( Xd_0__inst_mult_3_186  ) + ( Xd_0__inst_mult_3_185  ))
// Xd_0__inst_mult_3_178  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_185 ),
	.sharein(Xd_0__inst_mult_3_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_176 ),
	.cout(Xd_0__inst_mult_3_177 ),
	.shareout(Xd_0__inst_mult_3_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_172 (
// Equation(s):
// Xd_0__inst_mult_6_173  = SUM(( GND ) + ( Xd_0__inst_mult_6_246  ) + ( Xd_0__inst_mult_6_245  ))
// Xd_0__inst_mult_6_174  = CARRY(( GND ) + ( Xd_0__inst_mult_6_246  ) + ( Xd_0__inst_mult_6_245  ))
// Xd_0__inst_mult_6_175  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_245 ),
	.sharein(Xd_0__inst_mult_6_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_173 ),
	.cout(Xd_0__inst_mult_6_174 ),
	.shareout(Xd_0__inst_mult_6_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_168 (
// Equation(s):
// Xd_0__inst_mult_0_169  = SUM(( GND ) + ( Xd_0__inst_mult_0_175  ) + ( Xd_0__inst_mult_0_174  ))
// Xd_0__inst_mult_0_170  = CARRY(( GND ) + ( Xd_0__inst_mult_0_175  ) + ( Xd_0__inst_mult_0_174  ))
// Xd_0__inst_mult_0_171  = SHARE(GND)

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_174 ),
	.sharein(Xd_0__inst_mult_0_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_169 ),
	.cout(Xd_0__inst_mult_0_170 ),
	.shareout(Xd_0__inst_mult_0_171 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_67 (
// Equation(s):
// Xd_0__inst_mult_3_180  = SUM(( (!din_a[44] & (((din_a[43] & din_b[46])))) # (din_a[44] & (!din_b[45] $ (((!din_a[43]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_190  ) + ( Xd_0__inst_mult_3_189  ))
// Xd_0__inst_mult_3_181  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[46])))) # (din_a[44] & (!din_b[45] $ (((!din_a[43]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_190  ) + ( Xd_0__inst_mult_3_189  ))
// Xd_0__inst_mult_3_182  = SHARE((din_a[44] & (din_b[45] & (din_a[43] & din_b[46]))))

	.dataa(!din_a[44]),
	.datab(!din_b[45]),
	.datac(!din_a[43]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_189 ),
	.sharein(Xd_0__inst_mult_3_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_180 ),
	.cout(Xd_0__inst_mult_3_181 ),
	.shareout(Xd_0__inst_mult_3_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7 (
// Equation(s):
// Xd_0__inst_mult_7_177  = SUM(( !Xd_0__inst_mult_7_252  $ (((!din_b[88]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_258  ) + ( Xd_0__inst_mult_7_257  ))
// Xd_0__inst_mult_7_178  = CARRY(( !Xd_0__inst_mult_7_252  $ (((!din_b[88]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_258  ) + ( Xd_0__inst_mult_7_257  ))
// Xd_0__inst_mult_7_179  = SHARE((din_b[88] & (din_a[94] & Xd_0__inst_mult_7_252 )))

	.dataa(!din_b[88]),
	.datab(!din_a[94]),
	.datac(!Xd_0__inst_mult_7_252 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_257 ),
	.sharein(Xd_0__inst_mult_7_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_177 ),
	.cout(Xd_0__inst_mult_7_178 ),
	.shareout(Xd_0__inst_mult_7_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6 (
// Equation(s):
// Xd_0__inst_mult_6_177  = SUM(( !Xd_0__inst_mult_6_0_q  $ (!Xd_0__inst_mult_6_1_q ) ) + ( Xd_0__inst_mult_4_37  ) + ( Xd_0__inst_mult_4_36  ))
// Xd_0__inst_mult_6_178  = CARRY(( !Xd_0__inst_mult_6_0_q  $ (!Xd_0__inst_mult_6_1_q ) ) + ( Xd_0__inst_mult_4_37  ) + ( Xd_0__inst_mult_4_36  ))
// Xd_0__inst_mult_6_179  = SHARE((Xd_0__inst_mult_6_0_q  & Xd_0__inst_mult_6_1_q ))

	.dataa(!Xd_0__inst_mult_6_0_q ),
	.datab(!Xd_0__inst_mult_6_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_36 ),
	.sharein(Xd_0__inst_mult_4_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_177 ),
	.cout(Xd_0__inst_mult_6_178 ),
	.shareout(Xd_0__inst_mult_6_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_70 (
// Equation(s):
// Xd_0__inst_mult_7_180  = SUM(( !Xd_0__inst_mult_7_0_q  $ (!Xd_0__inst_mult_7_1_q ) ) + ( Xd_0__inst_mult_3_37  ) + ( Xd_0__inst_mult_3_36  ))
// Xd_0__inst_mult_7_181  = CARRY(( !Xd_0__inst_mult_7_0_q  $ (!Xd_0__inst_mult_7_1_q ) ) + ( Xd_0__inst_mult_3_37  ) + ( Xd_0__inst_mult_3_36  ))
// Xd_0__inst_mult_7_182  = SHARE((Xd_0__inst_mult_7_0_q  & Xd_0__inst_mult_7_1_q ))

	.dataa(!Xd_0__inst_mult_7_0_q ),
	.datab(!Xd_0__inst_mult_7_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_36 ),
	.sharein(Xd_0__inst_mult_3_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_180 ),
	.cout(Xd_0__inst_mult_7_181 ),
	.shareout(Xd_0__inst_mult_7_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_70 (
// Equation(s):
// Xd_0__inst_mult_6_180  = SUM(( !Xd_0__inst_mult_6_2_q  $ (!Xd_0__inst_mult_6_3_q ) ) + ( Xd_0__inst_mult_6_179  ) + ( Xd_0__inst_mult_6_178  ))
// Xd_0__inst_mult_6_181  = CARRY(( !Xd_0__inst_mult_6_2_q  $ (!Xd_0__inst_mult_6_3_q ) ) + ( Xd_0__inst_mult_6_179  ) + ( Xd_0__inst_mult_6_178  ))
// Xd_0__inst_mult_6_182  = SHARE((Xd_0__inst_mult_6_2_q  & Xd_0__inst_mult_6_3_q ))

	.dataa(!Xd_0__inst_mult_6_2_q ),
	.datab(!Xd_0__inst_mult_6_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_178 ),
	.sharein(Xd_0__inst_mult_6_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_180 ),
	.cout(Xd_0__inst_mult_6_181 ),
	.shareout(Xd_0__inst_mult_6_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_71 (
// Equation(s):
// Xd_0__inst_mult_7_184  = SUM(( !Xd_0__inst_mult_7_2_q  $ (!Xd_0__inst_mult_7_3_q ) ) + ( Xd_0__inst_mult_7_182  ) + ( Xd_0__inst_mult_7_181  ))
// Xd_0__inst_mult_7_185  = CARRY(( !Xd_0__inst_mult_7_2_q  $ (!Xd_0__inst_mult_7_3_q ) ) + ( Xd_0__inst_mult_7_182  ) + ( Xd_0__inst_mult_7_181  ))
// Xd_0__inst_mult_7_186  = SHARE((Xd_0__inst_mult_7_2_q  & Xd_0__inst_mult_7_3_q ))

	.dataa(!Xd_0__inst_mult_7_2_q ),
	.datab(!Xd_0__inst_mult_7_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_181 ),
	.sharein(Xd_0__inst_mult_7_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_184 ),
	.cout(Xd_0__inst_mult_7_185 ),
	.shareout(Xd_0__inst_mult_7_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_71 (
// Equation(s):
// Xd_0__inst_mult_6_184  = SUM(( !Xd_0__inst_mult_6_4_q  $ (!Xd_0__inst_mult_6_5_q ) ) + ( Xd_0__inst_mult_6_182  ) + ( Xd_0__inst_mult_6_181  ))
// Xd_0__inst_mult_6_185  = CARRY(( !Xd_0__inst_mult_6_4_q  $ (!Xd_0__inst_mult_6_5_q ) ) + ( Xd_0__inst_mult_6_182  ) + ( Xd_0__inst_mult_6_181  ))
// Xd_0__inst_mult_6_186  = SHARE((Xd_0__inst_mult_6_4_q  & Xd_0__inst_mult_6_5_q ))

	.dataa(!Xd_0__inst_mult_6_4_q ),
	.datab(!Xd_0__inst_mult_6_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_181 ),
	.sharein(Xd_0__inst_mult_6_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_184 ),
	.cout(Xd_0__inst_mult_6_185 ),
	.shareout(Xd_0__inst_mult_6_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_72 (
// Equation(s):
// Xd_0__inst_mult_7_188  = SUM(( !Xd_0__inst_mult_7_4_q  $ (!Xd_0__inst_mult_7_5_q ) ) + ( Xd_0__inst_mult_7_186  ) + ( Xd_0__inst_mult_7_185  ))
// Xd_0__inst_mult_7_189  = CARRY(( !Xd_0__inst_mult_7_4_q  $ (!Xd_0__inst_mult_7_5_q ) ) + ( Xd_0__inst_mult_7_186  ) + ( Xd_0__inst_mult_7_185  ))
// Xd_0__inst_mult_7_190  = SHARE((Xd_0__inst_mult_7_4_q  & Xd_0__inst_mult_7_5_q ))

	.dataa(!Xd_0__inst_mult_7_4_q ),
	.datab(!Xd_0__inst_mult_7_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_185 ),
	.sharein(Xd_0__inst_mult_7_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_188 ),
	.cout(Xd_0__inst_mult_7_189 ),
	.shareout(Xd_0__inst_mult_7_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_72 (
// Equation(s):
// Xd_0__inst_mult_6_188  = SUM(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_186  ) + ( Xd_0__inst_mult_6_185  ))
// Xd_0__inst_mult_6_189  = CARRY(( !Xd_0__inst_mult_6_6_q  $ (!Xd_0__inst_mult_6_7_q ) ) + ( Xd_0__inst_mult_6_186  ) + ( Xd_0__inst_mult_6_185  ))
// Xd_0__inst_mult_6_190  = SHARE((Xd_0__inst_mult_6_6_q  & Xd_0__inst_mult_6_7_q ))

	.dataa(!Xd_0__inst_mult_6_6_q ),
	.datab(!Xd_0__inst_mult_6_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_185 ),
	.sharein(Xd_0__inst_mult_6_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_188 ),
	.cout(Xd_0__inst_mult_6_189 ),
	.shareout(Xd_0__inst_mult_6_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_73 (
// Equation(s):
// Xd_0__inst_mult_7_192  = SUM(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_190  ) + ( Xd_0__inst_mult_7_189  ))
// Xd_0__inst_mult_7_193  = CARRY(( !Xd_0__inst_mult_7_6_q  $ (!Xd_0__inst_mult_7_7_q ) ) + ( Xd_0__inst_mult_7_190  ) + ( Xd_0__inst_mult_7_189  ))
// Xd_0__inst_mult_7_194  = SHARE((Xd_0__inst_mult_7_6_q  & Xd_0__inst_mult_7_7_q ))

	.dataa(!Xd_0__inst_mult_7_6_q ),
	.datab(!Xd_0__inst_mult_7_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_189 ),
	.sharein(Xd_0__inst_mult_7_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_192 ),
	.cout(Xd_0__inst_mult_7_193 ),
	.shareout(Xd_0__inst_mult_7_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_73 (
// Equation(s):
// Xd_0__inst_mult_6_192  = SUM(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_190  ) + ( Xd_0__inst_mult_6_189  ))
// Xd_0__inst_mult_6_193  = CARRY(( !Xd_0__inst_mult_6_8_q  $ (!Xd_0__inst_mult_6_9_q ) ) + ( Xd_0__inst_mult_6_190  ) + ( Xd_0__inst_mult_6_189  ))
// Xd_0__inst_mult_6_194  = SHARE((Xd_0__inst_mult_6_8_q  & Xd_0__inst_mult_6_9_q ))

	.dataa(!Xd_0__inst_mult_6_8_q ),
	.datab(!Xd_0__inst_mult_6_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_189 ),
	.sharein(Xd_0__inst_mult_6_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_192 ),
	.cout(Xd_0__inst_mult_6_193 ),
	.shareout(Xd_0__inst_mult_6_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_74 (
// Equation(s):
// Xd_0__inst_mult_7_196  = SUM(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_194  ) + ( Xd_0__inst_mult_7_193  ))
// Xd_0__inst_mult_7_197  = CARRY(( !Xd_0__inst_mult_7_8_q  $ (!Xd_0__inst_mult_7_9_q ) ) + ( Xd_0__inst_mult_7_194  ) + ( Xd_0__inst_mult_7_193  ))
// Xd_0__inst_mult_7_198  = SHARE((Xd_0__inst_mult_7_8_q  & Xd_0__inst_mult_7_9_q ))

	.dataa(!Xd_0__inst_mult_7_8_q ),
	.datab(!Xd_0__inst_mult_7_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_193 ),
	.sharein(Xd_0__inst_mult_7_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_196 ),
	.cout(Xd_0__inst_mult_7_197 ),
	.shareout(Xd_0__inst_mult_7_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_74 (
// Equation(s):
// Xd_0__inst_mult_6_196  = SUM(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q ) ) + ( Xd_0__inst_mult_6_194  ) + ( Xd_0__inst_mult_6_193  ))
// Xd_0__inst_mult_6_197  = CARRY(( !Xd_0__inst_mult_6_10_q  $ (!Xd_0__inst_mult_6_11_q ) ) + ( Xd_0__inst_mult_6_194  ) + ( Xd_0__inst_mult_6_193  ))
// Xd_0__inst_mult_6_198  = SHARE((Xd_0__inst_mult_6_10_q  & Xd_0__inst_mult_6_11_q ))

	.dataa(!Xd_0__inst_mult_6_10_q ),
	.datab(!Xd_0__inst_mult_6_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_193 ),
	.sharein(Xd_0__inst_mult_6_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_196 ),
	.cout(Xd_0__inst_mult_6_197 ),
	.shareout(Xd_0__inst_mult_6_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_75 (
// Equation(s):
// Xd_0__inst_mult_7_200  = SUM(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q ) ) + ( Xd_0__inst_mult_7_198  ) + ( Xd_0__inst_mult_7_197  ))
// Xd_0__inst_mult_7_201  = CARRY(( !Xd_0__inst_mult_7_10_q  $ (!Xd_0__inst_mult_7_11_q ) ) + ( Xd_0__inst_mult_7_198  ) + ( Xd_0__inst_mult_7_197  ))
// Xd_0__inst_mult_7_202  = SHARE((Xd_0__inst_mult_7_10_q  & Xd_0__inst_mult_7_11_q ))

	.dataa(!Xd_0__inst_mult_7_10_q ),
	.datab(!Xd_0__inst_mult_7_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_197 ),
	.sharein(Xd_0__inst_mult_7_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_200 ),
	.cout(Xd_0__inst_mult_7_201 ),
	.shareout(Xd_0__inst_mult_7_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_75 (
// Equation(s):
// Xd_0__inst_mult_6_200  = SUM(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_198  ) + ( Xd_0__inst_mult_6_197  ))
// Xd_0__inst_mult_6_201  = CARRY(( !Xd_0__inst_mult_6_12_q  $ (!Xd_0__inst_mult_6_13_q ) ) + ( Xd_0__inst_mult_6_198  ) + ( Xd_0__inst_mult_6_197  ))
// Xd_0__inst_mult_6_202  = SHARE((Xd_0__inst_mult_6_12_q  & Xd_0__inst_mult_6_13_q ))

	.dataa(!Xd_0__inst_mult_6_12_q ),
	.datab(!Xd_0__inst_mult_6_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_197 ),
	.sharein(Xd_0__inst_mult_6_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_200 ),
	.cout(Xd_0__inst_mult_6_201 ),
	.shareout(Xd_0__inst_mult_6_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_76 (
// Equation(s):
// Xd_0__inst_mult_7_204  = SUM(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_202  ) + ( Xd_0__inst_mult_7_201  ))
// Xd_0__inst_mult_7_205  = CARRY(( !Xd_0__inst_mult_7_12_q  $ (!Xd_0__inst_mult_7_13_q ) ) + ( Xd_0__inst_mult_7_202  ) + ( Xd_0__inst_mult_7_201  ))
// Xd_0__inst_mult_7_206  = SHARE((Xd_0__inst_mult_7_12_q  & Xd_0__inst_mult_7_13_q ))

	.dataa(!Xd_0__inst_mult_7_12_q ),
	.datab(!Xd_0__inst_mult_7_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_201 ),
	.sharein(Xd_0__inst_mult_7_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_204 ),
	.cout(Xd_0__inst_mult_7_205 ),
	.shareout(Xd_0__inst_mult_7_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_76 (
// Equation(s):
// Xd_0__inst_mult_6_204  = SUM(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_202  ) + ( Xd_0__inst_mult_6_201  ))
// Xd_0__inst_mult_6_205  = CARRY(( !Xd_0__inst_mult_6_14_q  $ (!Xd_0__inst_mult_6_15_q ) ) + ( Xd_0__inst_mult_6_202  ) + ( Xd_0__inst_mult_6_201  ))
// Xd_0__inst_mult_6_206  = SHARE((Xd_0__inst_mult_6_14_q  & Xd_0__inst_mult_6_15_q ))

	.dataa(!Xd_0__inst_mult_6_14_q ),
	.datab(!Xd_0__inst_mult_6_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_201 ),
	.sharein(Xd_0__inst_mult_6_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_204 ),
	.cout(Xd_0__inst_mult_6_205 ),
	.shareout(Xd_0__inst_mult_6_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_77 (
// Equation(s):
// Xd_0__inst_mult_7_208  = SUM(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_206  ) + ( Xd_0__inst_mult_7_205  ))
// Xd_0__inst_mult_7_209  = CARRY(( !Xd_0__inst_mult_7_14_q  $ (!Xd_0__inst_mult_7_15_q ) ) + ( Xd_0__inst_mult_7_206  ) + ( Xd_0__inst_mult_7_205  ))
// Xd_0__inst_mult_7_210  = SHARE((Xd_0__inst_mult_7_14_q  & Xd_0__inst_mult_7_15_q ))

	.dataa(!Xd_0__inst_mult_7_14_q ),
	.datab(!Xd_0__inst_mult_7_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_205 ),
	.sharein(Xd_0__inst_mult_7_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_208 ),
	.cout(Xd_0__inst_mult_7_209 ),
	.shareout(Xd_0__inst_mult_7_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_77 (
// Equation(s):
// Xd_0__inst_mult_6_208  = SUM(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q ) ) + ( Xd_0__inst_mult_6_206  ) + ( Xd_0__inst_mult_6_205  ))
// Xd_0__inst_mult_6_209  = CARRY(( !Xd_0__inst_mult_6_16_q  $ (!Xd_0__inst_mult_6_17_q ) ) + ( Xd_0__inst_mult_6_206  ) + ( Xd_0__inst_mult_6_205  ))
// Xd_0__inst_mult_6_210  = SHARE((Xd_0__inst_mult_6_16_q  & Xd_0__inst_mult_6_17_q ))

	.dataa(!Xd_0__inst_mult_6_16_q ),
	.datab(!Xd_0__inst_mult_6_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_205 ),
	.sharein(Xd_0__inst_mult_6_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_208 ),
	.cout(Xd_0__inst_mult_6_209 ),
	.shareout(Xd_0__inst_mult_6_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_78 (
// Equation(s):
// Xd_0__inst_mult_7_212  = SUM(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q ) ) + ( Xd_0__inst_mult_7_210  ) + ( Xd_0__inst_mult_7_209  ))
// Xd_0__inst_mult_7_213  = CARRY(( !Xd_0__inst_mult_7_16_q  $ (!Xd_0__inst_mult_7_17_q ) ) + ( Xd_0__inst_mult_7_210  ) + ( Xd_0__inst_mult_7_209  ))
// Xd_0__inst_mult_7_214  = SHARE((Xd_0__inst_mult_7_16_q  & Xd_0__inst_mult_7_17_q ))

	.dataa(!Xd_0__inst_mult_7_16_q ),
	.datab(!Xd_0__inst_mult_7_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_209 ),
	.sharein(Xd_0__inst_mult_7_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_212 ),
	.cout(Xd_0__inst_mult_7_213 ),
	.shareout(Xd_0__inst_mult_7_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_78 (
// Equation(s):
// Xd_0__inst_mult_6_212  = SUM(( !Xd_0__inst_mult_6_18_q  $ (!Xd_0__inst_mult_6_19_q ) ) + ( Xd_0__inst_mult_6_210  ) + ( Xd_0__inst_mult_6_209  ))
// Xd_0__inst_mult_6_213  = CARRY(( !Xd_0__inst_mult_6_18_q  $ (!Xd_0__inst_mult_6_19_q ) ) + ( Xd_0__inst_mult_6_210  ) + ( Xd_0__inst_mult_6_209  ))
// Xd_0__inst_mult_6_214  = SHARE((Xd_0__inst_mult_6_18_q  & Xd_0__inst_mult_6_19_q ))

	.dataa(!Xd_0__inst_mult_6_18_q ),
	.datab(!Xd_0__inst_mult_6_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_209 ),
	.sharein(Xd_0__inst_mult_6_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_212 ),
	.cout(Xd_0__inst_mult_6_213 ),
	.shareout(Xd_0__inst_mult_6_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_79 (
// Equation(s):
// Xd_0__inst_mult_7_216  = SUM(( !Xd_0__inst_mult_7_18_q  $ (!Xd_0__inst_mult_7_19_q ) ) + ( Xd_0__inst_mult_7_214  ) + ( Xd_0__inst_mult_7_213  ))
// Xd_0__inst_mult_7_217  = CARRY(( !Xd_0__inst_mult_7_18_q  $ (!Xd_0__inst_mult_7_19_q ) ) + ( Xd_0__inst_mult_7_214  ) + ( Xd_0__inst_mult_7_213  ))
// Xd_0__inst_mult_7_218  = SHARE((Xd_0__inst_mult_7_18_q  & Xd_0__inst_mult_7_19_q ))

	.dataa(!Xd_0__inst_mult_7_18_q ),
	.datab(!Xd_0__inst_mult_7_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_213 ),
	.sharein(Xd_0__inst_mult_7_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_216 ),
	.cout(Xd_0__inst_mult_7_217 ),
	.shareout(Xd_0__inst_mult_7_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_79 (
// Equation(s):
// Xd_0__inst_mult_6_216  = SUM(( !Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q  $ (((Xd_0__inst_mult_6_22_q  & Xd_0__inst_mult_6_23_q )))) ) + ( Xd_0__inst_mult_6_214  ) + ( Xd_0__inst_mult_6_213  ))
// Xd_0__inst_mult_6_217  = CARRY(( !Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q  $ (((Xd_0__inst_mult_6_22_q  & Xd_0__inst_mult_6_23_q )))) ) + ( Xd_0__inst_mult_6_214  ) + ( Xd_0__inst_mult_6_213  ))
// Xd_0__inst_mult_6_218  = SHARE((Xd_0__inst_mult_6_22_q  & (Xd_0__inst_mult_6_23_q  & (!Xd_0__inst_mult_6_20_q  $ (!Xd_0__inst_mult_6_21_q )))))

	.dataa(!Xd_0__inst_mult_6_20_q ),
	.datab(!Xd_0__inst_mult_6_21_q ),
	.datac(!Xd_0__inst_mult_6_22_q ),
	.datad(!Xd_0__inst_mult_6_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_213 ),
	.sharein(Xd_0__inst_mult_6_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_216 ),
	.cout(Xd_0__inst_mult_6_217 ),
	.shareout(Xd_0__inst_mult_6_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_80 (
// Equation(s):
// Xd_0__inst_mult_7_220  = SUM(( !Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q  $ (((Xd_0__inst_mult_7_22_q  & Xd_0__inst_mult_7_23_q )))) ) + ( Xd_0__inst_mult_7_218  ) + ( Xd_0__inst_mult_7_217  ))
// Xd_0__inst_mult_7_221  = CARRY(( !Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q  $ (((Xd_0__inst_mult_7_22_q  & Xd_0__inst_mult_7_23_q )))) ) + ( Xd_0__inst_mult_7_218  ) + ( Xd_0__inst_mult_7_217  ))
// Xd_0__inst_mult_7_222  = SHARE((Xd_0__inst_mult_7_22_q  & (Xd_0__inst_mult_7_23_q  & (!Xd_0__inst_mult_7_20_q  $ (!Xd_0__inst_mult_7_21_q )))))

	.dataa(!Xd_0__inst_mult_7_20_q ),
	.datab(!Xd_0__inst_mult_7_21_q ),
	.datac(!Xd_0__inst_mult_7_22_q ),
	.datad(!Xd_0__inst_mult_7_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_217 ),
	.sharein(Xd_0__inst_mult_7_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_220 ),
	.cout(Xd_0__inst_mult_7_221 ),
	.shareout(Xd_0__inst_mult_7_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_80 (
// Equation(s):
// Xd_0__inst_mult_6_220  = SUM(( !Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q  $ (((Xd_0__inst_mult_6_20_q  & Xd_0__inst_mult_6_21_q )))) ) + ( Xd_0__inst_mult_6_218  ) + ( Xd_0__inst_mult_6_217  ))
// Xd_0__inst_mult_6_221  = CARRY(( !Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q  $ (((Xd_0__inst_mult_6_20_q  & Xd_0__inst_mult_6_21_q )))) ) + ( Xd_0__inst_mult_6_218  ) + ( Xd_0__inst_mult_6_217  ))
// Xd_0__inst_mult_6_222  = SHARE((Xd_0__inst_mult_6_20_q  & (Xd_0__inst_mult_6_21_q  & (!Xd_0__inst_mult_6_24_q  $ (!Xd_0__inst_mult_6_25_q )))))

	.dataa(!Xd_0__inst_mult_6_24_q ),
	.datab(!Xd_0__inst_mult_6_25_q ),
	.datac(!Xd_0__inst_mult_6_20_q ),
	.datad(!Xd_0__inst_mult_6_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_217 ),
	.sharein(Xd_0__inst_mult_6_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_220 ),
	.cout(Xd_0__inst_mult_6_221 ),
	.shareout(Xd_0__inst_mult_6_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_81 (
// Equation(s):
// Xd_0__inst_mult_7_224  = SUM(( !Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q  $ (((Xd_0__inst_mult_7_20_q  & Xd_0__inst_mult_7_21_q )))) ) + ( Xd_0__inst_mult_7_222  ) + ( Xd_0__inst_mult_7_221  ))
// Xd_0__inst_mult_7_225  = CARRY(( !Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q  $ (((Xd_0__inst_mult_7_20_q  & Xd_0__inst_mult_7_21_q )))) ) + ( Xd_0__inst_mult_7_222  ) + ( Xd_0__inst_mult_7_221  ))
// Xd_0__inst_mult_7_226  = SHARE((Xd_0__inst_mult_7_20_q  & (Xd_0__inst_mult_7_21_q  & (!Xd_0__inst_mult_7_24_q  $ (!Xd_0__inst_mult_7_25_q )))))

	.dataa(!Xd_0__inst_mult_7_24_q ),
	.datab(!Xd_0__inst_mult_7_25_q ),
	.datac(!Xd_0__inst_mult_7_20_q ),
	.datad(!Xd_0__inst_mult_7_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_221 ),
	.sharein(Xd_0__inst_mult_7_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_224 ),
	.cout(Xd_0__inst_mult_7_225 ),
	.shareout(Xd_0__inst_mult_7_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_81 (
// Equation(s):
// Xd_0__inst_mult_6_224  = SUM(( !Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q  $ (((Xd_0__inst_mult_6_24_q  & Xd_0__inst_mult_6_25_q )))) ) + ( Xd_0__inst_mult_6_222  ) + ( Xd_0__inst_mult_6_221  ))
// Xd_0__inst_mult_6_225  = CARRY(( !Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q  $ (((Xd_0__inst_mult_6_24_q  & Xd_0__inst_mult_6_25_q )))) ) + ( Xd_0__inst_mult_6_222  ) + ( Xd_0__inst_mult_6_221  ))
// Xd_0__inst_mult_6_226  = SHARE((Xd_0__inst_mult_6_24_q  & (Xd_0__inst_mult_6_25_q  & (!Xd_0__inst_mult_6_26_q  $ (!Xd_0__inst_mult_6_27_q )))))

	.dataa(!Xd_0__inst_mult_6_26_q ),
	.datab(!Xd_0__inst_mult_6_27_q ),
	.datac(!Xd_0__inst_mult_6_24_q ),
	.datad(!Xd_0__inst_mult_6_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_221 ),
	.sharein(Xd_0__inst_mult_6_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_224 ),
	.cout(Xd_0__inst_mult_6_225 ),
	.shareout(Xd_0__inst_mult_6_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_82 (
// Equation(s):
// Xd_0__inst_mult_7_228  = SUM(( !Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q  $ (((Xd_0__inst_mult_7_24_q  & Xd_0__inst_mult_7_25_q )))) ) + ( Xd_0__inst_mult_7_226  ) + ( Xd_0__inst_mult_7_225  ))
// Xd_0__inst_mult_7_229  = CARRY(( !Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q  $ (((Xd_0__inst_mult_7_24_q  & Xd_0__inst_mult_7_25_q )))) ) + ( Xd_0__inst_mult_7_226  ) + ( Xd_0__inst_mult_7_225  ))
// Xd_0__inst_mult_7_230  = SHARE((Xd_0__inst_mult_7_24_q  & (Xd_0__inst_mult_7_25_q  & (!Xd_0__inst_mult_7_26_q  $ (!Xd_0__inst_mult_7_27_q )))))

	.dataa(!Xd_0__inst_mult_7_26_q ),
	.datab(!Xd_0__inst_mult_7_27_q ),
	.datac(!Xd_0__inst_mult_7_24_q ),
	.datad(!Xd_0__inst_mult_7_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_225 ),
	.sharein(Xd_0__inst_mult_7_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_228 ),
	.cout(Xd_0__inst_mult_7_229 ),
	.shareout(Xd_0__inst_mult_7_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_82 (
// Equation(s):
// Xd_0__inst_mult_6_228  = SUM(( !Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q  $ (((Xd_0__inst_mult_6_26_q  & Xd_0__inst_mult_6_27_q )))) ) + ( Xd_0__inst_mult_6_226  ) + ( Xd_0__inst_mult_6_225  ))
// Xd_0__inst_mult_6_229  = CARRY(( !Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q  $ (((Xd_0__inst_mult_6_26_q  & Xd_0__inst_mult_6_27_q )))) ) + ( Xd_0__inst_mult_6_226  ) + ( Xd_0__inst_mult_6_225  ))
// Xd_0__inst_mult_6_230  = SHARE((Xd_0__inst_mult_6_26_q  & (Xd_0__inst_mult_6_27_q  & (!Xd_0__inst_mult_6_28_q  $ (!Xd_0__inst_mult_6_29_q )))))

	.dataa(!Xd_0__inst_mult_6_28_q ),
	.datab(!Xd_0__inst_mult_6_29_q ),
	.datac(!Xd_0__inst_mult_6_26_q ),
	.datad(!Xd_0__inst_mult_6_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_225 ),
	.sharein(Xd_0__inst_mult_6_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_228 ),
	.cout(Xd_0__inst_mult_6_229 ),
	.shareout(Xd_0__inst_mult_6_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_83 (
// Equation(s):
// Xd_0__inst_mult_7_232  = SUM(( !Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q  $ (((Xd_0__inst_mult_7_26_q  & Xd_0__inst_mult_7_27_q )))) ) + ( Xd_0__inst_mult_7_230  ) + ( Xd_0__inst_mult_7_229  ))
// Xd_0__inst_mult_7_233  = CARRY(( !Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q  $ (((Xd_0__inst_mult_7_26_q  & Xd_0__inst_mult_7_27_q )))) ) + ( Xd_0__inst_mult_7_230  ) + ( Xd_0__inst_mult_7_229  ))
// Xd_0__inst_mult_7_234  = SHARE((Xd_0__inst_mult_7_26_q  & (Xd_0__inst_mult_7_27_q  & (!Xd_0__inst_mult_7_28_q  $ (!Xd_0__inst_mult_7_29_q )))))

	.dataa(!Xd_0__inst_mult_7_28_q ),
	.datab(!Xd_0__inst_mult_7_29_q ),
	.datac(!Xd_0__inst_mult_7_26_q ),
	.datad(!Xd_0__inst_mult_7_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_229 ),
	.sharein(Xd_0__inst_mult_7_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_232 ),
	.cout(Xd_0__inst_mult_7_233 ),
	.shareout(Xd_0__inst_mult_7_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_83 (
// Equation(s):
// Xd_0__inst_mult_6_232  = SUM(( !Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q  $ (((Xd_0__inst_mult_6_28_q  & Xd_0__inst_mult_6_29_q )))) ) + ( Xd_0__inst_mult_6_230  ) + ( Xd_0__inst_mult_6_229  ))
// Xd_0__inst_mult_6_233  = CARRY(( !Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q  $ (((Xd_0__inst_mult_6_28_q  & Xd_0__inst_mult_6_29_q )))) ) + ( Xd_0__inst_mult_6_230  ) + ( Xd_0__inst_mult_6_229  ))
// Xd_0__inst_mult_6_234  = SHARE((Xd_0__inst_mult_6_28_q  & (Xd_0__inst_mult_6_29_q  & (!Xd_0__inst_mult_6_30_q  $ (!Xd_0__inst_mult_6_31_q )))))

	.dataa(!Xd_0__inst_mult_6_30_q ),
	.datab(!Xd_0__inst_mult_6_31_q ),
	.datac(!Xd_0__inst_mult_6_28_q ),
	.datad(!Xd_0__inst_mult_6_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_229 ),
	.sharein(Xd_0__inst_mult_6_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_232 ),
	.cout(Xd_0__inst_mult_6_233 ),
	.shareout(Xd_0__inst_mult_6_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_84 (
// Equation(s):
// Xd_0__inst_mult_7_236  = SUM(( !Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q  $ (((Xd_0__inst_mult_7_28_q  & Xd_0__inst_mult_7_29_q )))) ) + ( Xd_0__inst_mult_7_234  ) + ( Xd_0__inst_mult_7_233  ))
// Xd_0__inst_mult_7_237  = CARRY(( !Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q  $ (((Xd_0__inst_mult_7_28_q  & Xd_0__inst_mult_7_29_q )))) ) + ( Xd_0__inst_mult_7_234  ) + ( Xd_0__inst_mult_7_233  ))
// Xd_0__inst_mult_7_238  = SHARE((Xd_0__inst_mult_7_28_q  & (Xd_0__inst_mult_7_29_q  & (!Xd_0__inst_mult_7_30_q  $ (!Xd_0__inst_mult_7_31_q )))))

	.dataa(!Xd_0__inst_mult_7_30_q ),
	.datab(!Xd_0__inst_mult_7_31_q ),
	.datac(!Xd_0__inst_mult_7_28_q ),
	.datad(!Xd_0__inst_mult_7_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_233 ),
	.sharein(Xd_0__inst_mult_7_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_236 ),
	.cout(Xd_0__inst_mult_7_237 ),
	.shareout(Xd_0__inst_mult_7_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_84 (
// Equation(s):
// Xd_0__inst_mult_6_236  = SUM(( !Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q  $ (((Xd_0__inst_mult_6_30_q  & Xd_0__inst_mult_6_31_q )))) ) + ( Xd_0__inst_mult_6_234  ) + ( Xd_0__inst_mult_6_233  ))
// Xd_0__inst_mult_6_237  = CARRY(( !Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q  $ (((Xd_0__inst_mult_6_30_q  & Xd_0__inst_mult_6_31_q )))) ) + ( Xd_0__inst_mult_6_234  ) + ( Xd_0__inst_mult_6_233  ))
// Xd_0__inst_mult_6_238  = SHARE((Xd_0__inst_mult_6_30_q  & (Xd_0__inst_mult_6_31_q  & (!Xd_0__inst_mult_6_32_q  $ (!Xd_0__inst_mult_6_33_q )))))

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(!Xd_0__inst_mult_6_30_q ),
	.datad(!Xd_0__inst_mult_6_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_233 ),
	.sharein(Xd_0__inst_mult_6_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_236 ),
	.cout(Xd_0__inst_mult_6_237 ),
	.shareout(Xd_0__inst_mult_6_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_85 (
// Equation(s):
// Xd_0__inst_mult_7_240  = SUM(( !Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q  $ (((Xd_0__inst_mult_7_30_q  & Xd_0__inst_mult_7_31_q )))) ) + ( Xd_0__inst_mult_7_238  ) + ( Xd_0__inst_mult_7_237  ))
// Xd_0__inst_mult_7_241  = CARRY(( !Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q  $ (((Xd_0__inst_mult_7_30_q  & Xd_0__inst_mult_7_31_q )))) ) + ( Xd_0__inst_mult_7_238  ) + ( Xd_0__inst_mult_7_237  ))
// Xd_0__inst_mult_7_242  = SHARE((Xd_0__inst_mult_7_30_q  & (Xd_0__inst_mult_7_31_q  & (!Xd_0__inst_mult_7_32_q  $ (!Xd_0__inst_mult_7_33_q )))))

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(!Xd_0__inst_mult_7_30_q ),
	.datad(!Xd_0__inst_mult_7_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_237 ),
	.sharein(Xd_0__inst_mult_7_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_240 ),
	.cout(Xd_0__inst_mult_7_241 ),
	.shareout(Xd_0__inst_mult_7_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_85 (
// Equation(s):
// Xd_0__inst_mult_6_240  = SUM(( (Xd_0__inst_mult_6_32_q  & Xd_0__inst_mult_6_33_q ) ) + ( Xd_0__inst_mult_6_238  ) + ( Xd_0__inst_mult_6_237  ))

	.dataa(!Xd_0__inst_mult_6_32_q ),
	.datab(!Xd_0__inst_mult_6_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_237 ),
	.sharein(Xd_0__inst_mult_6_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_240 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_86 (
// Equation(s):
// Xd_0__inst_mult_7_244  = SUM(( (Xd_0__inst_mult_7_32_q  & Xd_0__inst_mult_7_33_q ) ) + ( Xd_0__inst_mult_7_242  ) + ( Xd_0__inst_mult_7_241  ))

	.dataa(!Xd_0__inst_mult_7_32_q ),
	.datab(!Xd_0__inst_mult_7_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_241 ),
	.sharein(Xd_0__inst_mult_7_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_244 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_68 (
// Equation(s):
// Xd_0__inst_mult_3_184  = SUM(( !Xd_0__inst_mult_3_260  $ (((!din_b[40]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_266  ) + ( Xd_0__inst_mult_3_265  ))
// Xd_0__inst_mult_3_185  = CARRY(( !Xd_0__inst_mult_3_260  $ (((!din_b[40]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_266  ) + ( Xd_0__inst_mult_3_265  ))
// Xd_0__inst_mult_3_186  = SHARE((din_b[40] & (din_a[46] & Xd_0__inst_mult_3_260 )))

	.dataa(!din_b[40]),
	.datab(!din_a[46]),
	.datac(!Xd_0__inst_mult_3_260 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_265 ),
	.sharein(Xd_0__inst_mult_3_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_184 ),
	.cout(Xd_0__inst_mult_3_185 ),
	.shareout(Xd_0__inst_mult_3_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_86 (
// Equation(s):
// Xd_0__inst_mult_6_244  = SUM(( !Xd_0__inst_mult_6_268  $ (((!din_b[76]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_274  ) + ( Xd_0__inst_mult_6_273  ))
// Xd_0__inst_mult_6_245  = CARRY(( !Xd_0__inst_mult_6_268  $ (((!din_b[76]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_274  ) + ( Xd_0__inst_mult_6_273  ))
// Xd_0__inst_mult_6_246  = SHARE((din_b[76] & (din_a[82] & Xd_0__inst_mult_6_268 )))

	.dataa(!din_b[76]),
	.datab(!din_a[82]),
	.datac(!Xd_0__inst_mult_6_268 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_273 ),
	.sharein(Xd_0__inst_mult_6_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_244 ),
	.cout(Xd_0__inst_mult_6_245 ),
	.shareout(Xd_0__inst_mult_6_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0 (
// Equation(s):
// Xd_0__inst_mult_0_173  = SUM(( !Xd_0__inst_mult_0_248  $ (((!din_b[4]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_254  ) + ( Xd_0__inst_mult_0_253  ))
// Xd_0__inst_mult_0_174  = CARRY(( !Xd_0__inst_mult_0_248  $ (((!din_b[4]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_254  ) + ( Xd_0__inst_mult_0_253  ))
// Xd_0__inst_mult_0_175  = SHARE((din_b[4] & (din_a[10] & Xd_0__inst_mult_0_248 )))

	.dataa(!din_b[4]),
	.datab(!din_a[10]),
	.datac(!Xd_0__inst_mult_0_248 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_253 ),
	.sharein(Xd_0__inst_mult_0_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_173 ),
	.cout(Xd_0__inst_mult_0_174 ),
	.shareout(Xd_0__inst_mult_0_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_69 (
// Equation(s):
// Xd_0__inst_mult_3_188  = SUM(( (!din_a[43] & (((din_a[42] & din_b[46])))) # (din_a[43] & (!din_b[45] $ (((!din_a[42]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_274  ) + ( Xd_0__inst_mult_3_273  ))
// Xd_0__inst_mult_3_189  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[46])))) # (din_a[43] & (!din_b[45] $ (((!din_a[42]) # (!din_b[46]))))) ) + ( Xd_0__inst_mult_3_274  ) + ( Xd_0__inst_mult_3_273  ))
// Xd_0__inst_mult_3_190  = SHARE((din_a[43] & (din_b[45] & (din_a[42] & din_b[46]))))

	.dataa(!din_a[43]),
	.datab(!din_b[45]),
	.datac(!din_a[42]),
	.datad(!din_b[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_273 ),
	.sharein(Xd_0__inst_mult_3_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_188 ),
	.cout(Xd_0__inst_mult_3_189 ),
	.shareout(Xd_0__inst_mult_3_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_87 (
// Equation(s):
// Xd_0__inst_mult_6_248  = SUM(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_249  = CARRY(( (din_a[72] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_250  = SHARE((din_a[72] & din_b[73]))

	.dataa(!din_a[72]),
	.datab(!din_b[72]),
	.datac(!din_b[73]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_248 ),
	.cout(Xd_0__inst_mult_6_249 ),
	.shareout(Xd_0__inst_mult_6_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_87 (
// Equation(s):
// Xd_0__inst_mult_7_248  = SUM(( (din_a[84] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_249  = CARRY(( (din_a[84] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_250  = SHARE((din_a[84] & din_b[85]))

	.dataa(!din_a[84]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_248 ),
	.cout(Xd_0__inst_mult_7_249 ),
	.shareout(Xd_0__inst_mult_7_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_1 (
// Equation(s):
// Xd_0__inst_i29_1_sumout  = SUM(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i29_7  ) + ( Xd_0__inst_i29_6  ))
// Xd_0__inst_i29_2  = CARRY(( !din_a[83] $ (!din_b[83]) ) + ( Xd_0__inst_i29_7  ) + ( Xd_0__inst_i29_6  ))
// Xd_0__inst_i29_3  = SHARE(GND)

	.dataa(!din_a[83]),
	.datab(!din_b[83]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_6 ),
	.sharein(Xd_0__inst_i29_7 ),
	.combout(),
	.sumout(Xd_0__inst_i29_1_sumout ),
	.cout(Xd_0__inst_i29_2 ),
	.shareout(Xd_0__inst_i29_3 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_5 (
// Equation(s):
// Xd_0__inst_i29_5_sumout  = SUM(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i29_11  ) + ( Xd_0__inst_i29_10  ))
// Xd_0__inst_i29_6  = CARRY(( !din_a[95] $ (!din_b[95]) ) + ( Xd_0__inst_i29_11  ) + ( Xd_0__inst_i29_10  ))
// Xd_0__inst_i29_7  = SHARE(GND)

	.dataa(!din_a[95]),
	.datab(!din_b[95]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_10 ),
	.sharein(Xd_0__inst_i29_11 ),
	.combout(),
	.sumout(Xd_0__inst_i29_5_sumout ),
	.cout(Xd_0__inst_i29_6 ),
	.shareout(Xd_0__inst_i29_7 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_88 (
// Equation(s):
// Xd_0__inst_mult_7_252  = SUM(( GND ) + ( Xd_0__inst_mult_7_278  ) + ( Xd_0__inst_mult_7_277  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_277 ),
	.sharein(Xd_0__inst_mult_7_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_252 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_89 (
// Equation(s):
// Xd_0__inst_mult_7_256  = SUM(( !Xd_0__inst_mult_7_276  $ (((!din_b[87]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_282  ) + ( Xd_0__inst_mult_7_281  ))
// Xd_0__inst_mult_7_257  = CARRY(( !Xd_0__inst_mult_7_276  $ (((!din_b[87]) # (!din_a[94]))) ) + ( Xd_0__inst_mult_7_282  ) + ( Xd_0__inst_mult_7_281  ))
// Xd_0__inst_mult_7_258  = SHARE((din_b[87] & (din_a[94] & Xd_0__inst_mult_7_276 )))

	.dataa(!din_b[87]),
	.datab(!din_a[94]),
	.datac(!Xd_0__inst_mult_7_276 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_281 ),
	.sharein(Xd_0__inst_mult_7_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_256 ),
	.cout(Xd_0__inst_mult_7_257 ),
	.shareout(Xd_0__inst_mult_7_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_88 (
// Equation(s):
// Xd_0__inst_mult_6_252  = SUM(( (din_a[73] & din_b[72]) ) + ( Xd_0__inst_mult_6_250  ) + ( Xd_0__inst_mult_6_249  ))
// Xd_0__inst_mult_6_253  = CARRY(( (din_a[73] & din_b[72]) ) + ( Xd_0__inst_mult_6_250  ) + ( Xd_0__inst_mult_6_249  ))
// Xd_0__inst_mult_6_254  = SHARE((din_a[72] & din_b[74]))

	.dataa(!din_a[73]),
	.datab(!din_b[72]),
	.datac(!din_a[72]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_249 ),
	.sharein(Xd_0__inst_mult_6_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_252 ),
	.cout(Xd_0__inst_mult_6_253 ),
	.shareout(Xd_0__inst_mult_6_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_90 (
// Equation(s):
// Xd_0__inst_mult_7_260  = SUM(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_7_250  ) + ( Xd_0__inst_mult_7_249  ))
// Xd_0__inst_mult_7_261  = CARRY(( (din_a[85] & din_b[84]) ) + ( Xd_0__inst_mult_7_250  ) + ( Xd_0__inst_mult_7_249  ))
// Xd_0__inst_mult_7_262  = SHARE((din_a[84] & din_b[86]))

	.dataa(!din_a[85]),
	.datab(!din_b[84]),
	.datac(!din_a[84]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_249 ),
	.sharein(Xd_0__inst_mult_7_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_260 ),
	.cout(Xd_0__inst_mult_7_261 ),
	.shareout(Xd_0__inst_mult_7_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_89 (
// Equation(s):
// Xd_0__inst_mult_6_256  = SUM(( (!din_a[73] & (((din_a[74] & din_b[72])))) # (din_a[73] & (!din_b[73] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_254  ) + ( Xd_0__inst_mult_6_253  ))
// Xd_0__inst_mult_6_257  = CARRY(( (!din_a[73] & (((din_a[74] & din_b[72])))) # (din_a[73] & (!din_b[73] $ (((!din_a[74]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_254  ) + ( Xd_0__inst_mult_6_253  ))
// Xd_0__inst_mult_6_258  = SHARE((din_a[73] & (din_b[73] & (din_a[74] & din_b[72]))))

	.dataa(!din_a[73]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_253 ),
	.sharein(Xd_0__inst_mult_6_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_256 ),
	.cout(Xd_0__inst_mult_6_257 ),
	.shareout(Xd_0__inst_mult_6_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_91 (
// Equation(s):
// Xd_0__inst_mult_7_264  = SUM(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_262  ) + ( Xd_0__inst_mult_7_261  ))
// Xd_0__inst_mult_7_265  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[84])))) # (din_a[85] & (!din_b[85] $ (((!din_a[86]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_262  ) + ( Xd_0__inst_mult_7_261  ))
// Xd_0__inst_mult_7_266  = SHARE((din_a[85] & (din_b[85] & (din_a[86] & din_b[84]))))

	.dataa(!din_a[85]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_261 ),
	.sharein(Xd_0__inst_mult_7_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_264 ),
	.cout(Xd_0__inst_mult_7_265 ),
	.shareout(Xd_0__inst_mult_7_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_90 (
// Equation(s):
// Xd_0__inst_mult_6_260  = SUM(( (din_a[72] & din_b[75]) ) + ( Xd_0__inst_mult_6_278  ) + ( Xd_0__inst_mult_6_277  ))
// Xd_0__inst_mult_6_261  = CARRY(( (din_a[72] & din_b[75]) ) + ( Xd_0__inst_mult_6_278  ) + ( Xd_0__inst_mult_6_277  ))
// Xd_0__inst_mult_6_262  = SHARE((din_a[72] & din_b[76]))

	.dataa(!din_a[72]),
	.datab(!din_b[75]),
	.datac(!din_b[76]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_277 ),
	.sharein(Xd_0__inst_mult_6_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_260 ),
	.cout(Xd_0__inst_mult_6_261 ),
	.shareout(Xd_0__inst_mult_6_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_92 (
// Equation(s):
// Xd_0__inst_mult_7_268  = SUM(( (din_a[84] & din_b[87]) ) + ( Xd_0__inst_mult_7_286  ) + ( Xd_0__inst_mult_7_285  ))
// Xd_0__inst_mult_7_269  = CARRY(( (din_a[84] & din_b[87]) ) + ( Xd_0__inst_mult_7_286  ) + ( Xd_0__inst_mult_7_285  ))
// Xd_0__inst_mult_7_270  = SHARE((din_a[84] & din_b[88]))

	.dataa(!din_a[84]),
	.datab(!din_b[87]),
	.datac(!din_b[88]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_285 ),
	.sharein(Xd_0__inst_mult_7_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_268 ),
	.cout(Xd_0__inst_mult_7_269 ),
	.shareout(Xd_0__inst_mult_7_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_91 (
// Equation(s):
// Xd_0__inst_mult_6_264  = SUM(( !Xd_0__inst_mult_6_280  $ (!Xd_0__inst_mult_6_284 ) ) + ( Xd_0__inst_mult_6_262  ) + ( Xd_0__inst_mult_6_261  ))
// Xd_0__inst_mult_6_265  = CARRY(( !Xd_0__inst_mult_6_280  $ (!Xd_0__inst_mult_6_284 ) ) + ( Xd_0__inst_mult_6_262  ) + ( Xd_0__inst_mult_6_261  ))
// Xd_0__inst_mult_6_266  = SHARE((Xd_0__inst_mult_6_280  & Xd_0__inst_mult_6_284 ))

	.dataa(!Xd_0__inst_mult_6_280 ),
	.datab(!Xd_0__inst_mult_6_284 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_261 ),
	.sharein(Xd_0__inst_mult_6_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_264 ),
	.cout(Xd_0__inst_mult_6_265 ),
	.shareout(Xd_0__inst_mult_6_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_93 (
// Equation(s):
// Xd_0__inst_mult_7_272  = SUM(( !Xd_0__inst_mult_7_288  $ (!Xd_0__inst_mult_7_292 ) ) + ( Xd_0__inst_mult_7_270  ) + ( Xd_0__inst_mult_7_269  ))
// Xd_0__inst_mult_7_273  = CARRY(( !Xd_0__inst_mult_7_288  $ (!Xd_0__inst_mult_7_292 ) ) + ( Xd_0__inst_mult_7_270  ) + ( Xd_0__inst_mult_7_269  ))
// Xd_0__inst_mult_7_274  = SHARE((Xd_0__inst_mult_7_288  & Xd_0__inst_mult_7_292 ))

	.dataa(!Xd_0__inst_mult_7_288 ),
	.datab(!Xd_0__inst_mult_7_292 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_269 ),
	.sharein(Xd_0__inst_mult_7_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_272 ),
	.cout(Xd_0__inst_mult_7_273 ),
	.shareout(Xd_0__inst_mult_7_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_172 (
// Equation(s):
// Xd_0__inst_mult_4_173  = SUM(( !Xd_0__inst_mult_4_0_q  $ (!Xd_0__inst_mult_4_1_q ) ) + ( Xd_0__inst_mult_2_37  ) + ( Xd_0__inst_mult_2_36  ))
// Xd_0__inst_mult_4_174  = CARRY(( !Xd_0__inst_mult_4_0_q  $ (!Xd_0__inst_mult_4_1_q ) ) + ( Xd_0__inst_mult_2_37  ) + ( Xd_0__inst_mult_2_36  ))
// Xd_0__inst_mult_4_175  = SHARE((Xd_0__inst_mult_4_0_q  & Xd_0__inst_mult_4_1_q ))

	.dataa(!Xd_0__inst_mult_4_0_q ),
	.datab(!Xd_0__inst_mult_4_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_36 ),
	.sharein(Xd_0__inst_mult_2_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_173 ),
	.cout(Xd_0__inst_mult_4_174 ),
	.shareout(Xd_0__inst_mult_4_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_172 (
// Equation(s):
// Xd_0__inst_mult_5_173  = SUM(( !Xd_0__inst_mult_5_0_q  $ (!Xd_0__inst_mult_5_1_q ) ) + ( Xd_0__inst_mult_0_37  ) + ( Xd_0__inst_mult_0_36  ))
// Xd_0__inst_mult_5_174  = CARRY(( !Xd_0__inst_mult_5_0_q  $ (!Xd_0__inst_mult_5_1_q ) ) + ( Xd_0__inst_mult_0_37  ) + ( Xd_0__inst_mult_0_36  ))
// Xd_0__inst_mult_5_175  = SHARE((Xd_0__inst_mult_5_0_q  & Xd_0__inst_mult_5_1_q ))

	.dataa(!Xd_0__inst_mult_5_0_q ),
	.datab(!Xd_0__inst_mult_5_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_36 ),
	.sharein(Xd_0__inst_mult_0_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_173 ),
	.cout(Xd_0__inst_mult_5_174 ),
	.shareout(Xd_0__inst_mult_5_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_172 (
// Equation(s):
// Xd_0__inst_mult_2_173  = SUM(( !Xd_0__inst_mult_2_0_q  $ (!Xd_0__inst_mult_2_1_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_174  = CARRY(( !Xd_0__inst_mult_2_0_q  $ (!Xd_0__inst_mult_2_1_q ) ) + ( Xd_0__inst_mult_2_41  ) + ( Xd_0__inst_mult_2_40  ))
// Xd_0__inst_mult_2_175  = SHARE((Xd_0__inst_mult_2_0_q  & Xd_0__inst_mult_2_1_q ))

	.dataa(!Xd_0__inst_mult_2_0_q ),
	.datab(!Xd_0__inst_mult_2_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_40 ),
	.sharein(Xd_0__inst_mult_2_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_173 ),
	.cout(Xd_0__inst_mult_2_174 ),
	.shareout(Xd_0__inst_mult_2_175 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_70 (
// Equation(s):
// Xd_0__inst_mult_3_192  = SUM(( !Xd_0__inst_mult_3_0_q  $ (!Xd_0__inst_mult_3_1_q ) ) + ( Xd_0__inst_mult_1_37  ) + ( Xd_0__inst_mult_1_36  ))
// Xd_0__inst_mult_3_193  = CARRY(( !Xd_0__inst_mult_3_0_q  $ (!Xd_0__inst_mult_3_1_q ) ) + ( Xd_0__inst_mult_1_37  ) + ( Xd_0__inst_mult_1_36  ))
// Xd_0__inst_mult_3_194  = SHARE((Xd_0__inst_mult_3_0_q  & Xd_0__inst_mult_3_1_q ))

	.dataa(!Xd_0__inst_mult_3_0_q ),
	.datab(!Xd_0__inst_mult_3_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_36 ),
	.sharein(Xd_0__inst_mult_1_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_192 ),
	.cout(Xd_0__inst_mult_3_193 ),
	.shareout(Xd_0__inst_mult_3_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_66 (
// Equation(s):
// Xd_0__inst_mult_0_176  = SUM(( !Xd_0__inst_mult_0_0_q  $ (!Xd_0__inst_mult_0_1_q ) ) + ( Xd_0__inst_mult_2_45  ) + ( Xd_0__inst_mult_2_44  ))
// Xd_0__inst_mult_0_177  = CARRY(( !Xd_0__inst_mult_0_0_q  $ (!Xd_0__inst_mult_0_1_q ) ) + ( Xd_0__inst_mult_2_45  ) + ( Xd_0__inst_mult_2_44  ))
// Xd_0__inst_mult_0_178  = SHARE((Xd_0__inst_mult_0_0_q  & Xd_0__inst_mult_0_1_q ))

	.dataa(!Xd_0__inst_mult_0_0_q ),
	.datab(!Xd_0__inst_mult_0_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_44 ),
	.sharein(Xd_0__inst_mult_2_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_176 ),
	.cout(Xd_0__inst_mult_0_177 ),
	.shareout(Xd_0__inst_mult_0_178 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_69 (
// Equation(s):
// Xd_0__inst_mult_1_188  = SUM(( !Xd_0__inst_mult_1_0_q  $ (!Xd_0__inst_mult_1_1_q ) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_1_189  = CARRY(( !Xd_0__inst_mult_1_0_q  $ (!Xd_0__inst_mult_1_1_q ) ) + ( Xd_0__inst_mult_1_41  ) + ( Xd_0__inst_mult_1_40  ))
// Xd_0__inst_mult_1_190  = SHARE((Xd_0__inst_mult_1_0_q  & Xd_0__inst_mult_1_1_q ))

	.dataa(!Xd_0__inst_mult_1_0_q ),
	.datab(!Xd_0__inst_mult_1_1_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_40 ),
	.sharein(Xd_0__inst_mult_1_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_188 ),
	.cout(Xd_0__inst_mult_1_189 ),
	.shareout(Xd_0__inst_mult_1_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_35 (
// Equation(s):
// Xd_0__inst_mult_4_35_sumout  = SUM(( (din_a[58] & din_b[48]) ) + ( Xd_0__inst_mult_1_45  ) + ( Xd_0__inst_mult_1_44  ))
// Xd_0__inst_mult_4_36  = CARRY(( (din_a[58] & din_b[48]) ) + ( Xd_0__inst_mult_1_45  ) + ( Xd_0__inst_mult_1_44  ))
// Xd_0__inst_mult_4_37  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_44 ),
	.sharein(Xd_0__inst_mult_1_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_35_sumout ),
	.cout(Xd_0__inst_mult_4_36 ),
	.shareout(Xd_0__inst_mult_4_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_35 (
// Equation(s):
// Xd_0__inst_mult_3_35_sumout  = SUM(( (din_a[46] & din_b[36]) ) + ( Xd_0__inst_mult_2_49  ) + ( Xd_0__inst_mult_2_48  ))
// Xd_0__inst_mult_3_36  = CARRY(( (din_a[46] & din_b[36]) ) + ( Xd_0__inst_mult_2_49  ) + ( Xd_0__inst_mult_2_48  ))
// Xd_0__inst_mult_3_37  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_48 ),
	.sharein(Xd_0__inst_mult_2_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_35_sumout ),
	.cout(Xd_0__inst_mult_3_36 ),
	.shareout(Xd_0__inst_mult_3_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4 (
// Equation(s):
// Xd_0__inst_mult_4_177  = SUM(( !Xd_0__inst_mult_4_2_q  $ (!Xd_0__inst_mult_4_3_q ) ) + ( Xd_0__inst_mult_4_175  ) + ( Xd_0__inst_mult_4_174  ))
// Xd_0__inst_mult_4_178  = CARRY(( !Xd_0__inst_mult_4_2_q  $ (!Xd_0__inst_mult_4_3_q ) ) + ( Xd_0__inst_mult_4_175  ) + ( Xd_0__inst_mult_4_174  ))
// Xd_0__inst_mult_4_179  = SHARE((Xd_0__inst_mult_4_2_q  & Xd_0__inst_mult_4_3_q ))

	.dataa(!Xd_0__inst_mult_4_2_q ),
	.datab(!Xd_0__inst_mult_4_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_174 ),
	.sharein(Xd_0__inst_mult_4_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_177 ),
	.cout(Xd_0__inst_mult_4_178 ),
	.shareout(Xd_0__inst_mult_4_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5 (
// Equation(s):
// Xd_0__inst_mult_5_177  = SUM(( !Xd_0__inst_mult_5_2_q  $ (!Xd_0__inst_mult_5_3_q ) ) + ( Xd_0__inst_mult_5_175  ) + ( Xd_0__inst_mult_5_174  ))
// Xd_0__inst_mult_5_178  = CARRY(( !Xd_0__inst_mult_5_2_q  $ (!Xd_0__inst_mult_5_3_q ) ) + ( Xd_0__inst_mult_5_175  ) + ( Xd_0__inst_mult_5_174  ))
// Xd_0__inst_mult_5_179  = SHARE((Xd_0__inst_mult_5_2_q  & Xd_0__inst_mult_5_3_q ))

	.dataa(!Xd_0__inst_mult_5_2_q ),
	.datab(!Xd_0__inst_mult_5_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_174 ),
	.sharein(Xd_0__inst_mult_5_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_177 ),
	.cout(Xd_0__inst_mult_5_178 ),
	.shareout(Xd_0__inst_mult_5_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2 (
// Equation(s):
// Xd_0__inst_mult_2_177  = SUM(( !Xd_0__inst_mult_2_2_q  $ (!Xd_0__inst_mult_2_3_q ) ) + ( Xd_0__inst_mult_2_175  ) + ( Xd_0__inst_mult_2_174  ))
// Xd_0__inst_mult_2_178  = CARRY(( !Xd_0__inst_mult_2_2_q  $ (!Xd_0__inst_mult_2_3_q ) ) + ( Xd_0__inst_mult_2_175  ) + ( Xd_0__inst_mult_2_174  ))
// Xd_0__inst_mult_2_179  = SHARE((Xd_0__inst_mult_2_2_q  & Xd_0__inst_mult_2_3_q ))

	.dataa(!Xd_0__inst_mult_2_2_q ),
	.datab(!Xd_0__inst_mult_2_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_174 ),
	.sharein(Xd_0__inst_mult_2_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_177 ),
	.cout(Xd_0__inst_mult_2_178 ),
	.shareout(Xd_0__inst_mult_2_179 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_71 (
// Equation(s):
// Xd_0__inst_mult_3_196  = SUM(( !Xd_0__inst_mult_3_2_q  $ (!Xd_0__inst_mult_3_3_q ) ) + ( Xd_0__inst_mult_3_194  ) + ( Xd_0__inst_mult_3_193  ))
// Xd_0__inst_mult_3_197  = CARRY(( !Xd_0__inst_mult_3_2_q  $ (!Xd_0__inst_mult_3_3_q ) ) + ( Xd_0__inst_mult_3_194  ) + ( Xd_0__inst_mult_3_193  ))
// Xd_0__inst_mult_3_198  = SHARE((Xd_0__inst_mult_3_2_q  & Xd_0__inst_mult_3_3_q ))

	.dataa(!Xd_0__inst_mult_3_2_q ),
	.datab(!Xd_0__inst_mult_3_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_193 ),
	.sharein(Xd_0__inst_mult_3_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_196 ),
	.cout(Xd_0__inst_mult_3_197 ),
	.shareout(Xd_0__inst_mult_3_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_67 (
// Equation(s):
// Xd_0__inst_mult_0_180  = SUM(( !Xd_0__inst_mult_0_2_q  $ (!Xd_0__inst_mult_0_3_q ) ) + ( Xd_0__inst_mult_0_178  ) + ( Xd_0__inst_mult_0_177  ))
// Xd_0__inst_mult_0_181  = CARRY(( !Xd_0__inst_mult_0_2_q  $ (!Xd_0__inst_mult_0_3_q ) ) + ( Xd_0__inst_mult_0_178  ) + ( Xd_0__inst_mult_0_177  ))
// Xd_0__inst_mult_0_182  = SHARE((Xd_0__inst_mult_0_2_q  & Xd_0__inst_mult_0_3_q ))

	.dataa(!Xd_0__inst_mult_0_2_q ),
	.datab(!Xd_0__inst_mult_0_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_177 ),
	.sharein(Xd_0__inst_mult_0_178 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_180 ),
	.cout(Xd_0__inst_mult_0_181 ),
	.shareout(Xd_0__inst_mult_0_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_70 (
// Equation(s):
// Xd_0__inst_mult_1_192  = SUM(( !Xd_0__inst_mult_1_2_q  $ (!Xd_0__inst_mult_1_3_q ) ) + ( Xd_0__inst_mult_1_190  ) + ( Xd_0__inst_mult_1_189  ))
// Xd_0__inst_mult_1_193  = CARRY(( !Xd_0__inst_mult_1_2_q  $ (!Xd_0__inst_mult_1_3_q ) ) + ( Xd_0__inst_mult_1_190  ) + ( Xd_0__inst_mult_1_189  ))
// Xd_0__inst_mult_1_194  = SHARE((Xd_0__inst_mult_1_2_q  & Xd_0__inst_mult_1_3_q ))

	.dataa(!Xd_0__inst_mult_1_2_q ),
	.datab(!Xd_0__inst_mult_1_3_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_189 ),
	.sharein(Xd_0__inst_mult_1_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_192 ),
	.cout(Xd_0__inst_mult_1_193 ),
	.shareout(Xd_0__inst_mult_1_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_70 (
// Equation(s):
// Xd_0__inst_mult_4_180  = SUM(( !Xd_0__inst_mult_4_4_q  $ (!Xd_0__inst_mult_4_5_q ) ) + ( Xd_0__inst_mult_4_179  ) + ( Xd_0__inst_mult_4_178  ))
// Xd_0__inst_mult_4_181  = CARRY(( !Xd_0__inst_mult_4_4_q  $ (!Xd_0__inst_mult_4_5_q ) ) + ( Xd_0__inst_mult_4_179  ) + ( Xd_0__inst_mult_4_178  ))
// Xd_0__inst_mult_4_182  = SHARE((Xd_0__inst_mult_4_4_q  & Xd_0__inst_mult_4_5_q ))

	.dataa(!Xd_0__inst_mult_4_4_q ),
	.datab(!Xd_0__inst_mult_4_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_178 ),
	.sharein(Xd_0__inst_mult_4_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_180 ),
	.cout(Xd_0__inst_mult_4_181 ),
	.shareout(Xd_0__inst_mult_4_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_70 (
// Equation(s):
// Xd_0__inst_mult_5_180  = SUM(( !Xd_0__inst_mult_5_4_q  $ (!Xd_0__inst_mult_5_5_q ) ) + ( Xd_0__inst_mult_5_179  ) + ( Xd_0__inst_mult_5_178  ))
// Xd_0__inst_mult_5_181  = CARRY(( !Xd_0__inst_mult_5_4_q  $ (!Xd_0__inst_mult_5_5_q ) ) + ( Xd_0__inst_mult_5_179  ) + ( Xd_0__inst_mult_5_178  ))
// Xd_0__inst_mult_5_182  = SHARE((Xd_0__inst_mult_5_4_q  & Xd_0__inst_mult_5_5_q ))

	.dataa(!Xd_0__inst_mult_5_4_q ),
	.datab(!Xd_0__inst_mult_5_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_178 ),
	.sharein(Xd_0__inst_mult_5_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_180 ),
	.cout(Xd_0__inst_mult_5_181 ),
	.shareout(Xd_0__inst_mult_5_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_70 (
// Equation(s):
// Xd_0__inst_mult_2_180  = SUM(( !Xd_0__inst_mult_2_4_q  $ (!Xd_0__inst_mult_2_5_q ) ) + ( Xd_0__inst_mult_2_179  ) + ( Xd_0__inst_mult_2_178  ))
// Xd_0__inst_mult_2_181  = CARRY(( !Xd_0__inst_mult_2_4_q  $ (!Xd_0__inst_mult_2_5_q ) ) + ( Xd_0__inst_mult_2_179  ) + ( Xd_0__inst_mult_2_178  ))
// Xd_0__inst_mult_2_182  = SHARE((Xd_0__inst_mult_2_4_q  & Xd_0__inst_mult_2_5_q ))

	.dataa(!Xd_0__inst_mult_2_4_q ),
	.datab(!Xd_0__inst_mult_2_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_178 ),
	.sharein(Xd_0__inst_mult_2_179 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_180 ),
	.cout(Xd_0__inst_mult_2_181 ),
	.shareout(Xd_0__inst_mult_2_182 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_72 (
// Equation(s):
// Xd_0__inst_mult_3_200  = SUM(( !Xd_0__inst_mult_3_4_q  $ (!Xd_0__inst_mult_3_5_q ) ) + ( Xd_0__inst_mult_3_198  ) + ( Xd_0__inst_mult_3_197  ))
// Xd_0__inst_mult_3_201  = CARRY(( !Xd_0__inst_mult_3_4_q  $ (!Xd_0__inst_mult_3_5_q ) ) + ( Xd_0__inst_mult_3_198  ) + ( Xd_0__inst_mult_3_197  ))
// Xd_0__inst_mult_3_202  = SHARE((Xd_0__inst_mult_3_4_q  & Xd_0__inst_mult_3_5_q ))

	.dataa(!Xd_0__inst_mult_3_4_q ),
	.datab(!Xd_0__inst_mult_3_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_197 ),
	.sharein(Xd_0__inst_mult_3_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_200 ),
	.cout(Xd_0__inst_mult_3_201 ),
	.shareout(Xd_0__inst_mult_3_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_68 (
// Equation(s):
// Xd_0__inst_mult_0_184  = SUM(( !Xd_0__inst_mult_0_4_q  $ (!Xd_0__inst_mult_0_5_q ) ) + ( Xd_0__inst_mult_0_182  ) + ( Xd_0__inst_mult_0_181  ))
// Xd_0__inst_mult_0_185  = CARRY(( !Xd_0__inst_mult_0_4_q  $ (!Xd_0__inst_mult_0_5_q ) ) + ( Xd_0__inst_mult_0_182  ) + ( Xd_0__inst_mult_0_181  ))
// Xd_0__inst_mult_0_186  = SHARE((Xd_0__inst_mult_0_4_q  & Xd_0__inst_mult_0_5_q ))

	.dataa(!Xd_0__inst_mult_0_4_q ),
	.datab(!Xd_0__inst_mult_0_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_181 ),
	.sharein(Xd_0__inst_mult_0_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_184 ),
	.cout(Xd_0__inst_mult_0_185 ),
	.shareout(Xd_0__inst_mult_0_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_71 (
// Equation(s):
// Xd_0__inst_mult_1_196  = SUM(( !Xd_0__inst_mult_1_4_q  $ (!Xd_0__inst_mult_1_5_q ) ) + ( Xd_0__inst_mult_1_194  ) + ( Xd_0__inst_mult_1_193  ))
// Xd_0__inst_mult_1_197  = CARRY(( !Xd_0__inst_mult_1_4_q  $ (!Xd_0__inst_mult_1_5_q ) ) + ( Xd_0__inst_mult_1_194  ) + ( Xd_0__inst_mult_1_193  ))
// Xd_0__inst_mult_1_198  = SHARE((Xd_0__inst_mult_1_4_q  & Xd_0__inst_mult_1_5_q ))

	.dataa(!Xd_0__inst_mult_1_4_q ),
	.datab(!Xd_0__inst_mult_1_5_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_193 ),
	.sharein(Xd_0__inst_mult_1_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_196 ),
	.cout(Xd_0__inst_mult_1_197 ),
	.shareout(Xd_0__inst_mult_1_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_71 (
// Equation(s):
// Xd_0__inst_mult_4_184  = SUM(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_182  ) + ( Xd_0__inst_mult_4_181  ))
// Xd_0__inst_mult_4_185  = CARRY(( !Xd_0__inst_mult_4_6_q  $ (!Xd_0__inst_mult_4_7_q ) ) + ( Xd_0__inst_mult_4_182  ) + ( Xd_0__inst_mult_4_181  ))
// Xd_0__inst_mult_4_186  = SHARE((Xd_0__inst_mult_4_6_q  & Xd_0__inst_mult_4_7_q ))

	.dataa(!Xd_0__inst_mult_4_6_q ),
	.datab(!Xd_0__inst_mult_4_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_181 ),
	.sharein(Xd_0__inst_mult_4_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_184 ),
	.cout(Xd_0__inst_mult_4_185 ),
	.shareout(Xd_0__inst_mult_4_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_71 (
// Equation(s):
// Xd_0__inst_mult_5_184  = SUM(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_182  ) + ( Xd_0__inst_mult_5_181  ))
// Xd_0__inst_mult_5_185  = CARRY(( !Xd_0__inst_mult_5_6_q  $ (!Xd_0__inst_mult_5_7_q ) ) + ( Xd_0__inst_mult_5_182  ) + ( Xd_0__inst_mult_5_181  ))
// Xd_0__inst_mult_5_186  = SHARE((Xd_0__inst_mult_5_6_q  & Xd_0__inst_mult_5_7_q ))

	.dataa(!Xd_0__inst_mult_5_6_q ),
	.datab(!Xd_0__inst_mult_5_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_181 ),
	.sharein(Xd_0__inst_mult_5_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_184 ),
	.cout(Xd_0__inst_mult_5_185 ),
	.shareout(Xd_0__inst_mult_5_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_71 (
// Equation(s):
// Xd_0__inst_mult_2_184  = SUM(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_182  ) + ( Xd_0__inst_mult_2_181  ))
// Xd_0__inst_mult_2_185  = CARRY(( !Xd_0__inst_mult_2_6_q  $ (!Xd_0__inst_mult_2_7_q ) ) + ( Xd_0__inst_mult_2_182  ) + ( Xd_0__inst_mult_2_181  ))
// Xd_0__inst_mult_2_186  = SHARE((Xd_0__inst_mult_2_6_q  & Xd_0__inst_mult_2_7_q ))

	.dataa(!Xd_0__inst_mult_2_6_q ),
	.datab(!Xd_0__inst_mult_2_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_181 ),
	.sharein(Xd_0__inst_mult_2_182 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_184 ),
	.cout(Xd_0__inst_mult_2_185 ),
	.shareout(Xd_0__inst_mult_2_186 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_73 (
// Equation(s):
// Xd_0__inst_mult_3_204  = SUM(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_202  ) + ( Xd_0__inst_mult_3_201  ))
// Xd_0__inst_mult_3_205  = CARRY(( !Xd_0__inst_mult_3_6_q  $ (!Xd_0__inst_mult_3_7_q ) ) + ( Xd_0__inst_mult_3_202  ) + ( Xd_0__inst_mult_3_201  ))
// Xd_0__inst_mult_3_206  = SHARE((Xd_0__inst_mult_3_6_q  & Xd_0__inst_mult_3_7_q ))

	.dataa(!Xd_0__inst_mult_3_6_q ),
	.datab(!Xd_0__inst_mult_3_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_201 ),
	.sharein(Xd_0__inst_mult_3_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_204 ),
	.cout(Xd_0__inst_mult_3_205 ),
	.shareout(Xd_0__inst_mult_3_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_69 (
// Equation(s):
// Xd_0__inst_mult_0_188  = SUM(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_186  ) + ( Xd_0__inst_mult_0_185  ))
// Xd_0__inst_mult_0_189  = CARRY(( !Xd_0__inst_mult_0_6_q  $ (!Xd_0__inst_mult_0_7_q ) ) + ( Xd_0__inst_mult_0_186  ) + ( Xd_0__inst_mult_0_185  ))
// Xd_0__inst_mult_0_190  = SHARE((Xd_0__inst_mult_0_6_q  & Xd_0__inst_mult_0_7_q ))

	.dataa(!Xd_0__inst_mult_0_6_q ),
	.datab(!Xd_0__inst_mult_0_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_185 ),
	.sharein(Xd_0__inst_mult_0_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_188 ),
	.cout(Xd_0__inst_mult_0_189 ),
	.shareout(Xd_0__inst_mult_0_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_72 (
// Equation(s):
// Xd_0__inst_mult_1_200  = SUM(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_198  ) + ( Xd_0__inst_mult_1_197  ))
// Xd_0__inst_mult_1_201  = CARRY(( !Xd_0__inst_mult_1_6_q  $ (!Xd_0__inst_mult_1_7_q ) ) + ( Xd_0__inst_mult_1_198  ) + ( Xd_0__inst_mult_1_197  ))
// Xd_0__inst_mult_1_202  = SHARE((Xd_0__inst_mult_1_6_q  & Xd_0__inst_mult_1_7_q ))

	.dataa(!Xd_0__inst_mult_1_6_q ),
	.datab(!Xd_0__inst_mult_1_7_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_197 ),
	.sharein(Xd_0__inst_mult_1_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_200 ),
	.cout(Xd_0__inst_mult_1_201 ),
	.shareout(Xd_0__inst_mult_1_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_72 (
// Equation(s):
// Xd_0__inst_mult_4_188  = SUM(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_186  ) + ( Xd_0__inst_mult_4_185  ))
// Xd_0__inst_mult_4_189  = CARRY(( !Xd_0__inst_mult_4_8_q  $ (!Xd_0__inst_mult_4_9_q ) ) + ( Xd_0__inst_mult_4_186  ) + ( Xd_0__inst_mult_4_185  ))
// Xd_0__inst_mult_4_190  = SHARE((Xd_0__inst_mult_4_8_q  & Xd_0__inst_mult_4_9_q ))

	.dataa(!Xd_0__inst_mult_4_8_q ),
	.datab(!Xd_0__inst_mult_4_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_185 ),
	.sharein(Xd_0__inst_mult_4_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_188 ),
	.cout(Xd_0__inst_mult_4_189 ),
	.shareout(Xd_0__inst_mult_4_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_72 (
// Equation(s):
// Xd_0__inst_mult_5_188  = SUM(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_186  ) + ( Xd_0__inst_mult_5_185  ))
// Xd_0__inst_mult_5_189  = CARRY(( !Xd_0__inst_mult_5_8_q  $ (!Xd_0__inst_mult_5_9_q ) ) + ( Xd_0__inst_mult_5_186  ) + ( Xd_0__inst_mult_5_185  ))
// Xd_0__inst_mult_5_190  = SHARE((Xd_0__inst_mult_5_8_q  & Xd_0__inst_mult_5_9_q ))

	.dataa(!Xd_0__inst_mult_5_8_q ),
	.datab(!Xd_0__inst_mult_5_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_185 ),
	.sharein(Xd_0__inst_mult_5_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_188 ),
	.cout(Xd_0__inst_mult_5_189 ),
	.shareout(Xd_0__inst_mult_5_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_72 (
// Equation(s):
// Xd_0__inst_mult_2_188  = SUM(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_186  ) + ( Xd_0__inst_mult_2_185  ))
// Xd_0__inst_mult_2_189  = CARRY(( !Xd_0__inst_mult_2_8_q  $ (!Xd_0__inst_mult_2_9_q ) ) + ( Xd_0__inst_mult_2_186  ) + ( Xd_0__inst_mult_2_185  ))
// Xd_0__inst_mult_2_190  = SHARE((Xd_0__inst_mult_2_8_q  & Xd_0__inst_mult_2_9_q ))

	.dataa(!Xd_0__inst_mult_2_8_q ),
	.datab(!Xd_0__inst_mult_2_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_185 ),
	.sharein(Xd_0__inst_mult_2_186 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_188 ),
	.cout(Xd_0__inst_mult_2_189 ),
	.shareout(Xd_0__inst_mult_2_190 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_74 (
// Equation(s):
// Xd_0__inst_mult_3_208  = SUM(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_206  ) + ( Xd_0__inst_mult_3_205  ))
// Xd_0__inst_mult_3_209  = CARRY(( !Xd_0__inst_mult_3_8_q  $ (!Xd_0__inst_mult_3_9_q ) ) + ( Xd_0__inst_mult_3_206  ) + ( Xd_0__inst_mult_3_205  ))
// Xd_0__inst_mult_3_210  = SHARE((Xd_0__inst_mult_3_8_q  & Xd_0__inst_mult_3_9_q ))

	.dataa(!Xd_0__inst_mult_3_8_q ),
	.datab(!Xd_0__inst_mult_3_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_205 ),
	.sharein(Xd_0__inst_mult_3_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_208 ),
	.cout(Xd_0__inst_mult_3_209 ),
	.shareout(Xd_0__inst_mult_3_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_70 (
// Equation(s):
// Xd_0__inst_mult_0_192  = SUM(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_190  ) + ( Xd_0__inst_mult_0_189  ))
// Xd_0__inst_mult_0_193  = CARRY(( !Xd_0__inst_mult_0_8_q  $ (!Xd_0__inst_mult_0_9_q ) ) + ( Xd_0__inst_mult_0_190  ) + ( Xd_0__inst_mult_0_189  ))
// Xd_0__inst_mult_0_194  = SHARE((Xd_0__inst_mult_0_8_q  & Xd_0__inst_mult_0_9_q ))

	.dataa(!Xd_0__inst_mult_0_8_q ),
	.datab(!Xd_0__inst_mult_0_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_189 ),
	.sharein(Xd_0__inst_mult_0_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_192 ),
	.cout(Xd_0__inst_mult_0_193 ),
	.shareout(Xd_0__inst_mult_0_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_73 (
// Equation(s):
// Xd_0__inst_mult_1_204  = SUM(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_202  ) + ( Xd_0__inst_mult_1_201  ))
// Xd_0__inst_mult_1_205  = CARRY(( !Xd_0__inst_mult_1_8_q  $ (!Xd_0__inst_mult_1_9_q ) ) + ( Xd_0__inst_mult_1_202  ) + ( Xd_0__inst_mult_1_201  ))
// Xd_0__inst_mult_1_206  = SHARE((Xd_0__inst_mult_1_8_q  & Xd_0__inst_mult_1_9_q ))

	.dataa(!Xd_0__inst_mult_1_8_q ),
	.datab(!Xd_0__inst_mult_1_9_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_201 ),
	.sharein(Xd_0__inst_mult_1_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_204 ),
	.cout(Xd_0__inst_mult_1_205 ),
	.shareout(Xd_0__inst_mult_1_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_73 (
// Equation(s):
// Xd_0__inst_mult_4_192  = SUM(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q ) ) + ( Xd_0__inst_mult_4_190  ) + ( Xd_0__inst_mult_4_189  ))
// Xd_0__inst_mult_4_193  = CARRY(( !Xd_0__inst_mult_4_10_q  $ (!Xd_0__inst_mult_4_11_q ) ) + ( Xd_0__inst_mult_4_190  ) + ( Xd_0__inst_mult_4_189  ))
// Xd_0__inst_mult_4_194  = SHARE((Xd_0__inst_mult_4_10_q  & Xd_0__inst_mult_4_11_q ))

	.dataa(!Xd_0__inst_mult_4_10_q ),
	.datab(!Xd_0__inst_mult_4_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_189 ),
	.sharein(Xd_0__inst_mult_4_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_192 ),
	.cout(Xd_0__inst_mult_4_193 ),
	.shareout(Xd_0__inst_mult_4_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_73 (
// Equation(s):
// Xd_0__inst_mult_5_192  = SUM(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q ) ) + ( Xd_0__inst_mult_5_190  ) + ( Xd_0__inst_mult_5_189  ))
// Xd_0__inst_mult_5_193  = CARRY(( !Xd_0__inst_mult_5_10_q  $ (!Xd_0__inst_mult_5_11_q ) ) + ( Xd_0__inst_mult_5_190  ) + ( Xd_0__inst_mult_5_189  ))
// Xd_0__inst_mult_5_194  = SHARE((Xd_0__inst_mult_5_10_q  & Xd_0__inst_mult_5_11_q ))

	.dataa(!Xd_0__inst_mult_5_10_q ),
	.datab(!Xd_0__inst_mult_5_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_189 ),
	.sharein(Xd_0__inst_mult_5_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_192 ),
	.cout(Xd_0__inst_mult_5_193 ),
	.shareout(Xd_0__inst_mult_5_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_73 (
// Equation(s):
// Xd_0__inst_mult_2_192  = SUM(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q ) ) + ( Xd_0__inst_mult_2_190  ) + ( Xd_0__inst_mult_2_189  ))
// Xd_0__inst_mult_2_193  = CARRY(( !Xd_0__inst_mult_2_10_q  $ (!Xd_0__inst_mult_2_11_q ) ) + ( Xd_0__inst_mult_2_190  ) + ( Xd_0__inst_mult_2_189  ))
// Xd_0__inst_mult_2_194  = SHARE((Xd_0__inst_mult_2_10_q  & Xd_0__inst_mult_2_11_q ))

	.dataa(!Xd_0__inst_mult_2_10_q ),
	.datab(!Xd_0__inst_mult_2_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_189 ),
	.sharein(Xd_0__inst_mult_2_190 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_192 ),
	.cout(Xd_0__inst_mult_2_193 ),
	.shareout(Xd_0__inst_mult_2_194 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_75 (
// Equation(s):
// Xd_0__inst_mult_3_212  = SUM(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q ) ) + ( Xd_0__inst_mult_3_210  ) + ( Xd_0__inst_mult_3_209  ))
// Xd_0__inst_mult_3_213  = CARRY(( !Xd_0__inst_mult_3_10_q  $ (!Xd_0__inst_mult_3_11_q ) ) + ( Xd_0__inst_mult_3_210  ) + ( Xd_0__inst_mult_3_209  ))
// Xd_0__inst_mult_3_214  = SHARE((Xd_0__inst_mult_3_10_q  & Xd_0__inst_mult_3_11_q ))

	.dataa(!Xd_0__inst_mult_3_10_q ),
	.datab(!Xd_0__inst_mult_3_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_209 ),
	.sharein(Xd_0__inst_mult_3_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_212 ),
	.cout(Xd_0__inst_mult_3_213 ),
	.shareout(Xd_0__inst_mult_3_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_71 (
// Equation(s):
// Xd_0__inst_mult_0_196  = SUM(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q ) ) + ( Xd_0__inst_mult_0_194  ) + ( Xd_0__inst_mult_0_193  ))
// Xd_0__inst_mult_0_197  = CARRY(( !Xd_0__inst_mult_0_10_q  $ (!Xd_0__inst_mult_0_11_q ) ) + ( Xd_0__inst_mult_0_194  ) + ( Xd_0__inst_mult_0_193  ))
// Xd_0__inst_mult_0_198  = SHARE((Xd_0__inst_mult_0_10_q  & Xd_0__inst_mult_0_11_q ))

	.dataa(!Xd_0__inst_mult_0_10_q ),
	.datab(!Xd_0__inst_mult_0_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_193 ),
	.sharein(Xd_0__inst_mult_0_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_196 ),
	.cout(Xd_0__inst_mult_0_197 ),
	.shareout(Xd_0__inst_mult_0_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_74 (
// Equation(s):
// Xd_0__inst_mult_1_208  = SUM(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q ) ) + ( Xd_0__inst_mult_1_206  ) + ( Xd_0__inst_mult_1_205  ))
// Xd_0__inst_mult_1_209  = CARRY(( !Xd_0__inst_mult_1_10_q  $ (!Xd_0__inst_mult_1_11_q ) ) + ( Xd_0__inst_mult_1_206  ) + ( Xd_0__inst_mult_1_205  ))
// Xd_0__inst_mult_1_210  = SHARE((Xd_0__inst_mult_1_10_q  & Xd_0__inst_mult_1_11_q ))

	.dataa(!Xd_0__inst_mult_1_10_q ),
	.datab(!Xd_0__inst_mult_1_11_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_205 ),
	.sharein(Xd_0__inst_mult_1_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_208 ),
	.cout(Xd_0__inst_mult_1_209 ),
	.shareout(Xd_0__inst_mult_1_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_74 (
// Equation(s):
// Xd_0__inst_mult_4_196  = SUM(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_194  ) + ( Xd_0__inst_mult_4_193  ))
// Xd_0__inst_mult_4_197  = CARRY(( !Xd_0__inst_mult_4_12_q  $ (!Xd_0__inst_mult_4_13_q ) ) + ( Xd_0__inst_mult_4_194  ) + ( Xd_0__inst_mult_4_193  ))
// Xd_0__inst_mult_4_198  = SHARE((Xd_0__inst_mult_4_12_q  & Xd_0__inst_mult_4_13_q ))

	.dataa(!Xd_0__inst_mult_4_12_q ),
	.datab(!Xd_0__inst_mult_4_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_193 ),
	.sharein(Xd_0__inst_mult_4_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_196 ),
	.cout(Xd_0__inst_mult_4_197 ),
	.shareout(Xd_0__inst_mult_4_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_74 (
// Equation(s):
// Xd_0__inst_mult_5_196  = SUM(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_194  ) + ( Xd_0__inst_mult_5_193  ))
// Xd_0__inst_mult_5_197  = CARRY(( !Xd_0__inst_mult_5_12_q  $ (!Xd_0__inst_mult_5_13_q ) ) + ( Xd_0__inst_mult_5_194  ) + ( Xd_0__inst_mult_5_193  ))
// Xd_0__inst_mult_5_198  = SHARE((Xd_0__inst_mult_5_12_q  & Xd_0__inst_mult_5_13_q ))

	.dataa(!Xd_0__inst_mult_5_12_q ),
	.datab(!Xd_0__inst_mult_5_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_193 ),
	.sharein(Xd_0__inst_mult_5_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_196 ),
	.cout(Xd_0__inst_mult_5_197 ),
	.shareout(Xd_0__inst_mult_5_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_74 (
// Equation(s):
// Xd_0__inst_mult_2_196  = SUM(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_194  ) + ( Xd_0__inst_mult_2_193  ))
// Xd_0__inst_mult_2_197  = CARRY(( !Xd_0__inst_mult_2_12_q  $ (!Xd_0__inst_mult_2_13_q ) ) + ( Xd_0__inst_mult_2_194  ) + ( Xd_0__inst_mult_2_193  ))
// Xd_0__inst_mult_2_198  = SHARE((Xd_0__inst_mult_2_12_q  & Xd_0__inst_mult_2_13_q ))

	.dataa(!Xd_0__inst_mult_2_12_q ),
	.datab(!Xd_0__inst_mult_2_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_193 ),
	.sharein(Xd_0__inst_mult_2_194 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_196 ),
	.cout(Xd_0__inst_mult_2_197 ),
	.shareout(Xd_0__inst_mult_2_198 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_76 (
// Equation(s):
// Xd_0__inst_mult_3_216  = SUM(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_214  ) + ( Xd_0__inst_mult_3_213  ))
// Xd_0__inst_mult_3_217  = CARRY(( !Xd_0__inst_mult_3_12_q  $ (!Xd_0__inst_mult_3_13_q ) ) + ( Xd_0__inst_mult_3_214  ) + ( Xd_0__inst_mult_3_213  ))
// Xd_0__inst_mult_3_218  = SHARE((Xd_0__inst_mult_3_12_q  & Xd_0__inst_mult_3_13_q ))

	.dataa(!Xd_0__inst_mult_3_12_q ),
	.datab(!Xd_0__inst_mult_3_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_213 ),
	.sharein(Xd_0__inst_mult_3_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_216 ),
	.cout(Xd_0__inst_mult_3_217 ),
	.shareout(Xd_0__inst_mult_3_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_72 (
// Equation(s):
// Xd_0__inst_mult_0_200  = SUM(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_198  ) + ( Xd_0__inst_mult_0_197  ))
// Xd_0__inst_mult_0_201  = CARRY(( !Xd_0__inst_mult_0_12_q  $ (!Xd_0__inst_mult_0_13_q ) ) + ( Xd_0__inst_mult_0_198  ) + ( Xd_0__inst_mult_0_197  ))
// Xd_0__inst_mult_0_202  = SHARE((Xd_0__inst_mult_0_12_q  & Xd_0__inst_mult_0_13_q ))

	.dataa(!Xd_0__inst_mult_0_12_q ),
	.datab(!Xd_0__inst_mult_0_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_197 ),
	.sharein(Xd_0__inst_mult_0_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_200 ),
	.cout(Xd_0__inst_mult_0_201 ),
	.shareout(Xd_0__inst_mult_0_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_75 (
// Equation(s):
// Xd_0__inst_mult_1_212  = SUM(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_210  ) + ( Xd_0__inst_mult_1_209  ))
// Xd_0__inst_mult_1_213  = CARRY(( !Xd_0__inst_mult_1_12_q  $ (!Xd_0__inst_mult_1_13_q ) ) + ( Xd_0__inst_mult_1_210  ) + ( Xd_0__inst_mult_1_209  ))
// Xd_0__inst_mult_1_214  = SHARE((Xd_0__inst_mult_1_12_q  & Xd_0__inst_mult_1_13_q ))

	.dataa(!Xd_0__inst_mult_1_12_q ),
	.datab(!Xd_0__inst_mult_1_13_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_209 ),
	.sharein(Xd_0__inst_mult_1_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_212 ),
	.cout(Xd_0__inst_mult_1_213 ),
	.shareout(Xd_0__inst_mult_1_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_75 (
// Equation(s):
// Xd_0__inst_mult_4_200  = SUM(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_198  ) + ( Xd_0__inst_mult_4_197  ))
// Xd_0__inst_mult_4_201  = CARRY(( !Xd_0__inst_mult_4_14_q  $ (!Xd_0__inst_mult_4_15_q ) ) + ( Xd_0__inst_mult_4_198  ) + ( Xd_0__inst_mult_4_197  ))
// Xd_0__inst_mult_4_202  = SHARE((Xd_0__inst_mult_4_14_q  & Xd_0__inst_mult_4_15_q ))

	.dataa(!Xd_0__inst_mult_4_14_q ),
	.datab(!Xd_0__inst_mult_4_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_197 ),
	.sharein(Xd_0__inst_mult_4_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_200 ),
	.cout(Xd_0__inst_mult_4_201 ),
	.shareout(Xd_0__inst_mult_4_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_75 (
// Equation(s):
// Xd_0__inst_mult_5_200  = SUM(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_198  ) + ( Xd_0__inst_mult_5_197  ))
// Xd_0__inst_mult_5_201  = CARRY(( !Xd_0__inst_mult_5_14_q  $ (!Xd_0__inst_mult_5_15_q ) ) + ( Xd_0__inst_mult_5_198  ) + ( Xd_0__inst_mult_5_197  ))
// Xd_0__inst_mult_5_202  = SHARE((Xd_0__inst_mult_5_14_q  & Xd_0__inst_mult_5_15_q ))

	.dataa(!Xd_0__inst_mult_5_14_q ),
	.datab(!Xd_0__inst_mult_5_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_197 ),
	.sharein(Xd_0__inst_mult_5_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_200 ),
	.cout(Xd_0__inst_mult_5_201 ),
	.shareout(Xd_0__inst_mult_5_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_75 (
// Equation(s):
// Xd_0__inst_mult_2_200  = SUM(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_198  ) + ( Xd_0__inst_mult_2_197  ))
// Xd_0__inst_mult_2_201  = CARRY(( !Xd_0__inst_mult_2_14_q  $ (!Xd_0__inst_mult_2_15_q ) ) + ( Xd_0__inst_mult_2_198  ) + ( Xd_0__inst_mult_2_197  ))
// Xd_0__inst_mult_2_202  = SHARE((Xd_0__inst_mult_2_14_q  & Xd_0__inst_mult_2_15_q ))

	.dataa(!Xd_0__inst_mult_2_14_q ),
	.datab(!Xd_0__inst_mult_2_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_197 ),
	.sharein(Xd_0__inst_mult_2_198 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_200 ),
	.cout(Xd_0__inst_mult_2_201 ),
	.shareout(Xd_0__inst_mult_2_202 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_77 (
// Equation(s):
// Xd_0__inst_mult_3_220  = SUM(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_218  ) + ( Xd_0__inst_mult_3_217  ))
// Xd_0__inst_mult_3_221  = CARRY(( !Xd_0__inst_mult_3_14_q  $ (!Xd_0__inst_mult_3_15_q ) ) + ( Xd_0__inst_mult_3_218  ) + ( Xd_0__inst_mult_3_217  ))
// Xd_0__inst_mult_3_222  = SHARE((Xd_0__inst_mult_3_14_q  & Xd_0__inst_mult_3_15_q ))

	.dataa(!Xd_0__inst_mult_3_14_q ),
	.datab(!Xd_0__inst_mult_3_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_217 ),
	.sharein(Xd_0__inst_mult_3_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_220 ),
	.cout(Xd_0__inst_mult_3_221 ),
	.shareout(Xd_0__inst_mult_3_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_73 (
// Equation(s):
// Xd_0__inst_mult_0_204  = SUM(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_202  ) + ( Xd_0__inst_mult_0_201  ))
// Xd_0__inst_mult_0_205  = CARRY(( !Xd_0__inst_mult_0_14_q  $ (!Xd_0__inst_mult_0_15_q ) ) + ( Xd_0__inst_mult_0_202  ) + ( Xd_0__inst_mult_0_201  ))
// Xd_0__inst_mult_0_206  = SHARE((Xd_0__inst_mult_0_14_q  & Xd_0__inst_mult_0_15_q ))

	.dataa(!Xd_0__inst_mult_0_14_q ),
	.datab(!Xd_0__inst_mult_0_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_201 ),
	.sharein(Xd_0__inst_mult_0_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_204 ),
	.cout(Xd_0__inst_mult_0_205 ),
	.shareout(Xd_0__inst_mult_0_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_76 (
// Equation(s):
// Xd_0__inst_mult_1_216  = SUM(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_214  ) + ( Xd_0__inst_mult_1_213  ))
// Xd_0__inst_mult_1_217  = CARRY(( !Xd_0__inst_mult_1_14_q  $ (!Xd_0__inst_mult_1_15_q ) ) + ( Xd_0__inst_mult_1_214  ) + ( Xd_0__inst_mult_1_213  ))
// Xd_0__inst_mult_1_218  = SHARE((Xd_0__inst_mult_1_14_q  & Xd_0__inst_mult_1_15_q ))

	.dataa(!Xd_0__inst_mult_1_14_q ),
	.datab(!Xd_0__inst_mult_1_15_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_213 ),
	.sharein(Xd_0__inst_mult_1_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_216 ),
	.cout(Xd_0__inst_mult_1_217 ),
	.shareout(Xd_0__inst_mult_1_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_76 (
// Equation(s):
// Xd_0__inst_mult_4_204  = SUM(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q ) ) + ( Xd_0__inst_mult_4_202  ) + ( Xd_0__inst_mult_4_201  ))
// Xd_0__inst_mult_4_205  = CARRY(( !Xd_0__inst_mult_4_16_q  $ (!Xd_0__inst_mult_4_17_q ) ) + ( Xd_0__inst_mult_4_202  ) + ( Xd_0__inst_mult_4_201  ))
// Xd_0__inst_mult_4_206  = SHARE((Xd_0__inst_mult_4_16_q  & Xd_0__inst_mult_4_17_q ))

	.dataa(!Xd_0__inst_mult_4_16_q ),
	.datab(!Xd_0__inst_mult_4_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_201 ),
	.sharein(Xd_0__inst_mult_4_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_204 ),
	.cout(Xd_0__inst_mult_4_205 ),
	.shareout(Xd_0__inst_mult_4_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_76 (
// Equation(s):
// Xd_0__inst_mult_5_204  = SUM(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q ) ) + ( Xd_0__inst_mult_5_202  ) + ( Xd_0__inst_mult_5_201  ))
// Xd_0__inst_mult_5_205  = CARRY(( !Xd_0__inst_mult_5_16_q  $ (!Xd_0__inst_mult_5_17_q ) ) + ( Xd_0__inst_mult_5_202  ) + ( Xd_0__inst_mult_5_201  ))
// Xd_0__inst_mult_5_206  = SHARE((Xd_0__inst_mult_5_16_q  & Xd_0__inst_mult_5_17_q ))

	.dataa(!Xd_0__inst_mult_5_16_q ),
	.datab(!Xd_0__inst_mult_5_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_201 ),
	.sharein(Xd_0__inst_mult_5_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_204 ),
	.cout(Xd_0__inst_mult_5_205 ),
	.shareout(Xd_0__inst_mult_5_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_76 (
// Equation(s):
// Xd_0__inst_mult_2_204  = SUM(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q ) ) + ( Xd_0__inst_mult_2_202  ) + ( Xd_0__inst_mult_2_201  ))
// Xd_0__inst_mult_2_205  = CARRY(( !Xd_0__inst_mult_2_16_q  $ (!Xd_0__inst_mult_2_17_q ) ) + ( Xd_0__inst_mult_2_202  ) + ( Xd_0__inst_mult_2_201  ))
// Xd_0__inst_mult_2_206  = SHARE((Xd_0__inst_mult_2_16_q  & Xd_0__inst_mult_2_17_q ))

	.dataa(!Xd_0__inst_mult_2_16_q ),
	.datab(!Xd_0__inst_mult_2_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_201 ),
	.sharein(Xd_0__inst_mult_2_202 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_204 ),
	.cout(Xd_0__inst_mult_2_205 ),
	.shareout(Xd_0__inst_mult_2_206 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_78 (
// Equation(s):
// Xd_0__inst_mult_3_224  = SUM(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q ) ) + ( Xd_0__inst_mult_3_222  ) + ( Xd_0__inst_mult_3_221  ))
// Xd_0__inst_mult_3_225  = CARRY(( !Xd_0__inst_mult_3_16_q  $ (!Xd_0__inst_mult_3_17_q ) ) + ( Xd_0__inst_mult_3_222  ) + ( Xd_0__inst_mult_3_221  ))
// Xd_0__inst_mult_3_226  = SHARE((Xd_0__inst_mult_3_16_q  & Xd_0__inst_mult_3_17_q ))

	.dataa(!Xd_0__inst_mult_3_16_q ),
	.datab(!Xd_0__inst_mult_3_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_221 ),
	.sharein(Xd_0__inst_mult_3_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_224 ),
	.cout(Xd_0__inst_mult_3_225 ),
	.shareout(Xd_0__inst_mult_3_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_74 (
// Equation(s):
// Xd_0__inst_mult_0_208  = SUM(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q ) ) + ( Xd_0__inst_mult_0_206  ) + ( Xd_0__inst_mult_0_205  ))
// Xd_0__inst_mult_0_209  = CARRY(( !Xd_0__inst_mult_0_16_q  $ (!Xd_0__inst_mult_0_17_q ) ) + ( Xd_0__inst_mult_0_206  ) + ( Xd_0__inst_mult_0_205  ))
// Xd_0__inst_mult_0_210  = SHARE((Xd_0__inst_mult_0_16_q  & Xd_0__inst_mult_0_17_q ))

	.dataa(!Xd_0__inst_mult_0_16_q ),
	.datab(!Xd_0__inst_mult_0_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_205 ),
	.sharein(Xd_0__inst_mult_0_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_208 ),
	.cout(Xd_0__inst_mult_0_209 ),
	.shareout(Xd_0__inst_mult_0_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_77 (
// Equation(s):
// Xd_0__inst_mult_1_220  = SUM(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q ) ) + ( Xd_0__inst_mult_1_218  ) + ( Xd_0__inst_mult_1_217  ))
// Xd_0__inst_mult_1_221  = CARRY(( !Xd_0__inst_mult_1_16_q  $ (!Xd_0__inst_mult_1_17_q ) ) + ( Xd_0__inst_mult_1_218  ) + ( Xd_0__inst_mult_1_217  ))
// Xd_0__inst_mult_1_222  = SHARE((Xd_0__inst_mult_1_16_q  & Xd_0__inst_mult_1_17_q ))

	.dataa(!Xd_0__inst_mult_1_16_q ),
	.datab(!Xd_0__inst_mult_1_17_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_217 ),
	.sharein(Xd_0__inst_mult_1_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_220 ),
	.cout(Xd_0__inst_mult_1_221 ),
	.shareout(Xd_0__inst_mult_1_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_77 (
// Equation(s):
// Xd_0__inst_mult_4_208  = SUM(( !Xd_0__inst_mult_4_18_q  $ (!Xd_0__inst_mult_4_19_q ) ) + ( Xd_0__inst_mult_4_206  ) + ( Xd_0__inst_mult_4_205  ))
// Xd_0__inst_mult_4_209  = CARRY(( !Xd_0__inst_mult_4_18_q  $ (!Xd_0__inst_mult_4_19_q ) ) + ( Xd_0__inst_mult_4_206  ) + ( Xd_0__inst_mult_4_205  ))
// Xd_0__inst_mult_4_210  = SHARE((Xd_0__inst_mult_4_18_q  & Xd_0__inst_mult_4_19_q ))

	.dataa(!Xd_0__inst_mult_4_18_q ),
	.datab(!Xd_0__inst_mult_4_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_205 ),
	.sharein(Xd_0__inst_mult_4_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_208 ),
	.cout(Xd_0__inst_mult_4_209 ),
	.shareout(Xd_0__inst_mult_4_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_77 (
// Equation(s):
// Xd_0__inst_mult_5_208  = SUM(( !Xd_0__inst_mult_5_18_q  $ (!Xd_0__inst_mult_5_19_q ) ) + ( Xd_0__inst_mult_5_206  ) + ( Xd_0__inst_mult_5_205  ))
// Xd_0__inst_mult_5_209  = CARRY(( !Xd_0__inst_mult_5_18_q  $ (!Xd_0__inst_mult_5_19_q ) ) + ( Xd_0__inst_mult_5_206  ) + ( Xd_0__inst_mult_5_205  ))
// Xd_0__inst_mult_5_210  = SHARE((Xd_0__inst_mult_5_18_q  & Xd_0__inst_mult_5_19_q ))

	.dataa(!Xd_0__inst_mult_5_18_q ),
	.datab(!Xd_0__inst_mult_5_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_205 ),
	.sharein(Xd_0__inst_mult_5_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_208 ),
	.cout(Xd_0__inst_mult_5_209 ),
	.shareout(Xd_0__inst_mult_5_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_77 (
// Equation(s):
// Xd_0__inst_mult_2_208  = SUM(( !Xd_0__inst_mult_2_18_q  $ (!Xd_0__inst_mult_2_19_q ) ) + ( Xd_0__inst_mult_2_206  ) + ( Xd_0__inst_mult_2_205  ))
// Xd_0__inst_mult_2_209  = CARRY(( !Xd_0__inst_mult_2_18_q  $ (!Xd_0__inst_mult_2_19_q ) ) + ( Xd_0__inst_mult_2_206  ) + ( Xd_0__inst_mult_2_205  ))
// Xd_0__inst_mult_2_210  = SHARE((Xd_0__inst_mult_2_18_q  & Xd_0__inst_mult_2_19_q ))

	.dataa(!Xd_0__inst_mult_2_18_q ),
	.datab(!Xd_0__inst_mult_2_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_205 ),
	.sharein(Xd_0__inst_mult_2_206 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_208 ),
	.cout(Xd_0__inst_mult_2_209 ),
	.shareout(Xd_0__inst_mult_2_210 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_79 (
// Equation(s):
// Xd_0__inst_mult_3_228  = SUM(( !Xd_0__inst_mult_3_18_q  $ (!Xd_0__inst_mult_3_19_q ) ) + ( Xd_0__inst_mult_3_226  ) + ( Xd_0__inst_mult_3_225  ))
// Xd_0__inst_mult_3_229  = CARRY(( !Xd_0__inst_mult_3_18_q  $ (!Xd_0__inst_mult_3_19_q ) ) + ( Xd_0__inst_mult_3_226  ) + ( Xd_0__inst_mult_3_225  ))
// Xd_0__inst_mult_3_230  = SHARE((Xd_0__inst_mult_3_18_q  & Xd_0__inst_mult_3_19_q ))

	.dataa(!Xd_0__inst_mult_3_18_q ),
	.datab(!Xd_0__inst_mult_3_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_225 ),
	.sharein(Xd_0__inst_mult_3_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_228 ),
	.cout(Xd_0__inst_mult_3_229 ),
	.shareout(Xd_0__inst_mult_3_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_75 (
// Equation(s):
// Xd_0__inst_mult_0_212  = SUM(( !Xd_0__inst_mult_0_18_q  $ (!Xd_0__inst_mult_0_19_q ) ) + ( Xd_0__inst_mult_0_210  ) + ( Xd_0__inst_mult_0_209  ))
// Xd_0__inst_mult_0_213  = CARRY(( !Xd_0__inst_mult_0_18_q  $ (!Xd_0__inst_mult_0_19_q ) ) + ( Xd_0__inst_mult_0_210  ) + ( Xd_0__inst_mult_0_209  ))
// Xd_0__inst_mult_0_214  = SHARE((Xd_0__inst_mult_0_18_q  & Xd_0__inst_mult_0_19_q ))

	.dataa(!Xd_0__inst_mult_0_18_q ),
	.datab(!Xd_0__inst_mult_0_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_209 ),
	.sharein(Xd_0__inst_mult_0_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_212 ),
	.cout(Xd_0__inst_mult_0_213 ),
	.shareout(Xd_0__inst_mult_0_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_78 (
// Equation(s):
// Xd_0__inst_mult_1_224  = SUM(( !Xd_0__inst_mult_1_18_q  $ (!Xd_0__inst_mult_1_19_q ) ) + ( Xd_0__inst_mult_1_222  ) + ( Xd_0__inst_mult_1_221  ))
// Xd_0__inst_mult_1_225  = CARRY(( !Xd_0__inst_mult_1_18_q  $ (!Xd_0__inst_mult_1_19_q ) ) + ( Xd_0__inst_mult_1_222  ) + ( Xd_0__inst_mult_1_221  ))
// Xd_0__inst_mult_1_226  = SHARE((Xd_0__inst_mult_1_18_q  & Xd_0__inst_mult_1_19_q ))

	.dataa(!Xd_0__inst_mult_1_18_q ),
	.datab(!Xd_0__inst_mult_1_19_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_221 ),
	.sharein(Xd_0__inst_mult_1_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_224 ),
	.cout(Xd_0__inst_mult_1_225 ),
	.shareout(Xd_0__inst_mult_1_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_78 (
// Equation(s):
// Xd_0__inst_mult_4_212  = SUM(( !Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q  $ (((Xd_0__inst_mult_4_22_q  & Xd_0__inst_mult_4_23_q )))) ) + ( Xd_0__inst_mult_4_210  ) + ( Xd_0__inst_mult_4_209  ))
// Xd_0__inst_mult_4_213  = CARRY(( !Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q  $ (((Xd_0__inst_mult_4_22_q  & Xd_0__inst_mult_4_23_q )))) ) + ( Xd_0__inst_mult_4_210  ) + ( Xd_0__inst_mult_4_209  ))
// Xd_0__inst_mult_4_214  = SHARE((Xd_0__inst_mult_4_22_q  & (Xd_0__inst_mult_4_23_q  & (!Xd_0__inst_mult_4_20_q  $ (!Xd_0__inst_mult_4_21_q )))))

	.dataa(!Xd_0__inst_mult_4_20_q ),
	.datab(!Xd_0__inst_mult_4_21_q ),
	.datac(!Xd_0__inst_mult_4_22_q ),
	.datad(!Xd_0__inst_mult_4_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_209 ),
	.sharein(Xd_0__inst_mult_4_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_212 ),
	.cout(Xd_0__inst_mult_4_213 ),
	.shareout(Xd_0__inst_mult_4_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_78 (
// Equation(s):
// Xd_0__inst_mult_5_212  = SUM(( !Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q  $ (((Xd_0__inst_mult_5_22_q  & Xd_0__inst_mult_5_23_q )))) ) + ( Xd_0__inst_mult_5_210  ) + ( Xd_0__inst_mult_5_209  ))
// Xd_0__inst_mult_5_213  = CARRY(( !Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q  $ (((Xd_0__inst_mult_5_22_q  & Xd_0__inst_mult_5_23_q )))) ) + ( Xd_0__inst_mult_5_210  ) + ( Xd_0__inst_mult_5_209  ))
// Xd_0__inst_mult_5_214  = SHARE((Xd_0__inst_mult_5_22_q  & (Xd_0__inst_mult_5_23_q  & (!Xd_0__inst_mult_5_20_q  $ (!Xd_0__inst_mult_5_21_q )))))

	.dataa(!Xd_0__inst_mult_5_20_q ),
	.datab(!Xd_0__inst_mult_5_21_q ),
	.datac(!Xd_0__inst_mult_5_22_q ),
	.datad(!Xd_0__inst_mult_5_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_209 ),
	.sharein(Xd_0__inst_mult_5_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_212 ),
	.cout(Xd_0__inst_mult_5_213 ),
	.shareout(Xd_0__inst_mult_5_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_78 (
// Equation(s):
// Xd_0__inst_mult_2_212  = SUM(( !Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q  $ (((Xd_0__inst_mult_2_22_q  & Xd_0__inst_mult_2_23_q )))) ) + ( Xd_0__inst_mult_2_210  ) + ( Xd_0__inst_mult_2_209  ))
// Xd_0__inst_mult_2_213  = CARRY(( !Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q  $ (((Xd_0__inst_mult_2_22_q  & Xd_0__inst_mult_2_23_q )))) ) + ( Xd_0__inst_mult_2_210  ) + ( Xd_0__inst_mult_2_209  ))
// Xd_0__inst_mult_2_214  = SHARE((Xd_0__inst_mult_2_22_q  & (Xd_0__inst_mult_2_23_q  & (!Xd_0__inst_mult_2_20_q  $ (!Xd_0__inst_mult_2_21_q )))))

	.dataa(!Xd_0__inst_mult_2_20_q ),
	.datab(!Xd_0__inst_mult_2_21_q ),
	.datac(!Xd_0__inst_mult_2_22_q ),
	.datad(!Xd_0__inst_mult_2_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_209 ),
	.sharein(Xd_0__inst_mult_2_210 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_212 ),
	.cout(Xd_0__inst_mult_2_213 ),
	.shareout(Xd_0__inst_mult_2_214 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_80 (
// Equation(s):
// Xd_0__inst_mult_3_232  = SUM(( !Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q  $ (((Xd_0__inst_mult_3_22_q  & Xd_0__inst_mult_3_23_q )))) ) + ( Xd_0__inst_mult_3_230  ) + ( Xd_0__inst_mult_3_229  ))
// Xd_0__inst_mult_3_233  = CARRY(( !Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q  $ (((Xd_0__inst_mult_3_22_q  & Xd_0__inst_mult_3_23_q )))) ) + ( Xd_0__inst_mult_3_230  ) + ( Xd_0__inst_mult_3_229  ))
// Xd_0__inst_mult_3_234  = SHARE((Xd_0__inst_mult_3_22_q  & (Xd_0__inst_mult_3_23_q  & (!Xd_0__inst_mult_3_20_q  $ (!Xd_0__inst_mult_3_21_q )))))

	.dataa(!Xd_0__inst_mult_3_20_q ),
	.datab(!Xd_0__inst_mult_3_21_q ),
	.datac(!Xd_0__inst_mult_3_22_q ),
	.datad(!Xd_0__inst_mult_3_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_229 ),
	.sharein(Xd_0__inst_mult_3_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_232 ),
	.cout(Xd_0__inst_mult_3_233 ),
	.shareout(Xd_0__inst_mult_3_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_76 (
// Equation(s):
// Xd_0__inst_mult_0_216  = SUM(( !Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q  $ (((Xd_0__inst_mult_0_22_q  & Xd_0__inst_mult_0_23_q )))) ) + ( Xd_0__inst_mult_0_214  ) + ( Xd_0__inst_mult_0_213  ))
// Xd_0__inst_mult_0_217  = CARRY(( !Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q  $ (((Xd_0__inst_mult_0_22_q  & Xd_0__inst_mult_0_23_q )))) ) + ( Xd_0__inst_mult_0_214  ) + ( Xd_0__inst_mult_0_213  ))
// Xd_0__inst_mult_0_218  = SHARE((Xd_0__inst_mult_0_22_q  & (Xd_0__inst_mult_0_23_q  & (!Xd_0__inst_mult_0_20_q  $ (!Xd_0__inst_mult_0_21_q )))))

	.dataa(!Xd_0__inst_mult_0_20_q ),
	.datab(!Xd_0__inst_mult_0_21_q ),
	.datac(!Xd_0__inst_mult_0_22_q ),
	.datad(!Xd_0__inst_mult_0_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_213 ),
	.sharein(Xd_0__inst_mult_0_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_216 ),
	.cout(Xd_0__inst_mult_0_217 ),
	.shareout(Xd_0__inst_mult_0_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_79 (
// Equation(s):
// Xd_0__inst_mult_1_228  = SUM(( !Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q  $ (((Xd_0__inst_mult_1_22_q  & Xd_0__inst_mult_1_23_q )))) ) + ( Xd_0__inst_mult_1_226  ) + ( Xd_0__inst_mult_1_225  ))
// Xd_0__inst_mult_1_229  = CARRY(( !Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q  $ (((Xd_0__inst_mult_1_22_q  & Xd_0__inst_mult_1_23_q )))) ) + ( Xd_0__inst_mult_1_226  ) + ( Xd_0__inst_mult_1_225  ))
// Xd_0__inst_mult_1_230  = SHARE((Xd_0__inst_mult_1_22_q  & (Xd_0__inst_mult_1_23_q  & (!Xd_0__inst_mult_1_20_q  $ (!Xd_0__inst_mult_1_21_q )))))

	.dataa(!Xd_0__inst_mult_1_20_q ),
	.datab(!Xd_0__inst_mult_1_21_q ),
	.datac(!Xd_0__inst_mult_1_22_q ),
	.datad(!Xd_0__inst_mult_1_23_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_225 ),
	.sharein(Xd_0__inst_mult_1_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_228 ),
	.cout(Xd_0__inst_mult_1_229 ),
	.shareout(Xd_0__inst_mult_1_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_79 (
// Equation(s):
// Xd_0__inst_mult_4_216  = SUM(( !Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q  $ (((Xd_0__inst_mult_4_20_q  & Xd_0__inst_mult_4_21_q )))) ) + ( Xd_0__inst_mult_4_214  ) + ( Xd_0__inst_mult_4_213  ))
// Xd_0__inst_mult_4_217  = CARRY(( !Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q  $ (((Xd_0__inst_mult_4_20_q  & Xd_0__inst_mult_4_21_q )))) ) + ( Xd_0__inst_mult_4_214  ) + ( Xd_0__inst_mult_4_213  ))
// Xd_0__inst_mult_4_218  = SHARE((Xd_0__inst_mult_4_20_q  & (Xd_0__inst_mult_4_21_q  & (!Xd_0__inst_mult_4_24_q  $ (!Xd_0__inst_mult_4_25_q )))))

	.dataa(!Xd_0__inst_mult_4_24_q ),
	.datab(!Xd_0__inst_mult_4_25_q ),
	.datac(!Xd_0__inst_mult_4_20_q ),
	.datad(!Xd_0__inst_mult_4_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_213 ),
	.sharein(Xd_0__inst_mult_4_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_216 ),
	.cout(Xd_0__inst_mult_4_217 ),
	.shareout(Xd_0__inst_mult_4_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_79 (
// Equation(s):
// Xd_0__inst_mult_5_216  = SUM(( !Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q  $ (((Xd_0__inst_mult_5_20_q  & Xd_0__inst_mult_5_21_q )))) ) + ( Xd_0__inst_mult_5_214  ) + ( Xd_0__inst_mult_5_213  ))
// Xd_0__inst_mult_5_217  = CARRY(( !Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q  $ (((Xd_0__inst_mult_5_20_q  & Xd_0__inst_mult_5_21_q )))) ) + ( Xd_0__inst_mult_5_214  ) + ( Xd_0__inst_mult_5_213  ))
// Xd_0__inst_mult_5_218  = SHARE((Xd_0__inst_mult_5_20_q  & (Xd_0__inst_mult_5_21_q  & (!Xd_0__inst_mult_5_24_q  $ (!Xd_0__inst_mult_5_25_q )))))

	.dataa(!Xd_0__inst_mult_5_24_q ),
	.datab(!Xd_0__inst_mult_5_25_q ),
	.datac(!Xd_0__inst_mult_5_20_q ),
	.datad(!Xd_0__inst_mult_5_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_213 ),
	.sharein(Xd_0__inst_mult_5_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_216 ),
	.cout(Xd_0__inst_mult_5_217 ),
	.shareout(Xd_0__inst_mult_5_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_79 (
// Equation(s):
// Xd_0__inst_mult_2_216  = SUM(( !Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q  $ (((Xd_0__inst_mult_2_20_q  & Xd_0__inst_mult_2_21_q )))) ) + ( Xd_0__inst_mult_2_214  ) + ( Xd_0__inst_mult_2_213  ))
// Xd_0__inst_mult_2_217  = CARRY(( !Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q  $ (((Xd_0__inst_mult_2_20_q  & Xd_0__inst_mult_2_21_q )))) ) + ( Xd_0__inst_mult_2_214  ) + ( Xd_0__inst_mult_2_213  ))
// Xd_0__inst_mult_2_218  = SHARE((Xd_0__inst_mult_2_20_q  & (Xd_0__inst_mult_2_21_q  & (!Xd_0__inst_mult_2_24_q  $ (!Xd_0__inst_mult_2_25_q )))))

	.dataa(!Xd_0__inst_mult_2_24_q ),
	.datab(!Xd_0__inst_mult_2_25_q ),
	.datac(!Xd_0__inst_mult_2_20_q ),
	.datad(!Xd_0__inst_mult_2_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_213 ),
	.sharein(Xd_0__inst_mult_2_214 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_216 ),
	.cout(Xd_0__inst_mult_2_217 ),
	.shareout(Xd_0__inst_mult_2_218 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_81 (
// Equation(s):
// Xd_0__inst_mult_3_236  = SUM(( !Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q  $ (((Xd_0__inst_mult_3_20_q  & Xd_0__inst_mult_3_21_q )))) ) + ( Xd_0__inst_mult_3_234  ) + ( Xd_0__inst_mult_3_233  ))
// Xd_0__inst_mult_3_237  = CARRY(( !Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q  $ (((Xd_0__inst_mult_3_20_q  & Xd_0__inst_mult_3_21_q )))) ) + ( Xd_0__inst_mult_3_234  ) + ( Xd_0__inst_mult_3_233  ))
// Xd_0__inst_mult_3_238  = SHARE((Xd_0__inst_mult_3_20_q  & (Xd_0__inst_mult_3_21_q  & (!Xd_0__inst_mult_3_24_q  $ (!Xd_0__inst_mult_3_25_q )))))

	.dataa(!Xd_0__inst_mult_3_24_q ),
	.datab(!Xd_0__inst_mult_3_25_q ),
	.datac(!Xd_0__inst_mult_3_20_q ),
	.datad(!Xd_0__inst_mult_3_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_233 ),
	.sharein(Xd_0__inst_mult_3_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_236 ),
	.cout(Xd_0__inst_mult_3_237 ),
	.shareout(Xd_0__inst_mult_3_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_77 (
// Equation(s):
// Xd_0__inst_mult_0_220  = SUM(( !Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q  $ (((Xd_0__inst_mult_0_20_q  & Xd_0__inst_mult_0_21_q )))) ) + ( Xd_0__inst_mult_0_218  ) + ( Xd_0__inst_mult_0_217  ))
// Xd_0__inst_mult_0_221  = CARRY(( !Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q  $ (((Xd_0__inst_mult_0_20_q  & Xd_0__inst_mult_0_21_q )))) ) + ( Xd_0__inst_mult_0_218  ) + ( Xd_0__inst_mult_0_217  ))
// Xd_0__inst_mult_0_222  = SHARE((Xd_0__inst_mult_0_20_q  & (Xd_0__inst_mult_0_21_q  & (!Xd_0__inst_mult_0_24_q  $ (!Xd_0__inst_mult_0_25_q )))))

	.dataa(!Xd_0__inst_mult_0_24_q ),
	.datab(!Xd_0__inst_mult_0_25_q ),
	.datac(!Xd_0__inst_mult_0_20_q ),
	.datad(!Xd_0__inst_mult_0_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_217 ),
	.sharein(Xd_0__inst_mult_0_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_220 ),
	.cout(Xd_0__inst_mult_0_221 ),
	.shareout(Xd_0__inst_mult_0_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_80 (
// Equation(s):
// Xd_0__inst_mult_1_232  = SUM(( !Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q  $ (((Xd_0__inst_mult_1_20_q  & Xd_0__inst_mult_1_21_q )))) ) + ( Xd_0__inst_mult_1_230  ) + ( Xd_0__inst_mult_1_229  ))
// Xd_0__inst_mult_1_233  = CARRY(( !Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q  $ (((Xd_0__inst_mult_1_20_q  & Xd_0__inst_mult_1_21_q )))) ) + ( Xd_0__inst_mult_1_230  ) + ( Xd_0__inst_mult_1_229  ))
// Xd_0__inst_mult_1_234  = SHARE((Xd_0__inst_mult_1_20_q  & (Xd_0__inst_mult_1_21_q  & (!Xd_0__inst_mult_1_24_q  $ (!Xd_0__inst_mult_1_25_q )))))

	.dataa(!Xd_0__inst_mult_1_24_q ),
	.datab(!Xd_0__inst_mult_1_25_q ),
	.datac(!Xd_0__inst_mult_1_20_q ),
	.datad(!Xd_0__inst_mult_1_21_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_229 ),
	.sharein(Xd_0__inst_mult_1_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_232 ),
	.cout(Xd_0__inst_mult_1_233 ),
	.shareout(Xd_0__inst_mult_1_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_80 (
// Equation(s):
// Xd_0__inst_mult_4_220  = SUM(( !Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q  $ (((Xd_0__inst_mult_4_24_q  & Xd_0__inst_mult_4_25_q )))) ) + ( Xd_0__inst_mult_4_218  ) + ( Xd_0__inst_mult_4_217  ))
// Xd_0__inst_mult_4_221  = CARRY(( !Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q  $ (((Xd_0__inst_mult_4_24_q  & Xd_0__inst_mult_4_25_q )))) ) + ( Xd_0__inst_mult_4_218  ) + ( Xd_0__inst_mult_4_217  ))
// Xd_0__inst_mult_4_222  = SHARE((Xd_0__inst_mult_4_24_q  & (Xd_0__inst_mult_4_25_q  & (!Xd_0__inst_mult_4_26_q  $ (!Xd_0__inst_mult_4_27_q )))))

	.dataa(!Xd_0__inst_mult_4_26_q ),
	.datab(!Xd_0__inst_mult_4_27_q ),
	.datac(!Xd_0__inst_mult_4_24_q ),
	.datad(!Xd_0__inst_mult_4_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_217 ),
	.sharein(Xd_0__inst_mult_4_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_220 ),
	.cout(Xd_0__inst_mult_4_221 ),
	.shareout(Xd_0__inst_mult_4_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_80 (
// Equation(s):
// Xd_0__inst_mult_5_220  = SUM(( !Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q  $ (((Xd_0__inst_mult_5_24_q  & Xd_0__inst_mult_5_25_q )))) ) + ( Xd_0__inst_mult_5_218  ) + ( Xd_0__inst_mult_5_217  ))
// Xd_0__inst_mult_5_221  = CARRY(( !Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q  $ (((Xd_0__inst_mult_5_24_q  & Xd_0__inst_mult_5_25_q )))) ) + ( Xd_0__inst_mult_5_218  ) + ( Xd_0__inst_mult_5_217  ))
// Xd_0__inst_mult_5_222  = SHARE((Xd_0__inst_mult_5_24_q  & (Xd_0__inst_mult_5_25_q  & (!Xd_0__inst_mult_5_26_q  $ (!Xd_0__inst_mult_5_27_q )))))

	.dataa(!Xd_0__inst_mult_5_26_q ),
	.datab(!Xd_0__inst_mult_5_27_q ),
	.datac(!Xd_0__inst_mult_5_24_q ),
	.datad(!Xd_0__inst_mult_5_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_217 ),
	.sharein(Xd_0__inst_mult_5_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_220 ),
	.cout(Xd_0__inst_mult_5_221 ),
	.shareout(Xd_0__inst_mult_5_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_80 (
// Equation(s):
// Xd_0__inst_mult_2_220  = SUM(( !Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q  $ (((Xd_0__inst_mult_2_24_q  & Xd_0__inst_mult_2_25_q )))) ) + ( Xd_0__inst_mult_2_218  ) + ( Xd_0__inst_mult_2_217  ))
// Xd_0__inst_mult_2_221  = CARRY(( !Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q  $ (((Xd_0__inst_mult_2_24_q  & Xd_0__inst_mult_2_25_q )))) ) + ( Xd_0__inst_mult_2_218  ) + ( Xd_0__inst_mult_2_217  ))
// Xd_0__inst_mult_2_222  = SHARE((Xd_0__inst_mult_2_24_q  & (Xd_0__inst_mult_2_25_q  & (!Xd_0__inst_mult_2_26_q  $ (!Xd_0__inst_mult_2_27_q )))))

	.dataa(!Xd_0__inst_mult_2_26_q ),
	.datab(!Xd_0__inst_mult_2_27_q ),
	.datac(!Xd_0__inst_mult_2_24_q ),
	.datad(!Xd_0__inst_mult_2_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_217 ),
	.sharein(Xd_0__inst_mult_2_218 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_220 ),
	.cout(Xd_0__inst_mult_2_221 ),
	.shareout(Xd_0__inst_mult_2_222 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_82 (
// Equation(s):
// Xd_0__inst_mult_3_240  = SUM(( !Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q  $ (((Xd_0__inst_mult_3_24_q  & Xd_0__inst_mult_3_25_q )))) ) + ( Xd_0__inst_mult_3_238  ) + ( Xd_0__inst_mult_3_237  ))
// Xd_0__inst_mult_3_241  = CARRY(( !Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q  $ (((Xd_0__inst_mult_3_24_q  & Xd_0__inst_mult_3_25_q )))) ) + ( Xd_0__inst_mult_3_238  ) + ( Xd_0__inst_mult_3_237  ))
// Xd_0__inst_mult_3_242  = SHARE((Xd_0__inst_mult_3_24_q  & (Xd_0__inst_mult_3_25_q  & (!Xd_0__inst_mult_3_26_q  $ (!Xd_0__inst_mult_3_27_q )))))

	.dataa(!Xd_0__inst_mult_3_26_q ),
	.datab(!Xd_0__inst_mult_3_27_q ),
	.datac(!Xd_0__inst_mult_3_24_q ),
	.datad(!Xd_0__inst_mult_3_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_237 ),
	.sharein(Xd_0__inst_mult_3_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_240 ),
	.cout(Xd_0__inst_mult_3_241 ),
	.shareout(Xd_0__inst_mult_3_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_78 (
// Equation(s):
// Xd_0__inst_mult_0_224  = SUM(( !Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q  $ (((Xd_0__inst_mult_0_24_q  & Xd_0__inst_mult_0_25_q )))) ) + ( Xd_0__inst_mult_0_222  ) + ( Xd_0__inst_mult_0_221  ))
// Xd_0__inst_mult_0_225  = CARRY(( !Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q  $ (((Xd_0__inst_mult_0_24_q  & Xd_0__inst_mult_0_25_q )))) ) + ( Xd_0__inst_mult_0_222  ) + ( Xd_0__inst_mult_0_221  ))
// Xd_0__inst_mult_0_226  = SHARE((Xd_0__inst_mult_0_24_q  & (Xd_0__inst_mult_0_25_q  & (!Xd_0__inst_mult_0_26_q  $ (!Xd_0__inst_mult_0_27_q )))))

	.dataa(!Xd_0__inst_mult_0_26_q ),
	.datab(!Xd_0__inst_mult_0_27_q ),
	.datac(!Xd_0__inst_mult_0_24_q ),
	.datad(!Xd_0__inst_mult_0_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_221 ),
	.sharein(Xd_0__inst_mult_0_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_224 ),
	.cout(Xd_0__inst_mult_0_225 ),
	.shareout(Xd_0__inst_mult_0_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_81 (
// Equation(s):
// Xd_0__inst_mult_1_236  = SUM(( !Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q  $ (((Xd_0__inst_mult_1_24_q  & Xd_0__inst_mult_1_25_q )))) ) + ( Xd_0__inst_mult_1_234  ) + ( Xd_0__inst_mult_1_233  ))
// Xd_0__inst_mult_1_237  = CARRY(( !Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q  $ (((Xd_0__inst_mult_1_24_q  & Xd_0__inst_mult_1_25_q )))) ) + ( Xd_0__inst_mult_1_234  ) + ( Xd_0__inst_mult_1_233  ))
// Xd_0__inst_mult_1_238  = SHARE((Xd_0__inst_mult_1_24_q  & (Xd_0__inst_mult_1_25_q  & (!Xd_0__inst_mult_1_26_q  $ (!Xd_0__inst_mult_1_27_q )))))

	.dataa(!Xd_0__inst_mult_1_26_q ),
	.datab(!Xd_0__inst_mult_1_27_q ),
	.datac(!Xd_0__inst_mult_1_24_q ),
	.datad(!Xd_0__inst_mult_1_25_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_233 ),
	.sharein(Xd_0__inst_mult_1_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_236 ),
	.cout(Xd_0__inst_mult_1_237 ),
	.shareout(Xd_0__inst_mult_1_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_81 (
// Equation(s):
// Xd_0__inst_mult_4_224  = SUM(( !Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q  $ (((Xd_0__inst_mult_4_26_q  & Xd_0__inst_mult_4_27_q )))) ) + ( Xd_0__inst_mult_4_222  ) + ( Xd_0__inst_mult_4_221  ))
// Xd_0__inst_mult_4_225  = CARRY(( !Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q  $ (((Xd_0__inst_mult_4_26_q  & Xd_0__inst_mult_4_27_q )))) ) + ( Xd_0__inst_mult_4_222  ) + ( Xd_0__inst_mult_4_221  ))
// Xd_0__inst_mult_4_226  = SHARE((Xd_0__inst_mult_4_26_q  & (Xd_0__inst_mult_4_27_q  & (!Xd_0__inst_mult_4_28_q  $ (!Xd_0__inst_mult_4_29_q )))))

	.dataa(!Xd_0__inst_mult_4_28_q ),
	.datab(!Xd_0__inst_mult_4_29_q ),
	.datac(!Xd_0__inst_mult_4_26_q ),
	.datad(!Xd_0__inst_mult_4_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_221 ),
	.sharein(Xd_0__inst_mult_4_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_224 ),
	.cout(Xd_0__inst_mult_4_225 ),
	.shareout(Xd_0__inst_mult_4_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_81 (
// Equation(s):
// Xd_0__inst_mult_5_224  = SUM(( !Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q  $ (((Xd_0__inst_mult_5_26_q  & Xd_0__inst_mult_5_27_q )))) ) + ( Xd_0__inst_mult_5_222  ) + ( Xd_0__inst_mult_5_221  ))
// Xd_0__inst_mult_5_225  = CARRY(( !Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q  $ (((Xd_0__inst_mult_5_26_q  & Xd_0__inst_mult_5_27_q )))) ) + ( Xd_0__inst_mult_5_222  ) + ( Xd_0__inst_mult_5_221  ))
// Xd_0__inst_mult_5_226  = SHARE((Xd_0__inst_mult_5_26_q  & (Xd_0__inst_mult_5_27_q  & (!Xd_0__inst_mult_5_28_q  $ (!Xd_0__inst_mult_5_29_q )))))

	.dataa(!Xd_0__inst_mult_5_28_q ),
	.datab(!Xd_0__inst_mult_5_29_q ),
	.datac(!Xd_0__inst_mult_5_26_q ),
	.datad(!Xd_0__inst_mult_5_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_221 ),
	.sharein(Xd_0__inst_mult_5_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_224 ),
	.cout(Xd_0__inst_mult_5_225 ),
	.shareout(Xd_0__inst_mult_5_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_81 (
// Equation(s):
// Xd_0__inst_mult_2_224  = SUM(( !Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q  $ (((Xd_0__inst_mult_2_26_q  & Xd_0__inst_mult_2_27_q )))) ) + ( Xd_0__inst_mult_2_222  ) + ( Xd_0__inst_mult_2_221  ))
// Xd_0__inst_mult_2_225  = CARRY(( !Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q  $ (((Xd_0__inst_mult_2_26_q  & Xd_0__inst_mult_2_27_q )))) ) + ( Xd_0__inst_mult_2_222  ) + ( Xd_0__inst_mult_2_221  ))
// Xd_0__inst_mult_2_226  = SHARE((Xd_0__inst_mult_2_26_q  & (Xd_0__inst_mult_2_27_q  & (!Xd_0__inst_mult_2_28_q  $ (!Xd_0__inst_mult_2_29_q )))))

	.dataa(!Xd_0__inst_mult_2_28_q ),
	.datab(!Xd_0__inst_mult_2_29_q ),
	.datac(!Xd_0__inst_mult_2_26_q ),
	.datad(!Xd_0__inst_mult_2_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_221 ),
	.sharein(Xd_0__inst_mult_2_222 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_224 ),
	.cout(Xd_0__inst_mult_2_225 ),
	.shareout(Xd_0__inst_mult_2_226 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_83 (
// Equation(s):
// Xd_0__inst_mult_3_244  = SUM(( !Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q  $ (((Xd_0__inst_mult_3_26_q  & Xd_0__inst_mult_3_27_q )))) ) + ( Xd_0__inst_mult_3_242  ) + ( Xd_0__inst_mult_3_241  ))
// Xd_0__inst_mult_3_245  = CARRY(( !Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q  $ (((Xd_0__inst_mult_3_26_q  & Xd_0__inst_mult_3_27_q )))) ) + ( Xd_0__inst_mult_3_242  ) + ( Xd_0__inst_mult_3_241  ))
// Xd_0__inst_mult_3_246  = SHARE((Xd_0__inst_mult_3_26_q  & (Xd_0__inst_mult_3_27_q  & (!Xd_0__inst_mult_3_28_q  $ (!Xd_0__inst_mult_3_29_q )))))

	.dataa(!Xd_0__inst_mult_3_28_q ),
	.datab(!Xd_0__inst_mult_3_29_q ),
	.datac(!Xd_0__inst_mult_3_26_q ),
	.datad(!Xd_0__inst_mult_3_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_241 ),
	.sharein(Xd_0__inst_mult_3_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_244 ),
	.cout(Xd_0__inst_mult_3_245 ),
	.shareout(Xd_0__inst_mult_3_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_79 (
// Equation(s):
// Xd_0__inst_mult_0_228  = SUM(( !Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q  $ (((Xd_0__inst_mult_0_26_q  & Xd_0__inst_mult_0_27_q )))) ) + ( Xd_0__inst_mult_0_226  ) + ( Xd_0__inst_mult_0_225  ))
// Xd_0__inst_mult_0_229  = CARRY(( !Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q  $ (((Xd_0__inst_mult_0_26_q  & Xd_0__inst_mult_0_27_q )))) ) + ( Xd_0__inst_mult_0_226  ) + ( Xd_0__inst_mult_0_225  ))
// Xd_0__inst_mult_0_230  = SHARE((Xd_0__inst_mult_0_26_q  & (Xd_0__inst_mult_0_27_q  & (!Xd_0__inst_mult_0_28_q  $ (!Xd_0__inst_mult_0_29_q )))))

	.dataa(!Xd_0__inst_mult_0_28_q ),
	.datab(!Xd_0__inst_mult_0_29_q ),
	.datac(!Xd_0__inst_mult_0_26_q ),
	.datad(!Xd_0__inst_mult_0_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_225 ),
	.sharein(Xd_0__inst_mult_0_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_228 ),
	.cout(Xd_0__inst_mult_0_229 ),
	.shareout(Xd_0__inst_mult_0_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_82 (
// Equation(s):
// Xd_0__inst_mult_1_240  = SUM(( !Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q  $ (((Xd_0__inst_mult_1_26_q  & Xd_0__inst_mult_1_27_q )))) ) + ( Xd_0__inst_mult_1_238  ) + ( Xd_0__inst_mult_1_237  ))
// Xd_0__inst_mult_1_241  = CARRY(( !Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q  $ (((Xd_0__inst_mult_1_26_q  & Xd_0__inst_mult_1_27_q )))) ) + ( Xd_0__inst_mult_1_238  ) + ( Xd_0__inst_mult_1_237  ))
// Xd_0__inst_mult_1_242  = SHARE((Xd_0__inst_mult_1_26_q  & (Xd_0__inst_mult_1_27_q  & (!Xd_0__inst_mult_1_28_q  $ (!Xd_0__inst_mult_1_29_q )))))

	.dataa(!Xd_0__inst_mult_1_28_q ),
	.datab(!Xd_0__inst_mult_1_29_q ),
	.datac(!Xd_0__inst_mult_1_26_q ),
	.datad(!Xd_0__inst_mult_1_27_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_237 ),
	.sharein(Xd_0__inst_mult_1_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_240 ),
	.cout(Xd_0__inst_mult_1_241 ),
	.shareout(Xd_0__inst_mult_1_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_82 (
// Equation(s):
// Xd_0__inst_mult_4_228  = SUM(( !Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q  $ (((Xd_0__inst_mult_4_28_q  & Xd_0__inst_mult_4_29_q )))) ) + ( Xd_0__inst_mult_4_226  ) + ( Xd_0__inst_mult_4_225  ))
// Xd_0__inst_mult_4_229  = CARRY(( !Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q  $ (((Xd_0__inst_mult_4_28_q  & Xd_0__inst_mult_4_29_q )))) ) + ( Xd_0__inst_mult_4_226  ) + ( Xd_0__inst_mult_4_225  ))
// Xd_0__inst_mult_4_230  = SHARE((Xd_0__inst_mult_4_28_q  & (Xd_0__inst_mult_4_29_q  & (!Xd_0__inst_mult_4_30_q  $ (!Xd_0__inst_mult_4_31_q )))))

	.dataa(!Xd_0__inst_mult_4_30_q ),
	.datab(!Xd_0__inst_mult_4_31_q ),
	.datac(!Xd_0__inst_mult_4_28_q ),
	.datad(!Xd_0__inst_mult_4_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_225 ),
	.sharein(Xd_0__inst_mult_4_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_228 ),
	.cout(Xd_0__inst_mult_4_229 ),
	.shareout(Xd_0__inst_mult_4_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_82 (
// Equation(s):
// Xd_0__inst_mult_5_228  = SUM(( !Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q  $ (((Xd_0__inst_mult_5_28_q  & Xd_0__inst_mult_5_29_q )))) ) + ( Xd_0__inst_mult_5_226  ) + ( Xd_0__inst_mult_5_225  ))
// Xd_0__inst_mult_5_229  = CARRY(( !Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q  $ (((Xd_0__inst_mult_5_28_q  & Xd_0__inst_mult_5_29_q )))) ) + ( Xd_0__inst_mult_5_226  ) + ( Xd_0__inst_mult_5_225  ))
// Xd_0__inst_mult_5_230  = SHARE((Xd_0__inst_mult_5_28_q  & (Xd_0__inst_mult_5_29_q  & (!Xd_0__inst_mult_5_30_q  $ (!Xd_0__inst_mult_5_31_q )))))

	.dataa(!Xd_0__inst_mult_5_30_q ),
	.datab(!Xd_0__inst_mult_5_31_q ),
	.datac(!Xd_0__inst_mult_5_28_q ),
	.datad(!Xd_0__inst_mult_5_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_225 ),
	.sharein(Xd_0__inst_mult_5_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_228 ),
	.cout(Xd_0__inst_mult_5_229 ),
	.shareout(Xd_0__inst_mult_5_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_82 (
// Equation(s):
// Xd_0__inst_mult_2_228  = SUM(( !Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q  $ (((Xd_0__inst_mult_2_28_q  & Xd_0__inst_mult_2_29_q )))) ) + ( Xd_0__inst_mult_2_226  ) + ( Xd_0__inst_mult_2_225  ))
// Xd_0__inst_mult_2_229  = CARRY(( !Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q  $ (((Xd_0__inst_mult_2_28_q  & Xd_0__inst_mult_2_29_q )))) ) + ( Xd_0__inst_mult_2_226  ) + ( Xd_0__inst_mult_2_225  ))
// Xd_0__inst_mult_2_230  = SHARE((Xd_0__inst_mult_2_28_q  & (Xd_0__inst_mult_2_29_q  & (!Xd_0__inst_mult_2_30_q  $ (!Xd_0__inst_mult_2_31_q )))))

	.dataa(!Xd_0__inst_mult_2_30_q ),
	.datab(!Xd_0__inst_mult_2_31_q ),
	.datac(!Xd_0__inst_mult_2_28_q ),
	.datad(!Xd_0__inst_mult_2_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_225 ),
	.sharein(Xd_0__inst_mult_2_226 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_228 ),
	.cout(Xd_0__inst_mult_2_229 ),
	.shareout(Xd_0__inst_mult_2_230 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_84 (
// Equation(s):
// Xd_0__inst_mult_3_248  = SUM(( !Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q  $ (((Xd_0__inst_mult_3_28_q  & Xd_0__inst_mult_3_29_q )))) ) + ( Xd_0__inst_mult_3_246  ) + ( Xd_0__inst_mult_3_245  ))
// Xd_0__inst_mult_3_249  = CARRY(( !Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q  $ (((Xd_0__inst_mult_3_28_q  & Xd_0__inst_mult_3_29_q )))) ) + ( Xd_0__inst_mult_3_246  ) + ( Xd_0__inst_mult_3_245  ))
// Xd_0__inst_mult_3_250  = SHARE((Xd_0__inst_mult_3_28_q  & (Xd_0__inst_mult_3_29_q  & (!Xd_0__inst_mult_3_30_q  $ (!Xd_0__inst_mult_3_31_q )))))

	.dataa(!Xd_0__inst_mult_3_30_q ),
	.datab(!Xd_0__inst_mult_3_31_q ),
	.datac(!Xd_0__inst_mult_3_28_q ),
	.datad(!Xd_0__inst_mult_3_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_245 ),
	.sharein(Xd_0__inst_mult_3_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_248 ),
	.cout(Xd_0__inst_mult_3_249 ),
	.shareout(Xd_0__inst_mult_3_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_80 (
// Equation(s):
// Xd_0__inst_mult_0_232  = SUM(( !Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q  $ (((Xd_0__inst_mult_0_28_q  & Xd_0__inst_mult_0_29_q )))) ) + ( Xd_0__inst_mult_0_230  ) + ( Xd_0__inst_mult_0_229  ))
// Xd_0__inst_mult_0_233  = CARRY(( !Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q  $ (((Xd_0__inst_mult_0_28_q  & Xd_0__inst_mult_0_29_q )))) ) + ( Xd_0__inst_mult_0_230  ) + ( Xd_0__inst_mult_0_229  ))
// Xd_0__inst_mult_0_234  = SHARE((Xd_0__inst_mult_0_28_q  & (Xd_0__inst_mult_0_29_q  & (!Xd_0__inst_mult_0_30_q  $ (!Xd_0__inst_mult_0_31_q )))))

	.dataa(!Xd_0__inst_mult_0_30_q ),
	.datab(!Xd_0__inst_mult_0_31_q ),
	.datac(!Xd_0__inst_mult_0_28_q ),
	.datad(!Xd_0__inst_mult_0_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_229 ),
	.sharein(Xd_0__inst_mult_0_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_232 ),
	.cout(Xd_0__inst_mult_0_233 ),
	.shareout(Xd_0__inst_mult_0_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_83 (
// Equation(s):
// Xd_0__inst_mult_1_244  = SUM(( !Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q  $ (((Xd_0__inst_mult_1_28_q  & Xd_0__inst_mult_1_29_q )))) ) + ( Xd_0__inst_mult_1_242  ) + ( Xd_0__inst_mult_1_241  ))
// Xd_0__inst_mult_1_245  = CARRY(( !Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q  $ (((Xd_0__inst_mult_1_28_q  & Xd_0__inst_mult_1_29_q )))) ) + ( Xd_0__inst_mult_1_242  ) + ( Xd_0__inst_mult_1_241  ))
// Xd_0__inst_mult_1_246  = SHARE((Xd_0__inst_mult_1_28_q  & (Xd_0__inst_mult_1_29_q  & (!Xd_0__inst_mult_1_30_q  $ (!Xd_0__inst_mult_1_31_q )))))

	.dataa(!Xd_0__inst_mult_1_30_q ),
	.datab(!Xd_0__inst_mult_1_31_q ),
	.datac(!Xd_0__inst_mult_1_28_q ),
	.datad(!Xd_0__inst_mult_1_29_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_241 ),
	.sharein(Xd_0__inst_mult_1_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_244 ),
	.cout(Xd_0__inst_mult_1_245 ),
	.shareout(Xd_0__inst_mult_1_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_83 (
// Equation(s):
// Xd_0__inst_mult_4_232  = SUM(( !Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q  $ (((Xd_0__inst_mult_4_30_q  & Xd_0__inst_mult_4_31_q )))) ) + ( Xd_0__inst_mult_4_230  ) + ( Xd_0__inst_mult_4_229  ))
// Xd_0__inst_mult_4_233  = CARRY(( !Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q  $ (((Xd_0__inst_mult_4_30_q  & Xd_0__inst_mult_4_31_q )))) ) + ( Xd_0__inst_mult_4_230  ) + ( Xd_0__inst_mult_4_229  ))
// Xd_0__inst_mult_4_234  = SHARE((Xd_0__inst_mult_4_30_q  & (Xd_0__inst_mult_4_31_q  & (!Xd_0__inst_mult_4_32_q  $ (!Xd_0__inst_mult_4_33_q )))))

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(!Xd_0__inst_mult_4_30_q ),
	.datad(!Xd_0__inst_mult_4_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_229 ),
	.sharein(Xd_0__inst_mult_4_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_232 ),
	.cout(Xd_0__inst_mult_4_233 ),
	.shareout(Xd_0__inst_mult_4_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_83 (
// Equation(s):
// Xd_0__inst_mult_5_232  = SUM(( !Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q  $ (((Xd_0__inst_mult_5_30_q  & Xd_0__inst_mult_5_31_q )))) ) + ( Xd_0__inst_mult_5_230  ) + ( Xd_0__inst_mult_5_229  ))
// Xd_0__inst_mult_5_233  = CARRY(( !Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q  $ (((Xd_0__inst_mult_5_30_q  & Xd_0__inst_mult_5_31_q )))) ) + ( Xd_0__inst_mult_5_230  ) + ( Xd_0__inst_mult_5_229  ))
// Xd_0__inst_mult_5_234  = SHARE((Xd_0__inst_mult_5_30_q  & (Xd_0__inst_mult_5_31_q  & (!Xd_0__inst_mult_5_32_q  $ (!Xd_0__inst_mult_5_33_q )))))

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(!Xd_0__inst_mult_5_30_q ),
	.datad(!Xd_0__inst_mult_5_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_229 ),
	.sharein(Xd_0__inst_mult_5_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_232 ),
	.cout(Xd_0__inst_mult_5_233 ),
	.shareout(Xd_0__inst_mult_5_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_83 (
// Equation(s):
// Xd_0__inst_mult_2_232  = SUM(( !Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q  $ (((Xd_0__inst_mult_2_30_q  & Xd_0__inst_mult_2_31_q )))) ) + ( Xd_0__inst_mult_2_230  ) + ( Xd_0__inst_mult_2_229  ))
// Xd_0__inst_mult_2_233  = CARRY(( !Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q  $ (((Xd_0__inst_mult_2_30_q  & Xd_0__inst_mult_2_31_q )))) ) + ( Xd_0__inst_mult_2_230  ) + ( Xd_0__inst_mult_2_229  ))
// Xd_0__inst_mult_2_234  = SHARE((Xd_0__inst_mult_2_30_q  & (Xd_0__inst_mult_2_31_q  & (!Xd_0__inst_mult_2_32_q  $ (!Xd_0__inst_mult_2_33_q )))))

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(!Xd_0__inst_mult_2_30_q ),
	.datad(!Xd_0__inst_mult_2_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_229 ),
	.sharein(Xd_0__inst_mult_2_230 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_232 ),
	.cout(Xd_0__inst_mult_2_233 ),
	.shareout(Xd_0__inst_mult_2_234 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_85 (
// Equation(s):
// Xd_0__inst_mult_3_252  = SUM(( !Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q  $ (((Xd_0__inst_mult_3_30_q  & Xd_0__inst_mult_3_31_q )))) ) + ( Xd_0__inst_mult_3_250  ) + ( Xd_0__inst_mult_3_249  ))
// Xd_0__inst_mult_3_253  = CARRY(( !Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q  $ (((Xd_0__inst_mult_3_30_q  & Xd_0__inst_mult_3_31_q )))) ) + ( Xd_0__inst_mult_3_250  ) + ( Xd_0__inst_mult_3_249  ))
// Xd_0__inst_mult_3_254  = SHARE((Xd_0__inst_mult_3_30_q  & (Xd_0__inst_mult_3_31_q  & (!Xd_0__inst_mult_3_32_q  $ (!Xd_0__inst_mult_3_33_q )))))

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(!Xd_0__inst_mult_3_30_q ),
	.datad(!Xd_0__inst_mult_3_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_249 ),
	.sharein(Xd_0__inst_mult_3_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_252 ),
	.cout(Xd_0__inst_mult_3_253 ),
	.shareout(Xd_0__inst_mult_3_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_81 (
// Equation(s):
// Xd_0__inst_mult_0_236  = SUM(( !Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q  $ (((Xd_0__inst_mult_0_30_q  & Xd_0__inst_mult_0_31_q )))) ) + ( Xd_0__inst_mult_0_234  ) + ( Xd_0__inst_mult_0_233  ))
// Xd_0__inst_mult_0_237  = CARRY(( !Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q  $ (((Xd_0__inst_mult_0_30_q  & Xd_0__inst_mult_0_31_q )))) ) + ( Xd_0__inst_mult_0_234  ) + ( Xd_0__inst_mult_0_233  ))
// Xd_0__inst_mult_0_238  = SHARE((Xd_0__inst_mult_0_30_q  & (Xd_0__inst_mult_0_31_q  & (!Xd_0__inst_mult_0_32_q  $ (!Xd_0__inst_mult_0_33_q )))))

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(!Xd_0__inst_mult_0_30_q ),
	.datad(!Xd_0__inst_mult_0_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_233 ),
	.sharein(Xd_0__inst_mult_0_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_236 ),
	.cout(Xd_0__inst_mult_0_237 ),
	.shareout(Xd_0__inst_mult_0_238 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000600006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_84 (
// Equation(s):
// Xd_0__inst_mult_1_248  = SUM(( !Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q  $ (((Xd_0__inst_mult_1_30_q  & Xd_0__inst_mult_1_31_q )))) ) + ( Xd_0__inst_mult_1_246  ) + ( Xd_0__inst_mult_1_245  ))
// Xd_0__inst_mult_1_249  = CARRY(( !Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q  $ (((Xd_0__inst_mult_1_30_q  & Xd_0__inst_mult_1_31_q )))) ) + ( Xd_0__inst_mult_1_246  ) + ( Xd_0__inst_mult_1_245  ))
// Xd_0__inst_mult_1_250  = SHARE((Xd_0__inst_mult_1_30_q  & (Xd_0__inst_mult_1_31_q  & (!Xd_0__inst_mult_1_32_q  $ (!Xd_0__inst_mult_1_33_q )))))

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(!Xd_0__inst_mult_1_30_q ),
	.datad(!Xd_0__inst_mult_1_31_q ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_245 ),
	.sharein(Xd_0__inst_mult_1_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_248 ),
	.cout(Xd_0__inst_mult_1_249 ),
	.shareout(Xd_0__inst_mult_1_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_84 (
// Equation(s):
// Xd_0__inst_mult_4_236  = SUM(( (Xd_0__inst_mult_4_32_q  & Xd_0__inst_mult_4_33_q ) ) + ( Xd_0__inst_mult_4_234  ) + ( Xd_0__inst_mult_4_233  ))

	.dataa(!Xd_0__inst_mult_4_32_q ),
	.datab(!Xd_0__inst_mult_4_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_233 ),
	.sharein(Xd_0__inst_mult_4_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_84 (
// Equation(s):
// Xd_0__inst_mult_5_236  = SUM(( (Xd_0__inst_mult_5_32_q  & Xd_0__inst_mult_5_33_q ) ) + ( Xd_0__inst_mult_5_234  ) + ( Xd_0__inst_mult_5_233  ))

	.dataa(!Xd_0__inst_mult_5_32_q ),
	.datab(!Xd_0__inst_mult_5_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_233 ),
	.sharein(Xd_0__inst_mult_5_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_84 (
// Equation(s):
// Xd_0__inst_mult_2_236  = SUM(( (Xd_0__inst_mult_2_32_q  & Xd_0__inst_mult_2_33_q ) ) + ( Xd_0__inst_mult_2_234  ) + ( Xd_0__inst_mult_2_233  ))

	.dataa(!Xd_0__inst_mult_2_32_q ),
	.datab(!Xd_0__inst_mult_2_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_233 ),
	.sharein(Xd_0__inst_mult_2_234 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_236 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_86 (
// Equation(s):
// Xd_0__inst_mult_3_256  = SUM(( (Xd_0__inst_mult_3_32_q  & Xd_0__inst_mult_3_33_q ) ) + ( Xd_0__inst_mult_3_254  ) + ( Xd_0__inst_mult_3_253  ))

	.dataa(!Xd_0__inst_mult_3_32_q ),
	.datab(!Xd_0__inst_mult_3_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_253 ),
	.sharein(Xd_0__inst_mult_3_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_256 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_82 (
// Equation(s):
// Xd_0__inst_mult_0_240  = SUM(( (Xd_0__inst_mult_0_32_q  & Xd_0__inst_mult_0_33_q ) ) + ( Xd_0__inst_mult_0_238  ) + ( Xd_0__inst_mult_0_237  ))

	.dataa(!Xd_0__inst_mult_0_32_q ),
	.datab(!Xd_0__inst_mult_0_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_237 ),
	.sharein(Xd_0__inst_mult_0_238 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_240 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_85 (
// Equation(s):
// Xd_0__inst_mult_1_252  = SUM(( (Xd_0__inst_mult_1_32_q  & Xd_0__inst_mult_1_33_q ) ) + ( Xd_0__inst_mult_1_250  ) + ( Xd_0__inst_mult_1_249  ))

	.dataa(!Xd_0__inst_mult_1_32_q ),
	.datab(!Xd_0__inst_mult_1_33_q ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_249 ),
	.sharein(Xd_0__inst_mult_1_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_252 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_85 (
// Equation(s):
// Xd_0__inst_mult_4_240  = SUM(( (din_a[48] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_241  = CARRY(( (din_a[48] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_242  = SHARE((din_a[48] & din_b[49]))

	.dataa(!din_a[48]),
	.datab(!din_b[48]),
	.datac(!din_b[49]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_240 ),
	.cout(Xd_0__inst_mult_4_241 ),
	.shareout(Xd_0__inst_mult_4_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_85 (
// Equation(s):
// Xd_0__inst_mult_5_240  = SUM(( (din_a[60] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_241  = CARRY(( (din_a[60] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_242  = SHARE((din_a[60] & din_b[61]))

	.dataa(!din_a[60]),
	.datab(!din_b[60]),
	.datac(!din_b[61]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_240 ),
	.cout(Xd_0__inst_mult_5_241 ),
	.shareout(Xd_0__inst_mult_5_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_9 (
// Equation(s):
// Xd_0__inst_i29_9_sumout  = SUM(( !din_a[59] $ (!din_b[59]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_10  = CARRY(( !din_a[59] $ (!din_b[59]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_i29_11  = SHARE(GND)

	.dataa(!din_a[59]),
	.datab(!din_b[59]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_i29_9_sumout ),
	.cout(Xd_0__inst_i29_10 ),
	.shareout(Xd_0__inst_i29_11 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_13 (
// Equation(s):
// Xd_0__inst_i29_13_sumout  = SUM(( !din_a[71] $ (!din_b[71]) ) + ( Xd_0__inst_i29_19  ) + ( Xd_0__inst_i29_18  ))
// Xd_0__inst_i29_14  = CARRY(( !din_a[71] $ (!din_b[71]) ) + ( Xd_0__inst_i29_19  ) + ( Xd_0__inst_i29_18  ))
// Xd_0__inst_i29_15  = SHARE(GND)

	.dataa(!din_a[71]),
	.datab(!din_b[71]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_18 ),
	.sharein(Xd_0__inst_i29_19 ),
	.combout(),
	.sumout(Xd_0__inst_i29_13_sumout ),
	.cout(Xd_0__inst_i29_14 ),
	.shareout(Xd_0__inst_i29_15 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_87 (
// Equation(s):
// Xd_0__inst_mult_3_260  = SUM(( GND ) + ( Xd_0__inst_mult_3_294  ) + ( Xd_0__inst_mult_3_293  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_293 ),
	.sharein(Xd_0__inst_mult_3_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_260 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_88 (
// Equation(s):
// Xd_0__inst_mult_3_264  = SUM(( !Xd_0__inst_mult_3_292  $ (((!din_b[39]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_298  ) + ( Xd_0__inst_mult_3_297  ))
// Xd_0__inst_mult_3_265  = CARRY(( !Xd_0__inst_mult_3_292  $ (((!din_b[39]) # (!din_a[46]))) ) + ( Xd_0__inst_mult_3_298  ) + ( Xd_0__inst_mult_3_297  ))
// Xd_0__inst_mult_3_266  = SHARE((din_b[39] & (din_a[46] & Xd_0__inst_mult_3_292 )))

	.dataa(!din_b[39]),
	.datab(!din_a[46]),
	.datac(!Xd_0__inst_mult_3_292 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_297 ),
	.sharein(Xd_0__inst_mult_3_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_264 ),
	.cout(Xd_0__inst_mult_3_265 ),
	.shareout(Xd_0__inst_mult_3_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_85 (
// Equation(s):
// Xd_0__inst_mult_2_240  = SUM(( (din_a[24] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_241  = CARRY(( (din_a[24] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_242  = SHARE((din_a[24] & din_b[25]))

	.dataa(!din_a[24]),
	.datab(!din_b[24]),
	.datac(!din_b[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_240 ),
	.cout(Xd_0__inst_mult_2_241 ),
	.shareout(Xd_0__inst_mult_2_242 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_89 (
// Equation(s):
// Xd_0__inst_mult_3_268  = SUM(( (din_a[36] & din_b[36]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_269  = CARRY(( (din_a[36] & din_b[36]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_270  = SHARE((din_a[36] & din_b[37]))

	.dataa(!din_a[36]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_268 ),
	.cout(Xd_0__inst_mult_3_269 ),
	.shareout(Xd_0__inst_mult_3_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_17 (
// Equation(s):
// Xd_0__inst_i29_17_sumout  = SUM(( !din_a[35] $ (!din_b[35]) ) + ( Xd_0__inst_i29_23  ) + ( Xd_0__inst_i29_22  ))
// Xd_0__inst_i29_18  = CARRY(( !din_a[35] $ (!din_b[35]) ) + ( Xd_0__inst_i29_23  ) + ( Xd_0__inst_i29_22  ))
// Xd_0__inst_i29_19  = SHARE(GND)

	.dataa(!din_a[35]),
	.datab(!din_b[35]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_22 ),
	.sharein(Xd_0__inst_i29_23 ),
	.combout(),
	.sumout(Xd_0__inst_i29_17_sumout ),
	.cout(Xd_0__inst_i29_18 ),
	.shareout(Xd_0__inst_i29_19 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_21 (
// Equation(s):
// Xd_0__inst_i29_21_sumout  = SUM(( !din_a[47] $ (!din_b[47]) ) + ( Xd_0__inst_i29_27  ) + ( Xd_0__inst_i29_26  ))
// Xd_0__inst_i29_22  = CARRY(( !din_a[47] $ (!din_b[47]) ) + ( Xd_0__inst_i29_27  ) + ( Xd_0__inst_i29_26  ))
// Xd_0__inst_i29_23  = SHARE(GND)

	.dataa(!din_a[47]),
	.datab(!din_b[47]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_26 ),
	.sharein(Xd_0__inst_i29_27 ),
	.combout(),
	.sumout(Xd_0__inst_i29_21_sumout ),
	.cout(Xd_0__inst_i29_22 ),
	.shareout(Xd_0__inst_i29_23 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_92 (
// Equation(s):
// Xd_0__inst_mult_6_268  = SUM(( GND ) + ( Xd_0__inst_mult_6_386  ) + ( Xd_0__inst_mult_6_385  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_385 ),
	.sharein(Xd_0__inst_mult_6_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_268 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_93 (
// Equation(s):
// Xd_0__inst_mult_6_272  = SUM(( !Xd_0__inst_mult_6_384  $ (((!din_b[75]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_346  ) + ( Xd_0__inst_mult_6_345  ))
// Xd_0__inst_mult_6_273  = CARRY(( !Xd_0__inst_mult_6_384  $ (((!din_b[75]) # (!din_a[82]))) ) + ( Xd_0__inst_mult_6_346  ) + ( Xd_0__inst_mult_6_345  ))
// Xd_0__inst_mult_6_274  = SHARE((din_b[75] & (din_a[82] & Xd_0__inst_mult_6_384 )))

	.dataa(!din_b[75]),
	.datab(!din_a[82]),
	.datac(!Xd_0__inst_mult_6_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_345 ),
	.sharein(Xd_0__inst_mult_6_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_272 ),
	.cout(Xd_0__inst_mult_6_273 ),
	.shareout(Xd_0__inst_mult_6_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_83 (
// Equation(s):
// Xd_0__inst_mult_0_244  = SUM(( (din_a[0] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_245  = CARRY(( (din_a[0] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_246  = SHARE((din_a[0] & din_b[1]))

	.dataa(!din_a[0]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_244 ),
	.cout(Xd_0__inst_mult_0_245 ),
	.shareout(Xd_0__inst_mult_0_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_25 (
// Equation(s):
// Xd_0__inst_i29_25_sumout  = SUM(( !din_a[11] $ (!din_b[11]) ) + ( Xd_0__inst_i29_31  ) + ( Xd_0__inst_i29_30  ))
// Xd_0__inst_i29_26  = CARRY(( !din_a[11] $ (!din_b[11]) ) + ( Xd_0__inst_i29_31  ) + ( Xd_0__inst_i29_30  ))
// Xd_0__inst_i29_27  = SHARE(GND)

	.dataa(!din_a[11]),
	.datab(!din_b[11]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_30 ),
	.sharein(Xd_0__inst_i29_31 ),
	.combout(),
	.sumout(Xd_0__inst_i29_25_sumout ),
	.cout(Xd_0__inst_i29_26 ),
	.shareout(Xd_0__inst_i29_27 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000006666),
	.shared_arith("on")
) Xd_0__inst_i29_29 (
// Equation(s):
// Xd_0__inst_i29_29_sumout  = SUM(( !din_a[23] $ (!din_b[23]) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_i29_30  = CARRY(( !din_a[23] $ (!din_b[23]) ) + ( Xd_0__inst_mult_3_41  ) + ( Xd_0__inst_mult_3_40  ))
// Xd_0__inst_i29_31  = SHARE(GND)

	.dataa(!din_a[23]),
	.datab(!din_b[23]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_40 ),
	.sharein(Xd_0__inst_mult_3_41 ),
	.combout(),
	.sumout(Xd_0__inst_i29_29_sumout ),
	.cout(Xd_0__inst_i29_30 ),
	.shareout(Xd_0__inst_i29_31 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_84 (
// Equation(s):
// Xd_0__inst_mult_0_248  = SUM(( GND ) + ( Xd_0__inst_mult_0_274  ) + ( Xd_0__inst_mult_0_273  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_273 ),
	.sharein(Xd_0__inst_mult_0_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_248 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_85 (
// Equation(s):
// Xd_0__inst_mult_0_252  = SUM(( !Xd_0__inst_mult_0_272  $ (((!din_b[3]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_278  ) + ( Xd_0__inst_mult_0_277  ))
// Xd_0__inst_mult_0_253  = CARRY(( !Xd_0__inst_mult_0_272  $ (((!din_b[3]) # (!din_a[10]))) ) + ( Xd_0__inst_mult_0_278  ) + ( Xd_0__inst_mult_0_277  ))
// Xd_0__inst_mult_0_254  = SHARE((din_b[3] & (din_a[10] & Xd_0__inst_mult_0_272 )))

	.dataa(!din_b[3]),
	.datab(!din_a[10]),
	.datac(!Xd_0__inst_mult_0_272 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_277 ),
	.sharein(Xd_0__inst_mult_0_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_252 ),
	.cout(Xd_0__inst_mult_0_253 ),
	.shareout(Xd_0__inst_mult_0_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_90 (
// Equation(s):
// Xd_0__inst_mult_3_272  = SUM(( (!din_a[43] & (((din_a[42] & din_b[45])))) # (din_a[43] & (!din_b[44] $ (((!din_a[42]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_3_302  ) + ( Xd_0__inst_mult_3_301  ))
// Xd_0__inst_mult_3_273  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[45])))) # (din_a[43] & (!din_b[44] $ (((!din_a[42]) # (!din_b[45]))))) ) + ( Xd_0__inst_mult_3_302  ) + ( Xd_0__inst_mult_3_301  ))
// Xd_0__inst_mult_3_274  = SHARE((din_a[43] & (din_b[44] & (din_a[42] & din_b[45]))))

	.dataa(!din_a[43]),
	.datab(!din_b[44]),
	.datac(!din_a[42]),
	.datad(!din_b[45]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_301 ),
	.sharein(Xd_0__inst_mult_3_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_272 ),
	.cout(Xd_0__inst_mult_3_273 ),
	.shareout(Xd_0__inst_mult_3_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_94 (
// Equation(s):
// Xd_0__inst_mult_7_276  = SUM(( (din_a[93] & din_b[88]) ) + ( Xd_0__inst_mult_7_390  ) + ( Xd_0__inst_mult_7_389  ))
// Xd_0__inst_mult_7_277  = CARRY(( (din_a[93] & din_b[88]) ) + ( Xd_0__inst_mult_7_390  ) + ( Xd_0__inst_mult_7_389  ))
// Xd_0__inst_mult_7_278  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[88]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_389 ),
	.sharein(Xd_0__inst_mult_7_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_276 ),
	.cout(Xd_0__inst_mult_7_277 ),
	.shareout(Xd_0__inst_mult_7_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_95 (
// Equation(s):
// Xd_0__inst_mult_7_280  = SUM(( !Xd_0__inst_mult_7_392  $ (!Xd_0__inst_mult_7_388  $ (((din_b[86] & din_a[94])))) ) + ( Xd_0__inst_mult_7_346  ) + ( Xd_0__inst_mult_7_345  ))
// Xd_0__inst_mult_7_281  = CARRY(( !Xd_0__inst_mult_7_392  $ (!Xd_0__inst_mult_7_388  $ (((din_b[86] & din_a[94])))) ) + ( Xd_0__inst_mult_7_346  ) + ( Xd_0__inst_mult_7_345  ))
// Xd_0__inst_mult_7_282  = SHARE((!Xd_0__inst_mult_7_392  & (Xd_0__inst_mult_7_388  & (din_b[86] & din_a[94]))) # (Xd_0__inst_mult_7_392  & (((din_b[86] & din_a[94])) # (Xd_0__inst_mult_7_388 ))))

	.dataa(!Xd_0__inst_mult_7_392 ),
	.datab(!Xd_0__inst_mult_7_388 ),
	.datac(!din_b[86]),
	.datad(!din_a[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_345 ),
	.sharein(Xd_0__inst_mult_7_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_280 ),
	.cout(Xd_0__inst_mult_7_281 ),
	.shareout(Xd_0__inst_mult_7_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_86 (
// Equation(s):
// Xd_0__inst_mult_4_244  = SUM(( (din_a[49] & din_b[48]) ) + ( Xd_0__inst_mult_4_242  ) + ( Xd_0__inst_mult_4_241  ))
// Xd_0__inst_mult_4_245  = CARRY(( (din_a[49] & din_b[48]) ) + ( Xd_0__inst_mult_4_242  ) + ( Xd_0__inst_mult_4_241  ))
// Xd_0__inst_mult_4_246  = SHARE((din_a[48] & din_b[50]))

	.dataa(!din_a[49]),
	.datab(!din_b[48]),
	.datac(!din_a[48]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_241 ),
	.sharein(Xd_0__inst_mult_4_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_244 ),
	.cout(Xd_0__inst_mult_4_245 ),
	.shareout(Xd_0__inst_mult_4_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_86 (
// Equation(s):
// Xd_0__inst_mult_5_244  = SUM(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_5_242  ) + ( Xd_0__inst_mult_5_241  ))
// Xd_0__inst_mult_5_245  = CARRY(( (din_a[61] & din_b[60]) ) + ( Xd_0__inst_mult_5_242  ) + ( Xd_0__inst_mult_5_241  ))
// Xd_0__inst_mult_5_246  = SHARE((din_a[60] & din_b[62]))

	.dataa(!din_a[61]),
	.datab(!din_b[60]),
	.datac(!din_a[60]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_241 ),
	.sharein(Xd_0__inst_mult_5_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_244 ),
	.cout(Xd_0__inst_mult_5_245 ),
	.shareout(Xd_0__inst_mult_5_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_86 (
// Equation(s):
// Xd_0__inst_mult_2_244  = SUM(( (din_a[25] & din_b[24]) ) + ( Xd_0__inst_mult_2_242  ) + ( Xd_0__inst_mult_2_241  ))
// Xd_0__inst_mult_2_245  = CARRY(( (din_a[25] & din_b[24]) ) + ( Xd_0__inst_mult_2_242  ) + ( Xd_0__inst_mult_2_241  ))
// Xd_0__inst_mult_2_246  = SHARE((din_a[24] & din_b[26]))

	.dataa(!din_a[25]),
	.datab(!din_b[24]),
	.datac(!din_a[24]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_241 ),
	.sharein(Xd_0__inst_mult_2_242 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_244 ),
	.cout(Xd_0__inst_mult_2_245 ),
	.shareout(Xd_0__inst_mult_2_246 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_91 (
// Equation(s):
// Xd_0__inst_mult_3_276  = SUM(( (din_a[37] & din_b[36]) ) + ( Xd_0__inst_mult_3_270  ) + ( Xd_0__inst_mult_3_269  ))
// Xd_0__inst_mult_3_277  = CARRY(( (din_a[37] & din_b[36]) ) + ( Xd_0__inst_mult_3_270  ) + ( Xd_0__inst_mult_3_269  ))
// Xd_0__inst_mult_3_278  = SHARE((din_a[36] & din_b[38]))

	.dataa(!din_a[37]),
	.datab(!din_b[36]),
	.datac(!din_a[36]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_269 ),
	.sharein(Xd_0__inst_mult_3_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_276 ),
	.cout(Xd_0__inst_mult_3_277 ),
	.shareout(Xd_0__inst_mult_3_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_86 (
// Equation(s):
// Xd_0__inst_mult_0_256  = SUM(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_246  ) + ( Xd_0__inst_mult_0_245  ))
// Xd_0__inst_mult_0_257  = CARRY(( (din_a[1] & din_b[0]) ) + ( Xd_0__inst_mult_0_246  ) + ( Xd_0__inst_mult_0_245  ))
// Xd_0__inst_mult_0_258  = SHARE((din_a[0] & din_b[2]))

	.dataa(!din_a[1]),
	.datab(!din_b[0]),
	.datac(!din_a[0]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_245 ),
	.sharein(Xd_0__inst_mult_0_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_256 ),
	.cout(Xd_0__inst_mult_0_257 ),
	.shareout(Xd_0__inst_mult_0_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_87 (
// Equation(s):
// Xd_0__inst_mult_4_248  = SUM(( (!din_a[49] & (((din_a[50] & din_b[48])))) # (din_a[49] & (!din_b[49] $ (((!din_a[50]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_246  ) + ( Xd_0__inst_mult_4_245  ))
// Xd_0__inst_mult_4_249  = CARRY(( (!din_a[49] & (((din_a[50] & din_b[48])))) # (din_a[49] & (!din_b[49] $ (((!din_a[50]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_246  ) + ( Xd_0__inst_mult_4_245  ))
// Xd_0__inst_mult_4_250  = SHARE((din_a[49] & (din_b[49] & (din_a[50] & din_b[48]))))

	.dataa(!din_a[49]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_245 ),
	.sharein(Xd_0__inst_mult_4_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_248 ),
	.cout(Xd_0__inst_mult_4_249 ),
	.shareout(Xd_0__inst_mult_4_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_87 (
// Equation(s):
// Xd_0__inst_mult_5_248  = SUM(( (!din_a[61] & (((din_a[62] & din_b[60])))) # (din_a[61] & (!din_b[61] $ (((!din_a[62]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_246  ) + ( Xd_0__inst_mult_5_245  ))
// Xd_0__inst_mult_5_249  = CARRY(( (!din_a[61] & (((din_a[62] & din_b[60])))) # (din_a[61] & (!din_b[61] $ (((!din_a[62]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_246  ) + ( Xd_0__inst_mult_5_245  ))
// Xd_0__inst_mult_5_250  = SHARE((din_a[61] & (din_b[61] & (din_a[62] & din_b[60]))))

	.dataa(!din_a[61]),
	.datab(!din_b[61]),
	.datac(!din_a[62]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_245 ),
	.sharein(Xd_0__inst_mult_5_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_248 ),
	.cout(Xd_0__inst_mult_5_249 ),
	.shareout(Xd_0__inst_mult_5_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_87 (
// Equation(s):
// Xd_0__inst_mult_2_248  = SUM(( (!din_a[25] & (((din_a[26] & din_b[24])))) # (din_a[25] & (!din_b[25] $ (((!din_a[26]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_246  ) + ( Xd_0__inst_mult_2_245  ))
// Xd_0__inst_mult_2_249  = CARRY(( (!din_a[25] & (((din_a[26] & din_b[24])))) # (din_a[25] & (!din_b[25] $ (((!din_a[26]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_246  ) + ( Xd_0__inst_mult_2_245  ))
// Xd_0__inst_mult_2_250  = SHARE((din_a[25] & (din_b[25] & (din_a[26] & din_b[24]))))

	.dataa(!din_a[25]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_245 ),
	.sharein(Xd_0__inst_mult_2_246 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_248 ),
	.cout(Xd_0__inst_mult_2_249 ),
	.shareout(Xd_0__inst_mult_2_250 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_92 (
// Equation(s):
// Xd_0__inst_mult_3_280  = SUM(( (!din_a[37] & (((din_a[38] & din_b[36])))) # (din_a[37] & (!din_b[37] $ (((!din_a[38]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_278  ) + ( Xd_0__inst_mult_3_277  ))
// Xd_0__inst_mult_3_281  = CARRY(( (!din_a[37] & (((din_a[38] & din_b[36])))) # (din_a[37] & (!din_b[37] $ (((!din_a[38]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_278  ) + ( Xd_0__inst_mult_3_277  ))
// Xd_0__inst_mult_3_282  = SHARE((din_a[37] & (din_b[37] & (din_a[38] & din_b[36]))))

	.dataa(!din_a[37]),
	.datab(!din_b[37]),
	.datac(!din_a[38]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_277 ),
	.sharein(Xd_0__inst_mult_3_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_280 ),
	.cout(Xd_0__inst_mult_3_281 ),
	.shareout(Xd_0__inst_mult_3_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_87 (
// Equation(s):
// Xd_0__inst_mult_0_260  = SUM(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_258  ) + ( Xd_0__inst_mult_0_257  ))
// Xd_0__inst_mult_0_261  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[0])))) # (din_a[1] & (!din_b[1] $ (((!din_a[2]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_258  ) + ( Xd_0__inst_mult_0_257  ))
// Xd_0__inst_mult_0_262  = SHARE((din_a[1] & (din_b[1] & (din_a[2] & din_b[0]))))

	.dataa(!din_a[1]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_257 ),
	.sharein(Xd_0__inst_mult_0_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_260 ),
	.cout(Xd_0__inst_mult_0_261 ),
	.shareout(Xd_0__inst_mult_0_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_88 (
// Equation(s):
// Xd_0__inst_mult_4_252  = SUM(( (din_a[48] & din_b[51]) ) + ( Xd_0__inst_mult_4_262  ) + ( Xd_0__inst_mult_4_261  ))
// Xd_0__inst_mult_4_253  = CARRY(( (din_a[48] & din_b[51]) ) + ( Xd_0__inst_mult_4_262  ) + ( Xd_0__inst_mult_4_261  ))
// Xd_0__inst_mult_4_254  = SHARE((din_a[48] & din_b[52]))

	.dataa(!din_a[48]),
	.datab(!din_b[51]),
	.datac(!din_b[52]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_261 ),
	.sharein(Xd_0__inst_mult_4_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_252 ),
	.cout(Xd_0__inst_mult_4_253 ),
	.shareout(Xd_0__inst_mult_4_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_88 (
// Equation(s):
// Xd_0__inst_mult_5_252  = SUM(( (din_a[60] & din_b[63]) ) + ( Xd_0__inst_mult_5_262  ) + ( Xd_0__inst_mult_5_261  ))
// Xd_0__inst_mult_5_253  = CARRY(( (din_a[60] & din_b[63]) ) + ( Xd_0__inst_mult_5_262  ) + ( Xd_0__inst_mult_5_261  ))
// Xd_0__inst_mult_5_254  = SHARE((din_a[60] & din_b[64]))

	.dataa(!din_a[60]),
	.datab(!din_b[63]),
	.datac(!din_b[64]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_261 ),
	.sharein(Xd_0__inst_mult_5_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_252 ),
	.cout(Xd_0__inst_mult_5_253 ),
	.shareout(Xd_0__inst_mult_5_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_88 (
// Equation(s):
// Xd_0__inst_mult_2_252  = SUM(( (din_a[24] & din_b[27]) ) + ( Xd_0__inst_mult_2_262  ) + ( Xd_0__inst_mult_2_261  ))
// Xd_0__inst_mult_2_253  = CARRY(( (din_a[24] & din_b[27]) ) + ( Xd_0__inst_mult_2_262  ) + ( Xd_0__inst_mult_2_261  ))
// Xd_0__inst_mult_2_254  = SHARE((din_a[24] & din_b[28]))

	.dataa(!din_a[24]),
	.datab(!din_b[27]),
	.datac(!din_b[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_261 ),
	.sharein(Xd_0__inst_mult_2_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_252 ),
	.cout(Xd_0__inst_mult_2_253 ),
	.shareout(Xd_0__inst_mult_2_254 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_93 (
// Equation(s):
// Xd_0__inst_mult_3_284  = SUM(( (din_a[36] & din_b[39]) ) + ( Xd_0__inst_mult_3_306  ) + ( Xd_0__inst_mult_3_305  ))
// Xd_0__inst_mult_3_285  = CARRY(( (din_a[36] & din_b[39]) ) + ( Xd_0__inst_mult_3_306  ) + ( Xd_0__inst_mult_3_305  ))
// Xd_0__inst_mult_3_286  = SHARE((din_a[36] & din_b[40]))

	.dataa(!din_a[36]),
	.datab(!din_b[39]),
	.datac(!din_b[40]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_305 ),
	.sharein(Xd_0__inst_mult_3_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_284 ),
	.cout(Xd_0__inst_mult_3_285 ),
	.shareout(Xd_0__inst_mult_3_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_88 (
// Equation(s):
// Xd_0__inst_mult_0_264  = SUM(( (din_a[0] & din_b[3]) ) + ( Xd_0__inst_mult_0_282  ) + ( Xd_0__inst_mult_0_281  ))
// Xd_0__inst_mult_0_265  = CARRY(( (din_a[0] & din_b[3]) ) + ( Xd_0__inst_mult_0_282  ) + ( Xd_0__inst_mult_0_281  ))
// Xd_0__inst_mult_0_266  = SHARE((din_a[0] & din_b[4]))

	.dataa(!din_a[0]),
	.datab(!din_b[3]),
	.datac(!din_b[4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_281 ),
	.sharein(Xd_0__inst_mult_0_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_264 ),
	.cout(Xd_0__inst_mult_0_265 ),
	.shareout(Xd_0__inst_mult_0_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_86 (
// Equation(s):
// Xd_0__inst_mult_1_256  = SUM(( (din_a[12] & din_b[15]) ) + ( Xd_0__inst_mult_1_266  ) + ( Xd_0__inst_mult_1_265  ))
// Xd_0__inst_mult_1_257  = CARRY(( (din_a[12] & din_b[15]) ) + ( Xd_0__inst_mult_1_266  ) + ( Xd_0__inst_mult_1_265  ))
// Xd_0__inst_mult_1_258  = SHARE((din_a[12] & din_b[16]))

	.dataa(!din_a[12]),
	.datab(!din_b[15]),
	.datac(!din_b[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_265 ),
	.sharein(Xd_0__inst_mult_1_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_256 ),
	.cout(Xd_0__inst_mult_1_257 ),
	.shareout(Xd_0__inst_mult_1_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_6_94 (
// Equation(s):
// Xd_0__inst_mult_6_277  = CARRY(( Xd_0__inst_mult_6_388  ) + ( Xd_0__inst_mult_6_394  ) + ( Xd_0__inst_mult_6_393  ))
// Xd_0__inst_mult_6_278  = SHARE((din_a[73] & din_b[74]))

	.dataa(!Xd_0__inst_mult_6_388 ),
	.datab(!din_a[73]),
	.datac(!din_b[74]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_393 ),
	.sharein(Xd_0__inst_mult_6_394 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_277 ),
	.shareout(Xd_0__inst_mult_6_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_7_96 (
// Equation(s):
// Xd_0__inst_mult_7_285  = CARRY(( Xd_0__inst_mult_7_396  ) + ( Xd_0__inst_mult_7_402  ) + ( Xd_0__inst_mult_7_401  ))
// Xd_0__inst_mult_7_286  = SHARE((din_a[85] & din_b[86]))

	.dataa(!Xd_0__inst_mult_7_396 ),
	.datab(!din_a[85]),
	.datac(!din_b[86]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_401 ),
	.sharein(Xd_0__inst_mult_7_402 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_285 ),
	.shareout(Xd_0__inst_mult_7_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_89 (
// Equation(s):
// Xd_0__inst_mult_4_256  = SUM(( !Xd_0__inst_mult_4_264  $ (!Xd_0__inst_mult_4_268 ) ) + ( Xd_0__inst_mult_4_254  ) + ( Xd_0__inst_mult_4_253  ))
// Xd_0__inst_mult_4_257  = CARRY(( !Xd_0__inst_mult_4_264  $ (!Xd_0__inst_mult_4_268 ) ) + ( Xd_0__inst_mult_4_254  ) + ( Xd_0__inst_mult_4_253  ))
// Xd_0__inst_mult_4_258  = SHARE((Xd_0__inst_mult_4_264  & Xd_0__inst_mult_4_268 ))

	.dataa(!Xd_0__inst_mult_4_264 ),
	.datab(!Xd_0__inst_mult_4_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_253 ),
	.sharein(Xd_0__inst_mult_4_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_256 ),
	.cout(Xd_0__inst_mult_4_257 ),
	.shareout(Xd_0__inst_mult_4_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_89 (
// Equation(s):
// Xd_0__inst_mult_5_256  = SUM(( !Xd_0__inst_mult_5_264  $ (!Xd_0__inst_mult_5_268 ) ) + ( Xd_0__inst_mult_5_254  ) + ( Xd_0__inst_mult_5_253  ))
// Xd_0__inst_mult_5_257  = CARRY(( !Xd_0__inst_mult_5_264  $ (!Xd_0__inst_mult_5_268 ) ) + ( Xd_0__inst_mult_5_254  ) + ( Xd_0__inst_mult_5_253  ))
// Xd_0__inst_mult_5_258  = SHARE((Xd_0__inst_mult_5_264  & Xd_0__inst_mult_5_268 ))

	.dataa(!Xd_0__inst_mult_5_264 ),
	.datab(!Xd_0__inst_mult_5_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_253 ),
	.sharein(Xd_0__inst_mult_5_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_256 ),
	.cout(Xd_0__inst_mult_5_257 ),
	.shareout(Xd_0__inst_mult_5_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_89 (
// Equation(s):
// Xd_0__inst_mult_2_256  = SUM(( !Xd_0__inst_mult_2_264  $ (!Xd_0__inst_mult_2_268 ) ) + ( Xd_0__inst_mult_2_254  ) + ( Xd_0__inst_mult_2_253  ))
// Xd_0__inst_mult_2_257  = CARRY(( !Xd_0__inst_mult_2_264  $ (!Xd_0__inst_mult_2_268 ) ) + ( Xd_0__inst_mult_2_254  ) + ( Xd_0__inst_mult_2_253  ))
// Xd_0__inst_mult_2_258  = SHARE((Xd_0__inst_mult_2_264  & Xd_0__inst_mult_2_268 ))

	.dataa(!Xd_0__inst_mult_2_264 ),
	.datab(!Xd_0__inst_mult_2_268 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_253 ),
	.sharein(Xd_0__inst_mult_2_254 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_256 ),
	.cout(Xd_0__inst_mult_2_257 ),
	.shareout(Xd_0__inst_mult_2_258 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_94 (
// Equation(s):
// Xd_0__inst_mult_3_288  = SUM(( !Xd_0__inst_mult_3_308  $ (!Xd_0__inst_mult_3_312 ) ) + ( Xd_0__inst_mult_3_286  ) + ( Xd_0__inst_mult_3_285  ))
// Xd_0__inst_mult_3_289  = CARRY(( !Xd_0__inst_mult_3_308  $ (!Xd_0__inst_mult_3_312 ) ) + ( Xd_0__inst_mult_3_286  ) + ( Xd_0__inst_mult_3_285  ))
// Xd_0__inst_mult_3_290  = SHARE((Xd_0__inst_mult_3_308  & Xd_0__inst_mult_3_312 ))

	.dataa(!Xd_0__inst_mult_3_308 ),
	.datab(!Xd_0__inst_mult_3_312 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_285 ),
	.sharein(Xd_0__inst_mult_3_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_288 ),
	.cout(Xd_0__inst_mult_3_289 ),
	.shareout(Xd_0__inst_mult_3_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_89 (
// Equation(s):
// Xd_0__inst_mult_0_268  = SUM(( !Xd_0__inst_mult_0_284  $ (!Xd_0__inst_mult_0_288 ) ) + ( Xd_0__inst_mult_0_266  ) + ( Xd_0__inst_mult_0_265  ))
// Xd_0__inst_mult_0_269  = CARRY(( !Xd_0__inst_mult_0_284  $ (!Xd_0__inst_mult_0_288 ) ) + ( Xd_0__inst_mult_0_266  ) + ( Xd_0__inst_mult_0_265  ))
// Xd_0__inst_mult_0_270  = SHARE((Xd_0__inst_mult_0_284  & Xd_0__inst_mult_0_288 ))

	.dataa(!Xd_0__inst_mult_0_284 ),
	.datab(!Xd_0__inst_mult_0_288 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_265 ),
	.sharein(Xd_0__inst_mult_0_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_268 ),
	.cout(Xd_0__inst_mult_0_269 ),
	.shareout(Xd_0__inst_mult_0_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_87 (
// Equation(s):
// Xd_0__inst_mult_1_260  = SUM(( !Xd_0__inst_mult_1_268  $ (!Xd_0__inst_mult_1_272 ) ) + ( Xd_0__inst_mult_1_258  ) + ( Xd_0__inst_mult_1_257  ))
// Xd_0__inst_mult_1_261  = CARRY(( !Xd_0__inst_mult_1_268  $ (!Xd_0__inst_mult_1_272 ) ) + ( Xd_0__inst_mult_1_258  ) + ( Xd_0__inst_mult_1_257  ))
// Xd_0__inst_mult_1_262  = SHARE((Xd_0__inst_mult_1_268  & Xd_0__inst_mult_1_272 ))

	.dataa(!Xd_0__inst_mult_1_268 ),
	.datab(!Xd_0__inst_mult_1_272 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_257 ),
	.sharein(Xd_0__inst_mult_1_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_260 ),
	.cout(Xd_0__inst_mult_1_261 ),
	.shareout(Xd_0__inst_mult_1_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_95 (
// Equation(s):
// Xd_0__inst_mult_6_280  = SUM(( (din_a[76] & din_b[72]) ) + ( Xd_0__inst_mult_6_390  ) + ( Xd_0__inst_mult_6_389  ))
// Xd_0__inst_mult_6_281  = CARRY(( (din_a[76] & din_b[72]) ) + ( Xd_0__inst_mult_6_390  ) + ( Xd_0__inst_mult_6_389  ))
// Xd_0__inst_mult_6_282  = SHARE((din_a[76] & din_b[73]))

	.dataa(!din_a[76]),
	.datab(!din_b[72]),
	.datac(!din_b[73]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_389 ),
	.sharein(Xd_0__inst_mult_6_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_280 ),
	.cout(Xd_0__inst_mult_6_281 ),
	.shareout(Xd_0__inst_mult_6_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_96 (
// Equation(s):
// Xd_0__inst_mult_6_284  = SUM(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_6_398  ) + ( Xd_0__inst_mult_6_397  ))
// Xd_0__inst_mult_6_285  = CARRY(( (din_a[73] & din_b[75]) ) + ( Xd_0__inst_mult_6_398  ) + ( Xd_0__inst_mult_6_397  ))
// Xd_0__inst_mult_6_286  = SHARE((din_b[75] & din_a[74]))

	.dataa(!din_a[73]),
	.datab(!din_b[75]),
	.datac(!din_a[74]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_397 ),
	.sharein(Xd_0__inst_mult_6_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_284 ),
	.cout(Xd_0__inst_mult_6_285 ),
	.shareout(Xd_0__inst_mult_6_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_97 (
// Equation(s):
// Xd_0__inst_mult_7_288  = SUM(( (din_a[88] & din_b[84]) ) + ( Xd_0__inst_mult_7_398  ) + ( Xd_0__inst_mult_7_397  ))
// Xd_0__inst_mult_7_289  = CARRY(( (din_a[88] & din_b[84]) ) + ( Xd_0__inst_mult_7_398  ) + ( Xd_0__inst_mult_7_397  ))
// Xd_0__inst_mult_7_290  = SHARE((din_a[88] & din_b[85]))

	.dataa(!din_a[88]),
	.datab(!din_b[84]),
	.datac(!din_b[85]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_397 ),
	.sharein(Xd_0__inst_mult_7_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_288 ),
	.cout(Xd_0__inst_mult_7_289 ),
	.shareout(Xd_0__inst_mult_7_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_98 (
// Equation(s):
// Xd_0__inst_mult_7_292  = SUM(( (din_a[85] & din_b[87]) ) + ( Xd_0__inst_mult_7_406  ) + ( Xd_0__inst_mult_7_405  ))
// Xd_0__inst_mult_7_293  = CARRY(( (din_a[85] & din_b[87]) ) + ( Xd_0__inst_mult_7_406  ) + ( Xd_0__inst_mult_7_405  ))
// Xd_0__inst_mult_7_294  = SHARE((din_b[87] & din_a[86]))

	.dataa(!din_a[85]),
	.datab(!din_b[87]),
	.datac(!din_a[86]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_405 ),
	.sharein(Xd_0__inst_mult_7_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_292 ),
	.cout(Xd_0__inst_mult_7_293 ),
	.shareout(Xd_0__inst_mult_7_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_35 (
// Equation(s):
// Xd_0__inst_mult_2_35_sumout  = SUM(( (din_a[34] & din_b[32]) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_2_36  = CARRY(( (din_a[34] & din_b[32]) ) + ( Xd_0__inst_mult_5_37  ) + ( Xd_0__inst_mult_5_36  ))
// Xd_0__inst_mult_2_37  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_36 ),
	.sharein(Xd_0__inst_mult_5_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_35_sumout ),
	.cout(Xd_0__inst_mult_2_36 ),
	.shareout(Xd_0__inst_mult_2_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_35 (
// Equation(s):
// Xd_0__inst_mult_0_35_sumout  = SUM(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_49  ) + ( Xd_0__inst_mult_1_48  ))
// Xd_0__inst_mult_0_36  = CARRY(( (din_a[10] & din_b[8]) ) + ( Xd_0__inst_mult_1_49  ) + ( Xd_0__inst_mult_1_48  ))
// Xd_0__inst_mult_0_37  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_48 ),
	.sharein(Xd_0__inst_mult_1_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_35_sumout ),
	.cout(Xd_0__inst_mult_0_36 ),
	.shareout(Xd_0__inst_mult_0_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_39 (
// Equation(s):
// Xd_0__inst_mult_2_39_sumout  = SUM(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_2_40  = CARRY(( (din_a[34] & din_b[33]) ) + ( Xd_0__inst_mult_5_41  ) + ( Xd_0__inst_mult_5_40  ))
// Xd_0__inst_mult_2_41  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[33]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_40 ),
	.sharein(Xd_0__inst_mult_5_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_39_sumout ),
	.cout(Xd_0__inst_mult_2_40 ),
	.shareout(Xd_0__inst_mult_2_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_35 (
// Equation(s):
// Xd_0__inst_mult_1_35_sumout  = SUM(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_0_41  ) + ( Xd_0__inst_mult_0_40  ))
// Xd_0__inst_mult_1_36  = CARRY(( (din_a[22] & din_b[21]) ) + ( Xd_0__inst_mult_0_41  ) + ( Xd_0__inst_mult_0_40  ))
// Xd_0__inst_mult_1_37  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[21]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_40 ),
	.sharein(Xd_0__inst_mult_0_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_35_sumout ),
	.cout(Xd_0__inst_mult_1_36 ),
	.shareout(Xd_0__inst_mult_1_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_43 (
// Equation(s):
// Xd_0__inst_mult_2_43_sumout  = SUM(( (din_a[34] & din_b[34]) ) + ( Xd_0__inst_mult_5_45  ) + ( Xd_0__inst_mult_5_44  ))
// Xd_0__inst_mult_2_44  = CARRY(( (din_a[34] & din_b[34]) ) + ( Xd_0__inst_mult_5_45  ) + ( Xd_0__inst_mult_5_44  ))
// Xd_0__inst_mult_2_45  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_44 ),
	.sharein(Xd_0__inst_mult_5_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_43_sumout ),
	.cout(Xd_0__inst_mult_2_44 ),
	.shareout(Xd_0__inst_mult_2_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_39 (
// Equation(s):
// Xd_0__inst_mult_1_39_sumout  = SUM(( (din_a[22] & din_b[22]) ) + ( Xd_0__inst_mult_0_45  ) + ( Xd_0__inst_mult_0_44  ))
// Xd_0__inst_mult_1_40  = CARRY(( (din_a[22] & din_b[22]) ) + ( Xd_0__inst_mult_0_45  ) + ( Xd_0__inst_mult_0_44  ))
// Xd_0__inst_mult_1_41  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_44 ),
	.sharein(Xd_0__inst_mult_0_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_39_sumout ),
	.cout(Xd_0__inst_mult_1_40 ),
	.shareout(Xd_0__inst_mult_1_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_97 (
// Equation(s):
// Xd_0__inst_mult_6_288  = SUM(( !Xd_0__inst_mult_6_400  $ (!Xd_0__inst_mult_6_404  $ (((din_b[76] & din_a[73])))) ) + ( Xd_0__inst_mult_6_266  ) + ( Xd_0__inst_mult_6_265  ))
// Xd_0__inst_mult_6_289  = CARRY(( !Xd_0__inst_mult_6_400  $ (!Xd_0__inst_mult_6_404  $ (((din_b[76] & din_a[73])))) ) + ( Xd_0__inst_mult_6_266  ) + ( Xd_0__inst_mult_6_265  ))
// Xd_0__inst_mult_6_290  = SHARE((!Xd_0__inst_mult_6_400  & (Xd_0__inst_mult_6_404  & (din_b[76] & din_a[73]))) # (Xd_0__inst_mult_6_400  & (((din_b[76] & din_a[73])) # (Xd_0__inst_mult_6_404 ))))

	.dataa(!Xd_0__inst_mult_6_400 ),
	.datab(!Xd_0__inst_mult_6_404 ),
	.datac(!din_b[76]),
	.datad(!din_a[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_265 ),
	.sharein(Xd_0__inst_mult_6_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_288 ),
	.cout(Xd_0__inst_mult_6_289 ),
	.shareout(Xd_0__inst_mult_6_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_98 (
// Equation(s):
// Xd_0__inst_mult_6_292  = SUM(( (din_a[72] & din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_293  = CARRY(( (din_a[72] & din_b[77]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_294  = SHARE((din_a[72] & din_b[78]))

	.dataa(!din_a[72]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_292 ),
	.cout(Xd_0__inst_mult_6_293 ),
	.shareout(Xd_0__inst_mult_6_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_43 (
// Equation(s):
// Xd_0__inst_mult_1_43_sumout  = SUM(( (din_a[21] & din_b[12]) ) + ( Xd_0__inst_mult_0_49  ) + ( Xd_0__inst_mult_0_48  ))
// Xd_0__inst_mult_1_44  = CARRY(( (din_a[21] & din_b[12]) ) + ( Xd_0__inst_mult_0_49  ) + ( Xd_0__inst_mult_0_48  ))
// Xd_0__inst_mult_1_45  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_48 ),
	.sharein(Xd_0__inst_mult_0_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_43_sumout ),
	.cout(Xd_0__inst_mult_1_44 ),
	.shareout(Xd_0__inst_mult_1_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_99 (
// Equation(s):
// Xd_0__inst_mult_7_296  = SUM(( !Xd_0__inst_mult_7_408  $ (!Xd_0__inst_mult_7_412  $ (((din_b[88] & din_a[85])))) ) + ( Xd_0__inst_mult_7_274  ) + ( Xd_0__inst_mult_7_273  ))
// Xd_0__inst_mult_7_297  = CARRY(( !Xd_0__inst_mult_7_408  $ (!Xd_0__inst_mult_7_412  $ (((din_b[88] & din_a[85])))) ) + ( Xd_0__inst_mult_7_274  ) + ( Xd_0__inst_mult_7_273  ))
// Xd_0__inst_mult_7_298  = SHARE((!Xd_0__inst_mult_7_408  & (Xd_0__inst_mult_7_412  & (din_b[88] & din_a[85]))) # (Xd_0__inst_mult_7_408  & (((din_b[88] & din_a[85])) # (Xd_0__inst_mult_7_412 ))))

	.dataa(!Xd_0__inst_mult_7_408 ),
	.datab(!Xd_0__inst_mult_7_412 ),
	.datac(!din_b[88]),
	.datad(!din_a[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_273 ),
	.sharein(Xd_0__inst_mult_7_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_296 ),
	.cout(Xd_0__inst_mult_7_297 ),
	.shareout(Xd_0__inst_mult_7_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_100 (
// Equation(s):
// Xd_0__inst_mult_7_300  = SUM(( (din_a[84] & din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_301  = CARRY(( (din_a[84] & din_b[89]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_302  = SHARE((din_a[84] & din_b[90]))

	.dataa(!din_a[84]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_300 ),
	.cout(Xd_0__inst_mult_7_301 ),
	.shareout(Xd_0__inst_mult_7_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_47 (
// Equation(s):
// Xd_0__inst_mult_2_47_sumout  = SUM(( (din_a[34] & din_b[24]) ) + ( Xd_0__inst_mult_5_49  ) + ( Xd_0__inst_mult_5_48  ))
// Xd_0__inst_mult_2_48  = CARRY(( (din_a[34] & din_b[24]) ) + ( Xd_0__inst_mult_5_49  ) + ( Xd_0__inst_mult_5_48  ))
// Xd_0__inst_mult_2_49  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_48 ),
	.sharein(Xd_0__inst_mult_5_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_47_sumout ),
	.cout(Xd_0__inst_mult_2_48 ),
	.shareout(Xd_0__inst_mult_2_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_99 (
// Equation(s):
// Xd_0__inst_mult_6_296  = SUM(( !Xd_0__inst_mult_6_408  $ (!Xd_0__inst_mult_6_412 ) ) + ( Xd_0__inst_mult_6_290  ) + ( Xd_0__inst_mult_6_289  ))
// Xd_0__inst_mult_6_297  = CARRY(( !Xd_0__inst_mult_6_408  $ (!Xd_0__inst_mult_6_412 ) ) + ( Xd_0__inst_mult_6_290  ) + ( Xd_0__inst_mult_6_289  ))
// Xd_0__inst_mult_6_298  = SHARE((Xd_0__inst_mult_6_408  & Xd_0__inst_mult_6_412 ))

	.dataa(!Xd_0__inst_mult_6_408 ),
	.datab(!Xd_0__inst_mult_6_412 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_289 ),
	.sharein(Xd_0__inst_mult_6_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_296 ),
	.cout(Xd_0__inst_mult_6_297 ),
	.shareout(Xd_0__inst_mult_6_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_100 (
// Equation(s):
// Xd_0__inst_mult_6_300  = SUM(( (din_a[73] & din_b[77]) ) + ( Xd_0__inst_mult_6_294  ) + ( Xd_0__inst_mult_6_293  ))
// Xd_0__inst_mult_6_301  = CARRY(( (din_a[73] & din_b[77]) ) + ( Xd_0__inst_mult_6_294  ) + ( Xd_0__inst_mult_6_293  ))
// Xd_0__inst_mult_6_302  = SHARE((din_a[72] & din_b[79]))

	.dataa(!din_a[73]),
	.datab(!din_b[77]),
	.datac(!din_a[72]),
	.datad(!din_b[79]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_293 ),
	.sharein(Xd_0__inst_mult_6_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_300 ),
	.cout(Xd_0__inst_mult_6_301 ),
	.shareout(Xd_0__inst_mult_6_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_101 (
// Equation(s):
// Xd_0__inst_mult_7_304  = SUM(( !Xd_0__inst_mult_7_416  $ (!Xd_0__inst_mult_7_420 ) ) + ( Xd_0__inst_mult_7_298  ) + ( Xd_0__inst_mult_7_297  ))
// Xd_0__inst_mult_7_305  = CARRY(( !Xd_0__inst_mult_7_416  $ (!Xd_0__inst_mult_7_420 ) ) + ( Xd_0__inst_mult_7_298  ) + ( Xd_0__inst_mult_7_297  ))
// Xd_0__inst_mult_7_306  = SHARE((Xd_0__inst_mult_7_416  & Xd_0__inst_mult_7_420 ))

	.dataa(!Xd_0__inst_mult_7_416 ),
	.datab(!Xd_0__inst_mult_7_420 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_297 ),
	.sharein(Xd_0__inst_mult_7_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_304 ),
	.cout(Xd_0__inst_mult_7_305 ),
	.shareout(Xd_0__inst_mult_7_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_102 (
// Equation(s):
// Xd_0__inst_mult_7_308  = SUM(( (din_a[85] & din_b[89]) ) + ( Xd_0__inst_mult_7_302  ) + ( Xd_0__inst_mult_7_301  ))
// Xd_0__inst_mult_7_309  = CARRY(( (din_a[85] & din_b[89]) ) + ( Xd_0__inst_mult_7_302  ) + ( Xd_0__inst_mult_7_301  ))
// Xd_0__inst_mult_7_310  = SHARE((din_a[84] & din_b[91]))

	.dataa(!din_a[85]),
	.datab(!din_b[89]),
	.datac(!din_a[84]),
	.datad(!din_b[91]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_301 ),
	.sharein(Xd_0__inst_mult_7_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_308 ),
	.cout(Xd_0__inst_mult_7_309 ),
	.shareout(Xd_0__inst_mult_7_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_101 (
// Equation(s):
// Xd_0__inst_mult_6_304  = SUM(( !Xd_0__inst_mult_6_416  $ (!Xd_0__inst_mult_6_420  $ (Xd_0__inst_mult_6_55_sumout )) ) + ( Xd_0__inst_mult_6_298  ) + ( Xd_0__inst_mult_6_297  ))
// Xd_0__inst_mult_6_305  = CARRY(( !Xd_0__inst_mult_6_416  $ (!Xd_0__inst_mult_6_420  $ (Xd_0__inst_mult_6_55_sumout )) ) + ( Xd_0__inst_mult_6_298  ) + ( Xd_0__inst_mult_6_297  ))
// Xd_0__inst_mult_6_306  = SHARE((!Xd_0__inst_mult_6_416  & (Xd_0__inst_mult_6_420  & Xd_0__inst_mult_6_55_sumout )) # (Xd_0__inst_mult_6_416  & ((Xd_0__inst_mult_6_55_sumout ) # (Xd_0__inst_mult_6_420 ))))

	.dataa(!Xd_0__inst_mult_6_416 ),
	.datab(!Xd_0__inst_mult_6_420 ),
	.datac(!Xd_0__inst_mult_6_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_297 ),
	.sharein(Xd_0__inst_mult_6_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_304 ),
	.cout(Xd_0__inst_mult_6_305 ),
	.shareout(Xd_0__inst_mult_6_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_102 (
// Equation(s):
// Xd_0__inst_mult_6_308  = SUM(( (!din_a[73] & (((din_a[74] & din_b[77])))) # (din_a[73] & (!din_b[78] $ (((!din_a[74]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_302  ) + ( Xd_0__inst_mult_6_301  ))
// Xd_0__inst_mult_6_309  = CARRY(( (!din_a[73] & (((din_a[74] & din_b[77])))) # (din_a[73] & (!din_b[78] $ (((!din_a[74]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_302  ) + ( Xd_0__inst_mult_6_301  ))
// Xd_0__inst_mult_6_310  = SHARE((din_a[73] & (din_b[78] & (din_a[74] & din_b[77]))))

	.dataa(!din_a[73]),
	.datab(!din_b[78]),
	.datac(!din_a[74]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_301 ),
	.sharein(Xd_0__inst_mult_6_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_308 ),
	.cout(Xd_0__inst_mult_6_309 ),
	.shareout(Xd_0__inst_mult_6_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_103 (
// Equation(s):
// Xd_0__inst_mult_7_312  = SUM(( !Xd_0__inst_mult_7_424  $ (!Xd_0__inst_mult_7_428  $ (Xd_0__inst_mult_7_55_sumout )) ) + ( Xd_0__inst_mult_7_306  ) + ( Xd_0__inst_mult_7_305  ))
// Xd_0__inst_mult_7_313  = CARRY(( !Xd_0__inst_mult_7_424  $ (!Xd_0__inst_mult_7_428  $ (Xd_0__inst_mult_7_55_sumout )) ) + ( Xd_0__inst_mult_7_306  ) + ( Xd_0__inst_mult_7_305  ))
// Xd_0__inst_mult_7_314  = SHARE((!Xd_0__inst_mult_7_424  & (Xd_0__inst_mult_7_428  & Xd_0__inst_mult_7_55_sumout )) # (Xd_0__inst_mult_7_424  & ((Xd_0__inst_mult_7_55_sumout ) # (Xd_0__inst_mult_7_428 ))))

	.dataa(!Xd_0__inst_mult_7_424 ),
	.datab(!Xd_0__inst_mult_7_428 ),
	.datac(!Xd_0__inst_mult_7_55_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_305 ),
	.sharein(Xd_0__inst_mult_7_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_312 ),
	.cout(Xd_0__inst_mult_7_313 ),
	.shareout(Xd_0__inst_mult_7_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_104 (
// Equation(s):
// Xd_0__inst_mult_7_316  = SUM(( (!din_a[85] & (((din_a[86] & din_b[89])))) # (din_a[85] & (!din_b[90] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_310  ) + ( Xd_0__inst_mult_7_309  ))
// Xd_0__inst_mult_7_317  = CARRY(( (!din_a[85] & (((din_a[86] & din_b[89])))) # (din_a[85] & (!din_b[90] $ (((!din_a[86]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_310  ) + ( Xd_0__inst_mult_7_309  ))
// Xd_0__inst_mult_7_318  = SHARE((din_a[85] & (din_b[90] & (din_a[86] & din_b[89]))))

	.dataa(!din_a[85]),
	.datab(!din_b[90]),
	.datac(!din_a[86]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_309 ),
	.sharein(Xd_0__inst_mult_7_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_316 ),
	.cout(Xd_0__inst_mult_7_317 ),
	.shareout(Xd_0__inst_mult_7_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_103 (
// Equation(s):
// Xd_0__inst_mult_6_312  = SUM(( !Xd_0__inst_mult_6_424  $ (!Xd_0__inst_mult_6_428  $ (Xd_0__inst_mult_6_59_sumout )) ) + ( Xd_0__inst_mult_6_306  ) + ( Xd_0__inst_mult_6_305  ))
// Xd_0__inst_mult_6_313  = CARRY(( !Xd_0__inst_mult_6_424  $ (!Xd_0__inst_mult_6_428  $ (Xd_0__inst_mult_6_59_sumout )) ) + ( Xd_0__inst_mult_6_306  ) + ( Xd_0__inst_mult_6_305  ))
// Xd_0__inst_mult_6_314  = SHARE((!Xd_0__inst_mult_6_424  & (Xd_0__inst_mult_6_428  & Xd_0__inst_mult_6_59_sumout )) # (Xd_0__inst_mult_6_424  & ((Xd_0__inst_mult_6_59_sumout ) # (Xd_0__inst_mult_6_428 ))))

	.dataa(!Xd_0__inst_mult_6_424 ),
	.datab(!Xd_0__inst_mult_6_428 ),
	.datac(!Xd_0__inst_mult_6_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_305 ),
	.sharein(Xd_0__inst_mult_6_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_312 ),
	.cout(Xd_0__inst_mult_6_313 ),
	.shareout(Xd_0__inst_mult_6_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_104 (
// Equation(s):
// Xd_0__inst_mult_6_316  = SUM(( !Xd_0__inst_mult_6_432  $ (((!din_a[73]) # (!din_b[79]))) ) + ( Xd_0__inst_mult_6_438  ) + ( Xd_0__inst_mult_6_437  ))
// Xd_0__inst_mult_6_317  = CARRY(( !Xd_0__inst_mult_6_432  $ (((!din_a[73]) # (!din_b[79]))) ) + ( Xd_0__inst_mult_6_438  ) + ( Xd_0__inst_mult_6_437  ))
// Xd_0__inst_mult_6_318  = SHARE((din_a[73] & (din_b[79] & Xd_0__inst_mult_6_432 )))

	.dataa(!din_a[73]),
	.datab(!din_b[79]),
	.datac(!Xd_0__inst_mult_6_432 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_437 ),
	.sharein(Xd_0__inst_mult_6_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_316 ),
	.cout(Xd_0__inst_mult_6_317 ),
	.shareout(Xd_0__inst_mult_6_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_105 (
// Equation(s):
// Xd_0__inst_mult_7_320  = SUM(( !Xd_0__inst_mult_7_432  $ (!Xd_0__inst_mult_7_436  $ (Xd_0__inst_mult_7_59_sumout )) ) + ( Xd_0__inst_mult_7_314  ) + ( Xd_0__inst_mult_7_313  ))
// Xd_0__inst_mult_7_321  = CARRY(( !Xd_0__inst_mult_7_432  $ (!Xd_0__inst_mult_7_436  $ (Xd_0__inst_mult_7_59_sumout )) ) + ( Xd_0__inst_mult_7_314  ) + ( Xd_0__inst_mult_7_313  ))
// Xd_0__inst_mult_7_322  = SHARE((!Xd_0__inst_mult_7_432  & (Xd_0__inst_mult_7_436  & Xd_0__inst_mult_7_59_sumout )) # (Xd_0__inst_mult_7_432  & ((Xd_0__inst_mult_7_59_sumout ) # (Xd_0__inst_mult_7_436 ))))

	.dataa(!Xd_0__inst_mult_7_432 ),
	.datab(!Xd_0__inst_mult_7_436 ),
	.datac(!Xd_0__inst_mult_7_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_313 ),
	.sharein(Xd_0__inst_mult_7_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_320 ),
	.cout(Xd_0__inst_mult_7_321 ),
	.shareout(Xd_0__inst_mult_7_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_106 (
// Equation(s):
// Xd_0__inst_mult_7_324  = SUM(( !Xd_0__inst_mult_7_440  $ (((!din_a[85]) # (!din_b[91]))) ) + ( Xd_0__inst_mult_7_446  ) + ( Xd_0__inst_mult_7_445  ))
// Xd_0__inst_mult_7_325  = CARRY(( !Xd_0__inst_mult_7_440  $ (((!din_a[85]) # (!din_b[91]))) ) + ( Xd_0__inst_mult_7_446  ) + ( Xd_0__inst_mult_7_445  ))
// Xd_0__inst_mult_7_326  = SHARE((din_a[85] & (din_b[91] & Xd_0__inst_mult_7_440 )))

	.dataa(!din_a[85]),
	.datab(!din_b[91]),
	.datac(!Xd_0__inst_mult_7_440 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_445 ),
	.sharein(Xd_0__inst_mult_7_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_324 ),
	.cout(Xd_0__inst_mult_7_325 ),
	.shareout(Xd_0__inst_mult_7_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_105 (
// Equation(s):
// Xd_0__inst_mult_6_320  = SUM(( !Xd_0__inst_mult_6_440  $ (!Xd_0__inst_mult_6_444  $ (Xd_0__inst_mult_6_63_sumout )) ) + ( Xd_0__inst_mult_6_314  ) + ( Xd_0__inst_mult_6_313  ))
// Xd_0__inst_mult_6_321  = CARRY(( !Xd_0__inst_mult_6_440  $ (!Xd_0__inst_mult_6_444  $ (Xd_0__inst_mult_6_63_sumout )) ) + ( Xd_0__inst_mult_6_314  ) + ( Xd_0__inst_mult_6_313  ))
// Xd_0__inst_mult_6_322  = SHARE((!Xd_0__inst_mult_6_440  & (Xd_0__inst_mult_6_444  & Xd_0__inst_mult_6_63_sumout )) # (Xd_0__inst_mult_6_440  & ((Xd_0__inst_mult_6_63_sumout ) # (Xd_0__inst_mult_6_444 ))))

	.dataa(!Xd_0__inst_mult_6_440 ),
	.datab(!Xd_0__inst_mult_6_444 ),
	.datac(!Xd_0__inst_mult_6_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_313 ),
	.sharein(Xd_0__inst_mult_6_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_320 ),
	.cout(Xd_0__inst_mult_6_321 ),
	.shareout(Xd_0__inst_mult_6_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_106 (
// Equation(s):
// Xd_0__inst_mult_6_324  = SUM(( !Xd_0__inst_mult_6_448  $ (!Xd_0__inst_mult_6_452 ) ) + ( Xd_0__inst_mult_6_318  ) + ( Xd_0__inst_mult_6_317  ))
// Xd_0__inst_mult_6_325  = CARRY(( !Xd_0__inst_mult_6_448  $ (!Xd_0__inst_mult_6_452 ) ) + ( Xd_0__inst_mult_6_318  ) + ( Xd_0__inst_mult_6_317  ))
// Xd_0__inst_mult_6_326  = SHARE((Xd_0__inst_mult_6_448  & Xd_0__inst_mult_6_452 ))

	.dataa(!Xd_0__inst_mult_6_448 ),
	.datab(!Xd_0__inst_mult_6_452 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_317 ),
	.sharein(Xd_0__inst_mult_6_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_324 ),
	.cout(Xd_0__inst_mult_6_325 ),
	.shareout(Xd_0__inst_mult_6_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_107 (
// Equation(s):
// Xd_0__inst_mult_7_328  = SUM(( !Xd_0__inst_mult_7_448  $ (!Xd_0__inst_mult_7_452  $ (Xd_0__inst_mult_7_63_sumout )) ) + ( Xd_0__inst_mult_7_322  ) + ( Xd_0__inst_mult_7_321  ))
// Xd_0__inst_mult_7_329  = CARRY(( !Xd_0__inst_mult_7_448  $ (!Xd_0__inst_mult_7_452  $ (Xd_0__inst_mult_7_63_sumout )) ) + ( Xd_0__inst_mult_7_322  ) + ( Xd_0__inst_mult_7_321  ))
// Xd_0__inst_mult_7_330  = SHARE((!Xd_0__inst_mult_7_448  & (Xd_0__inst_mult_7_452  & Xd_0__inst_mult_7_63_sumout )) # (Xd_0__inst_mult_7_448  & ((Xd_0__inst_mult_7_63_sumout ) # (Xd_0__inst_mult_7_452 ))))

	.dataa(!Xd_0__inst_mult_7_448 ),
	.datab(!Xd_0__inst_mult_7_452 ),
	.datac(!Xd_0__inst_mult_7_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_321 ),
	.sharein(Xd_0__inst_mult_7_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_328 ),
	.cout(Xd_0__inst_mult_7_329 ),
	.shareout(Xd_0__inst_mult_7_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_108 (
// Equation(s):
// Xd_0__inst_mult_7_332  = SUM(( !Xd_0__inst_mult_7_456  $ (!Xd_0__inst_mult_7_460 ) ) + ( Xd_0__inst_mult_7_326  ) + ( Xd_0__inst_mult_7_325  ))
// Xd_0__inst_mult_7_333  = CARRY(( !Xd_0__inst_mult_7_456  $ (!Xd_0__inst_mult_7_460 ) ) + ( Xd_0__inst_mult_7_326  ) + ( Xd_0__inst_mult_7_325  ))
// Xd_0__inst_mult_7_334  = SHARE((Xd_0__inst_mult_7_456  & Xd_0__inst_mult_7_460 ))

	.dataa(!Xd_0__inst_mult_7_456 ),
	.datab(!Xd_0__inst_mult_7_460 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_325 ),
	.sharein(Xd_0__inst_mult_7_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_332 ),
	.cout(Xd_0__inst_mult_7_333 ),
	.shareout(Xd_0__inst_mult_7_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_107 (
// Equation(s):
// Xd_0__inst_mult_6_328  = SUM(( !Xd_0__inst_mult_6_456  $ (!Xd_0__inst_mult_6_460  $ (Xd_0__inst_mult_6_67_sumout )) ) + ( Xd_0__inst_mult_6_322  ) + ( Xd_0__inst_mult_6_321  ))
// Xd_0__inst_mult_6_329  = CARRY(( !Xd_0__inst_mult_6_456  $ (!Xd_0__inst_mult_6_460  $ (Xd_0__inst_mult_6_67_sumout )) ) + ( Xd_0__inst_mult_6_322  ) + ( Xd_0__inst_mult_6_321  ))
// Xd_0__inst_mult_6_330  = SHARE((!Xd_0__inst_mult_6_456  & (Xd_0__inst_mult_6_460  & Xd_0__inst_mult_6_67_sumout )) # (Xd_0__inst_mult_6_456  & ((Xd_0__inst_mult_6_67_sumout ) # (Xd_0__inst_mult_6_460 ))))

	.dataa(!Xd_0__inst_mult_6_456 ),
	.datab(!Xd_0__inst_mult_6_460 ),
	.datac(!Xd_0__inst_mult_6_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_321 ),
	.sharein(Xd_0__inst_mult_6_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_328 ),
	.cout(Xd_0__inst_mult_6_329 ),
	.shareout(Xd_0__inst_mult_6_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_108 (
// Equation(s):
// Xd_0__inst_mult_6_332  = SUM(( !Xd_0__inst_mult_6_464  $ (!Xd_0__inst_mult_6_468  $ (Xd_0__inst_mult_6_472 )) ) + ( Xd_0__inst_mult_6_326  ) + ( Xd_0__inst_mult_6_325  ))
// Xd_0__inst_mult_6_333  = CARRY(( !Xd_0__inst_mult_6_464  $ (!Xd_0__inst_mult_6_468  $ (Xd_0__inst_mult_6_472 )) ) + ( Xd_0__inst_mult_6_326  ) + ( Xd_0__inst_mult_6_325  ))
// Xd_0__inst_mult_6_334  = SHARE((!Xd_0__inst_mult_6_464  & (Xd_0__inst_mult_6_468  & Xd_0__inst_mult_6_472 )) # (Xd_0__inst_mult_6_464  & ((Xd_0__inst_mult_6_472 ) # (Xd_0__inst_mult_6_468 ))))

	.dataa(!Xd_0__inst_mult_6_464 ),
	.datab(!Xd_0__inst_mult_6_468 ),
	.datac(!Xd_0__inst_mult_6_472 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_325 ),
	.sharein(Xd_0__inst_mult_6_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_332 ),
	.cout(Xd_0__inst_mult_6_333 ),
	.shareout(Xd_0__inst_mult_6_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_109 (
// Equation(s):
// Xd_0__inst_mult_7_336  = SUM(( !Xd_0__inst_mult_7_464  $ (!Xd_0__inst_mult_7_468  $ (Xd_0__inst_mult_7_67_sumout )) ) + ( Xd_0__inst_mult_7_330  ) + ( Xd_0__inst_mult_7_329  ))
// Xd_0__inst_mult_7_337  = CARRY(( !Xd_0__inst_mult_7_464  $ (!Xd_0__inst_mult_7_468  $ (Xd_0__inst_mult_7_67_sumout )) ) + ( Xd_0__inst_mult_7_330  ) + ( Xd_0__inst_mult_7_329  ))
// Xd_0__inst_mult_7_338  = SHARE((!Xd_0__inst_mult_7_464  & (Xd_0__inst_mult_7_468  & Xd_0__inst_mult_7_67_sumout )) # (Xd_0__inst_mult_7_464  & ((Xd_0__inst_mult_7_67_sumout ) # (Xd_0__inst_mult_7_468 ))))

	.dataa(!Xd_0__inst_mult_7_464 ),
	.datab(!Xd_0__inst_mult_7_468 ),
	.datac(!Xd_0__inst_mult_7_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_329 ),
	.sharein(Xd_0__inst_mult_7_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_336 ),
	.cout(Xd_0__inst_mult_7_337 ),
	.shareout(Xd_0__inst_mult_7_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_110 (
// Equation(s):
// Xd_0__inst_mult_7_340  = SUM(( !Xd_0__inst_mult_7_472  $ (!Xd_0__inst_mult_7_476  $ (Xd_0__inst_mult_7_480 )) ) + ( Xd_0__inst_mult_7_334  ) + ( Xd_0__inst_mult_7_333  ))
// Xd_0__inst_mult_7_341  = CARRY(( !Xd_0__inst_mult_7_472  $ (!Xd_0__inst_mult_7_476  $ (Xd_0__inst_mult_7_480 )) ) + ( Xd_0__inst_mult_7_334  ) + ( Xd_0__inst_mult_7_333  ))
// Xd_0__inst_mult_7_342  = SHARE((!Xd_0__inst_mult_7_472  & (Xd_0__inst_mult_7_476  & Xd_0__inst_mult_7_480 )) # (Xd_0__inst_mult_7_472  & ((Xd_0__inst_mult_7_480 ) # (Xd_0__inst_mult_7_476 ))))

	.dataa(!Xd_0__inst_mult_7_472 ),
	.datab(!Xd_0__inst_mult_7_476 ),
	.datac(!Xd_0__inst_mult_7_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_333 ),
	.sharein(Xd_0__inst_mult_7_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_340 ),
	.cout(Xd_0__inst_mult_7_341 ),
	.shareout(Xd_0__inst_mult_7_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_109 (
// Equation(s):
// Xd_0__inst_mult_6_336  = SUM(( !Xd_0__inst_mult_6_476  $ (!Xd_0__inst_mult_6_480 ) ) + ( Xd_0__inst_mult_6_330  ) + ( Xd_0__inst_mult_6_329  ))
// Xd_0__inst_mult_6_337  = CARRY(( !Xd_0__inst_mult_6_476  $ (!Xd_0__inst_mult_6_480 ) ) + ( Xd_0__inst_mult_6_330  ) + ( Xd_0__inst_mult_6_329  ))
// Xd_0__inst_mult_6_338  = SHARE((Xd_0__inst_mult_6_476  & Xd_0__inst_mult_6_480 ))

	.dataa(!Xd_0__inst_mult_6_476 ),
	.datab(!Xd_0__inst_mult_6_480 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_329 ),
	.sharein(Xd_0__inst_mult_6_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_336 ),
	.cout(Xd_0__inst_mult_6_337 ),
	.shareout(Xd_0__inst_mult_6_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_110 (
// Equation(s):
// Xd_0__inst_mult_6_340  = SUM(( !Xd_0__inst_mult_6_484  $ (!Xd_0__inst_mult_6_488  $ (Xd_0__inst_mult_6_492 )) ) + ( Xd_0__inst_mult_6_334  ) + ( Xd_0__inst_mult_6_333  ))
// Xd_0__inst_mult_6_341  = CARRY(( !Xd_0__inst_mult_6_484  $ (!Xd_0__inst_mult_6_488  $ (Xd_0__inst_mult_6_492 )) ) + ( Xd_0__inst_mult_6_334  ) + ( Xd_0__inst_mult_6_333  ))
// Xd_0__inst_mult_6_342  = SHARE((!Xd_0__inst_mult_6_484  & (Xd_0__inst_mult_6_488  & Xd_0__inst_mult_6_492 )) # (Xd_0__inst_mult_6_484  & ((Xd_0__inst_mult_6_492 ) # (Xd_0__inst_mult_6_488 ))))

	.dataa(!Xd_0__inst_mult_6_484 ),
	.datab(!Xd_0__inst_mult_6_488 ),
	.datac(!Xd_0__inst_mult_6_492 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_333 ),
	.sharein(Xd_0__inst_mult_6_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_340 ),
	.cout(Xd_0__inst_mult_6_341 ),
	.shareout(Xd_0__inst_mult_6_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_111 (
// Equation(s):
// Xd_0__inst_mult_7_344  = SUM(( !Xd_0__inst_mult_7_484  $ (!Xd_0__inst_mult_7_488 ) ) + ( Xd_0__inst_mult_7_338  ) + ( Xd_0__inst_mult_7_337  ))
// Xd_0__inst_mult_7_345  = CARRY(( !Xd_0__inst_mult_7_484  $ (!Xd_0__inst_mult_7_488 ) ) + ( Xd_0__inst_mult_7_338  ) + ( Xd_0__inst_mult_7_337  ))
// Xd_0__inst_mult_7_346  = SHARE((Xd_0__inst_mult_7_484  & Xd_0__inst_mult_7_488 ))

	.dataa(!Xd_0__inst_mult_7_484 ),
	.datab(!Xd_0__inst_mult_7_488 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_337 ),
	.sharein(Xd_0__inst_mult_7_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_344 ),
	.cout(Xd_0__inst_mult_7_345 ),
	.shareout(Xd_0__inst_mult_7_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_112 (
// Equation(s):
// Xd_0__inst_mult_7_348  = SUM(( !Xd_0__inst_mult_7_492  $ (!Xd_0__inst_mult_7_496  $ (Xd_0__inst_mult_7_500 )) ) + ( Xd_0__inst_mult_7_342  ) + ( Xd_0__inst_mult_7_341  ))
// Xd_0__inst_mult_7_349  = CARRY(( !Xd_0__inst_mult_7_492  $ (!Xd_0__inst_mult_7_496  $ (Xd_0__inst_mult_7_500 )) ) + ( Xd_0__inst_mult_7_342  ) + ( Xd_0__inst_mult_7_341  ))
// Xd_0__inst_mult_7_350  = SHARE((!Xd_0__inst_mult_7_492  & (Xd_0__inst_mult_7_496  & Xd_0__inst_mult_7_500 )) # (Xd_0__inst_mult_7_492  & ((Xd_0__inst_mult_7_500 ) # (Xd_0__inst_mult_7_496 ))))

	.dataa(!Xd_0__inst_mult_7_492 ),
	.datab(!Xd_0__inst_mult_7_496 ),
	.datac(!Xd_0__inst_mult_7_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_341 ),
	.sharein(Xd_0__inst_mult_7_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_348 ),
	.cout(Xd_0__inst_mult_7_349 ),
	.shareout(Xd_0__inst_mult_7_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_111 (
// Equation(s):
// Xd_0__inst_mult_6_344  = SUM(( !Xd_0__inst_mult_6_496  $ (!Xd_0__inst_mult_6_500  $ (((din_b[74] & din_a[82])))) ) + ( Xd_0__inst_mult_6_338  ) + ( Xd_0__inst_mult_6_337  ))
// Xd_0__inst_mult_6_345  = CARRY(( !Xd_0__inst_mult_6_496  $ (!Xd_0__inst_mult_6_500  $ (((din_b[74] & din_a[82])))) ) + ( Xd_0__inst_mult_6_338  ) + ( Xd_0__inst_mult_6_337  ))
// Xd_0__inst_mult_6_346  = SHARE((!Xd_0__inst_mult_6_496  & (Xd_0__inst_mult_6_500  & (din_b[74] & din_a[82]))) # (Xd_0__inst_mult_6_496  & (((din_b[74] & din_a[82])) # (Xd_0__inst_mult_6_500 ))))

	.dataa(!Xd_0__inst_mult_6_496 ),
	.datab(!Xd_0__inst_mult_6_500 ),
	.datac(!din_b[74]),
	.datad(!din_a[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_337 ),
	.sharein(Xd_0__inst_mult_6_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_344 ),
	.cout(Xd_0__inst_mult_6_345 ),
	.shareout(Xd_0__inst_mult_6_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_112 (
// Equation(s):
// Xd_0__inst_mult_6_348  = SUM(( !Xd_0__inst_mult_6_504  $ (!Xd_0__inst_mult_6_508  $ (Xd_0__inst_mult_6_512 )) ) + ( Xd_0__inst_mult_6_342  ) + ( Xd_0__inst_mult_6_341  ))
// Xd_0__inst_mult_6_349  = CARRY(( !Xd_0__inst_mult_6_504  $ (!Xd_0__inst_mult_6_508  $ (Xd_0__inst_mult_6_512 )) ) + ( Xd_0__inst_mult_6_342  ) + ( Xd_0__inst_mult_6_341  ))
// Xd_0__inst_mult_6_350  = SHARE((!Xd_0__inst_mult_6_504  & (Xd_0__inst_mult_6_508  & Xd_0__inst_mult_6_512 )) # (Xd_0__inst_mult_6_504  & ((Xd_0__inst_mult_6_512 ) # (Xd_0__inst_mult_6_508 ))))

	.dataa(!Xd_0__inst_mult_6_504 ),
	.datab(!Xd_0__inst_mult_6_508 ),
	.datac(!Xd_0__inst_mult_6_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_341 ),
	.sharein(Xd_0__inst_mult_6_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_348 ),
	.cout(Xd_0__inst_mult_6_349 ),
	.shareout(Xd_0__inst_mult_6_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_113 (
// Equation(s):
// Xd_0__inst_mult_7_352  = SUM(( !Xd_0__inst_mult_7_504  $ (!Xd_0__inst_mult_7_508  $ (Xd_0__inst_mult_7_512 )) ) + ( Xd_0__inst_mult_7_350  ) + ( Xd_0__inst_mult_7_349  ))
// Xd_0__inst_mult_7_353  = CARRY(( !Xd_0__inst_mult_7_504  $ (!Xd_0__inst_mult_7_508  $ (Xd_0__inst_mult_7_512 )) ) + ( Xd_0__inst_mult_7_350  ) + ( Xd_0__inst_mult_7_349  ))
// Xd_0__inst_mult_7_354  = SHARE((!Xd_0__inst_mult_7_504  & (Xd_0__inst_mult_7_508  & Xd_0__inst_mult_7_512 )) # (Xd_0__inst_mult_7_504  & ((Xd_0__inst_mult_7_512 ) # (Xd_0__inst_mult_7_508 ))))

	.dataa(!Xd_0__inst_mult_7_504 ),
	.datab(!Xd_0__inst_mult_7_508 ),
	.datac(!Xd_0__inst_mult_7_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_349 ),
	.sharein(Xd_0__inst_mult_7_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_352 ),
	.cout(Xd_0__inst_mult_7_353 ),
	.shareout(Xd_0__inst_mult_7_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_113 (
// Equation(s):
// Xd_0__inst_mult_6_352  = SUM(( !Xd_0__inst_mult_6_516  $ (!Xd_0__inst_mult_6_520  $ (Xd_0__inst_mult_6_524 )) ) + ( Xd_0__inst_mult_6_350  ) + ( Xd_0__inst_mult_6_349  ))
// Xd_0__inst_mult_6_353  = CARRY(( !Xd_0__inst_mult_6_516  $ (!Xd_0__inst_mult_6_520  $ (Xd_0__inst_mult_6_524 )) ) + ( Xd_0__inst_mult_6_350  ) + ( Xd_0__inst_mult_6_349  ))
// Xd_0__inst_mult_6_354  = SHARE((!Xd_0__inst_mult_6_516  & (Xd_0__inst_mult_6_520  & Xd_0__inst_mult_6_524 )) # (Xd_0__inst_mult_6_516  & ((Xd_0__inst_mult_6_524 ) # (Xd_0__inst_mult_6_520 ))))

	.dataa(!Xd_0__inst_mult_6_516 ),
	.datab(!Xd_0__inst_mult_6_520 ),
	.datac(!Xd_0__inst_mult_6_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_349 ),
	.sharein(Xd_0__inst_mult_6_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_352 ),
	.cout(Xd_0__inst_mult_6_353 ),
	.shareout(Xd_0__inst_mult_6_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_114 (
// Equation(s):
// Xd_0__inst_mult_7_356  = SUM(( !Xd_0__inst_mult_7_516  $ (!Xd_0__inst_mult_7_520  $ (Xd_0__inst_mult_7_524 )) ) + ( Xd_0__inst_mult_7_354  ) + ( Xd_0__inst_mult_7_353  ))
// Xd_0__inst_mult_7_357  = CARRY(( !Xd_0__inst_mult_7_516  $ (!Xd_0__inst_mult_7_520  $ (Xd_0__inst_mult_7_524 )) ) + ( Xd_0__inst_mult_7_354  ) + ( Xd_0__inst_mult_7_353  ))
// Xd_0__inst_mult_7_358  = SHARE((!Xd_0__inst_mult_7_516  & (Xd_0__inst_mult_7_520  & Xd_0__inst_mult_7_524 )) # (Xd_0__inst_mult_7_516  & ((Xd_0__inst_mult_7_524 ) # (Xd_0__inst_mult_7_520 ))))

	.dataa(!Xd_0__inst_mult_7_516 ),
	.datab(!Xd_0__inst_mult_7_520 ),
	.datac(!Xd_0__inst_mult_7_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_353 ),
	.sharein(Xd_0__inst_mult_7_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_356 ),
	.cout(Xd_0__inst_mult_7_357 ),
	.shareout(Xd_0__inst_mult_7_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_114 (
// Equation(s):
// Xd_0__inst_mult_6_356  = SUM(( !Xd_0__inst_mult_6_528  $ (!Xd_0__inst_mult_6_532  $ (Xd_0__inst_mult_6_536 )) ) + ( Xd_0__inst_mult_6_354  ) + ( Xd_0__inst_mult_6_353  ))
// Xd_0__inst_mult_6_357  = CARRY(( !Xd_0__inst_mult_6_528  $ (!Xd_0__inst_mult_6_532  $ (Xd_0__inst_mult_6_536 )) ) + ( Xd_0__inst_mult_6_354  ) + ( Xd_0__inst_mult_6_353  ))
// Xd_0__inst_mult_6_358  = SHARE((!Xd_0__inst_mult_6_528  & (Xd_0__inst_mult_6_532  & Xd_0__inst_mult_6_536 )) # (Xd_0__inst_mult_6_528  & ((Xd_0__inst_mult_6_536 ) # (Xd_0__inst_mult_6_532 ))))

	.dataa(!Xd_0__inst_mult_6_528 ),
	.datab(!Xd_0__inst_mult_6_532 ),
	.datac(!Xd_0__inst_mult_6_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_353 ),
	.sharein(Xd_0__inst_mult_6_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_356 ),
	.cout(Xd_0__inst_mult_6_357 ),
	.shareout(Xd_0__inst_mult_6_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_115 (
// Equation(s):
// Xd_0__inst_mult_7_360  = SUM(( !Xd_0__inst_mult_7_528  $ (!Xd_0__inst_mult_7_532  $ (Xd_0__inst_mult_7_536 )) ) + ( Xd_0__inst_mult_7_358  ) + ( Xd_0__inst_mult_7_357  ))
// Xd_0__inst_mult_7_361  = CARRY(( !Xd_0__inst_mult_7_528  $ (!Xd_0__inst_mult_7_532  $ (Xd_0__inst_mult_7_536 )) ) + ( Xd_0__inst_mult_7_358  ) + ( Xd_0__inst_mult_7_357  ))
// Xd_0__inst_mult_7_362  = SHARE((!Xd_0__inst_mult_7_528  & (Xd_0__inst_mult_7_532  & Xd_0__inst_mult_7_536 )) # (Xd_0__inst_mult_7_528  & ((Xd_0__inst_mult_7_536 ) # (Xd_0__inst_mult_7_532 ))))

	.dataa(!Xd_0__inst_mult_7_528 ),
	.datab(!Xd_0__inst_mult_7_532 ),
	.datac(!Xd_0__inst_mult_7_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_357 ),
	.sharein(Xd_0__inst_mult_7_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_360 ),
	.cout(Xd_0__inst_mult_7_361 ),
	.shareout(Xd_0__inst_mult_7_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_6_115 (
// Equation(s):
// Xd_0__inst_mult_6_360  = SUM(( !Xd_0__inst_mult_6_540  $ (!Xd_0__inst_mult_6_544  $ (Xd_0__inst_mult_6_548 )) ) + ( Xd_0__inst_mult_6_358  ) + ( Xd_0__inst_mult_6_357  ))
// Xd_0__inst_mult_6_361  = CARRY(( !Xd_0__inst_mult_6_540  $ (!Xd_0__inst_mult_6_544  $ (Xd_0__inst_mult_6_548 )) ) + ( Xd_0__inst_mult_6_358  ) + ( Xd_0__inst_mult_6_357  ))
// Xd_0__inst_mult_6_362  = SHARE((!Xd_0__inst_mult_6_540  & (Xd_0__inst_mult_6_544  & Xd_0__inst_mult_6_548 )) # (Xd_0__inst_mult_6_540  & ((Xd_0__inst_mult_6_548 ) # (Xd_0__inst_mult_6_544 ))))

	.dataa(!Xd_0__inst_mult_6_540 ),
	.datab(!Xd_0__inst_mult_6_544 ),
	.datac(!Xd_0__inst_mult_6_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_357 ),
	.sharein(Xd_0__inst_mult_6_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_360 ),
	.cout(Xd_0__inst_mult_6_361 ),
	.shareout(Xd_0__inst_mult_6_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_7_116 (
// Equation(s):
// Xd_0__inst_mult_7_364  = SUM(( !Xd_0__inst_mult_7_540  $ (!Xd_0__inst_mult_7_544  $ (Xd_0__inst_mult_4_360 )) ) + ( Xd_0__inst_mult_7_362  ) + ( Xd_0__inst_mult_7_361  ))
// Xd_0__inst_mult_7_365  = CARRY(( !Xd_0__inst_mult_7_540  $ (!Xd_0__inst_mult_7_544  $ (Xd_0__inst_mult_4_360 )) ) + ( Xd_0__inst_mult_7_362  ) + ( Xd_0__inst_mult_7_361  ))
// Xd_0__inst_mult_7_366  = SHARE((!Xd_0__inst_mult_7_540  & (Xd_0__inst_mult_7_544  & Xd_0__inst_mult_4_360 )) # (Xd_0__inst_mult_7_540  & ((Xd_0__inst_mult_4_360 ) # (Xd_0__inst_mult_7_544 ))))

	.dataa(!Xd_0__inst_mult_7_540 ),
	.datab(!Xd_0__inst_mult_7_544 ),
	.datac(!Xd_0__inst_mult_4_360 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_361 ),
	.sharein(Xd_0__inst_mult_7_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_364 ),
	.cout(Xd_0__inst_mult_7_365 ),
	.shareout(Xd_0__inst_mult_7_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_6_116 (
// Equation(s):
// Xd_0__inst_mult_6_364  = SUM(( !Xd_0__inst_mult_6_552  $ (!Xd_0__inst_mult_6_556 ) ) + ( Xd_0__inst_mult_6_362  ) + ( Xd_0__inst_mult_6_361  ))
// Xd_0__inst_mult_6_365  = CARRY(( !Xd_0__inst_mult_6_552  $ (!Xd_0__inst_mult_6_556 ) ) + ( Xd_0__inst_mult_6_362  ) + ( Xd_0__inst_mult_6_361  ))
// Xd_0__inst_mult_6_366  = SHARE((Xd_0__inst_mult_6_552  & Xd_0__inst_mult_6_556 ))

	.dataa(!Xd_0__inst_mult_6_552 ),
	.datab(!Xd_0__inst_mult_6_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_361 ),
	.sharein(Xd_0__inst_mult_6_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_364 ),
	.cout(Xd_0__inst_mult_6_365 ),
	.shareout(Xd_0__inst_mult_6_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_35 (
// Equation(s):
// Xd_0__inst_mult_6_35_sumout  = SUM(( (din_a[82] & din_b[78]) ) + ( Xd_0__inst_i29_3  ) + ( Xd_0__inst_i29_2  ))
// Xd_0__inst_mult_6_36  = CARRY(( (din_a[82] & din_b[78]) ) + ( Xd_0__inst_i29_3  ) + ( Xd_0__inst_i29_2  ))
// Xd_0__inst_mult_6_37  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_2 ),
	.sharein(Xd_0__inst_i29_3 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_35_sumout ),
	.cout(Xd_0__inst_mult_6_36 ),
	.shareout(Xd_0__inst_mult_6_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_7_117 (
// Equation(s):
// Xd_0__inst_mult_7_368  = SUM(( !Xd_0__inst_mult_7_548  $ (!Xd_0__inst_mult_7_552 ) ) + ( Xd_0__inst_mult_7_366  ) + ( Xd_0__inst_mult_7_365  ))
// Xd_0__inst_mult_7_369  = CARRY(( !Xd_0__inst_mult_7_548  $ (!Xd_0__inst_mult_7_552 ) ) + ( Xd_0__inst_mult_7_366  ) + ( Xd_0__inst_mult_7_365  ))
// Xd_0__inst_mult_7_370  = SHARE((Xd_0__inst_mult_7_548  & Xd_0__inst_mult_7_552 ))

	.dataa(!Xd_0__inst_mult_7_548 ),
	.datab(!Xd_0__inst_mult_7_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_365 ),
	.sharein(Xd_0__inst_mult_7_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_368 ),
	.cout(Xd_0__inst_mult_7_369 ),
	.shareout(Xd_0__inst_mult_7_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_35 (
// Equation(s):
// Xd_0__inst_mult_7_35_sumout  = SUM(( (din_a[94] & din_b[90]) ) + ( Xd_0__inst_mult_6_57  ) + ( Xd_0__inst_mult_6_56  ))
// Xd_0__inst_mult_7_36  = CARRY(( (din_a[94] & din_b[90]) ) + ( Xd_0__inst_mult_6_57  ) + ( Xd_0__inst_mult_6_56  ))
// Xd_0__inst_mult_7_37  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_56 ),
	.sharein(Xd_0__inst_mult_6_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_35_sumout ),
	.cout(Xd_0__inst_mult_7_36 ),
	.shareout(Xd_0__inst_mult_7_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_6_117 (
// Equation(s):
// Xd_0__inst_mult_6_368  = SUM(( !Xd_0__inst_mult_6_560  $ (!Xd_0__inst_mult_6_564  $ (((din_a[81] & din_b[80])))) ) + ( Xd_0__inst_mult_6_366  ) + ( Xd_0__inst_mult_6_365  ))
// Xd_0__inst_mult_6_369  = CARRY(( !Xd_0__inst_mult_6_560  $ (!Xd_0__inst_mult_6_564  $ (((din_a[81] & din_b[80])))) ) + ( Xd_0__inst_mult_6_366  ) + ( Xd_0__inst_mult_6_365  ))
// Xd_0__inst_mult_6_370  = SHARE((!Xd_0__inst_mult_6_560  & (Xd_0__inst_mult_6_564  & (din_a[81] & din_b[80]))) # (Xd_0__inst_mult_6_560  & (((din_a[81] & din_b[80])) # (Xd_0__inst_mult_6_564 ))))

	.dataa(!Xd_0__inst_mult_6_560 ),
	.datab(!Xd_0__inst_mult_6_564 ),
	.datac(!din_a[81]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_365 ),
	.sharein(Xd_0__inst_mult_6_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_368 ),
	.cout(Xd_0__inst_mult_6_369 ),
	.shareout(Xd_0__inst_mult_6_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_39 (
// Equation(s):
// Xd_0__inst_mult_6_39_sumout  = SUM(( (din_a[82] & din_b[79]) ) + ( Xd_0__inst_mult_7_57  ) + ( Xd_0__inst_mult_7_56  ))
// Xd_0__inst_mult_6_40  = CARRY(( (din_a[82] & din_b[79]) ) + ( Xd_0__inst_mult_7_57  ) + ( Xd_0__inst_mult_7_56  ))
// Xd_0__inst_mult_6_41  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_56 ),
	.sharein(Xd_0__inst_mult_7_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_39_sumout ),
	.cout(Xd_0__inst_mult_6_40 ),
	.shareout(Xd_0__inst_mult_6_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_7_118 (
// Equation(s):
// Xd_0__inst_mult_7_372  = SUM(( !Xd_0__inst_mult_7_556  $ (!Xd_0__inst_mult_7_560  $ (((din_a[93] & din_b[92])))) ) + ( Xd_0__inst_mult_7_370  ) + ( Xd_0__inst_mult_7_369  ))
// Xd_0__inst_mult_7_373  = CARRY(( !Xd_0__inst_mult_7_556  $ (!Xd_0__inst_mult_7_560  $ (((din_a[93] & din_b[92])))) ) + ( Xd_0__inst_mult_7_370  ) + ( Xd_0__inst_mult_7_369  ))
// Xd_0__inst_mult_7_374  = SHARE((!Xd_0__inst_mult_7_556  & (Xd_0__inst_mult_7_560  & (din_a[93] & din_b[92]))) # (Xd_0__inst_mult_7_556  & (((din_a[93] & din_b[92])) # (Xd_0__inst_mult_7_560 ))))

	.dataa(!Xd_0__inst_mult_7_556 ),
	.datab(!Xd_0__inst_mult_7_560 ),
	.datac(!din_a[93]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_369 ),
	.sharein(Xd_0__inst_mult_7_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_372 ),
	.cout(Xd_0__inst_mult_7_373 ),
	.shareout(Xd_0__inst_mult_7_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_39 (
// Equation(s):
// Xd_0__inst_mult_7_39_sumout  = SUM(( (din_a[94] & din_b[91]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_40  = CARRY(( (din_a[94] & din_b[91]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_41  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_39_sumout ),
	.cout(Xd_0__inst_mult_7_40 ),
	.shareout(Xd_0__inst_mult_7_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_118 (
// Equation(s):
// Xd_0__inst_mult_6_372  = SUM(( !Xd_0__inst_mult_6_568  $ (((!din_a[81]) # (!din_b[81]))) ) + ( Xd_0__inst_mult_6_370  ) + ( Xd_0__inst_mult_6_369  ))
// Xd_0__inst_mult_6_373  = CARRY(( !Xd_0__inst_mult_6_568  $ (((!din_a[81]) # (!din_b[81]))) ) + ( Xd_0__inst_mult_6_370  ) + ( Xd_0__inst_mult_6_369  ))
// Xd_0__inst_mult_6_374  = SHARE((din_a[81] & (din_b[81] & Xd_0__inst_mult_6_568 )))

	.dataa(!din_a[81]),
	.datab(!din_b[81]),
	.datac(!Xd_0__inst_mult_6_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_369 ),
	.sharein(Xd_0__inst_mult_6_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_372 ),
	.cout(Xd_0__inst_mult_6_373 ),
	.shareout(Xd_0__inst_mult_6_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_43 (
// Equation(s):
// Xd_0__inst_mult_6_43_sumout  = SUM(( (din_a[82] & din_b[80]) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_6_44  = CARRY(( (din_a[82] & din_b[80]) ) + ( Xd_0__inst_mult_7_41  ) + ( Xd_0__inst_mult_7_40  ))
// Xd_0__inst_mult_6_45  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_40 ),
	.sharein(Xd_0__inst_mult_7_41 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_43_sumout ),
	.cout(Xd_0__inst_mult_6_44 ),
	.shareout(Xd_0__inst_mult_6_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_119 (
// Equation(s):
// Xd_0__inst_mult_7_376  = SUM(( !Xd_0__inst_mult_7_564  $ (((!din_a[93]) # (!din_b[93]))) ) + ( Xd_0__inst_mult_7_374  ) + ( Xd_0__inst_mult_7_373  ))
// Xd_0__inst_mult_7_377  = CARRY(( !Xd_0__inst_mult_7_564  $ (((!din_a[93]) # (!din_b[93]))) ) + ( Xd_0__inst_mult_7_374  ) + ( Xd_0__inst_mult_7_373  ))
// Xd_0__inst_mult_7_378  = SHARE((din_a[93] & (din_b[93] & Xd_0__inst_mult_7_564 )))

	.dataa(!din_a[93]),
	.datab(!din_b[93]),
	.datac(!Xd_0__inst_mult_7_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_373 ),
	.sharein(Xd_0__inst_mult_7_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_376 ),
	.cout(Xd_0__inst_mult_7_377 ),
	.shareout(Xd_0__inst_mult_7_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_43 (
// Equation(s):
// Xd_0__inst_mult_7_43_sumout  = SUM(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_6_45  ) + ( Xd_0__inst_mult_6_44  ))
// Xd_0__inst_mult_7_44  = CARRY(( (din_a[94] & din_b[92]) ) + ( Xd_0__inst_mult_6_45  ) + ( Xd_0__inst_mult_6_44  ))
// Xd_0__inst_mult_7_45  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_44 ),
	.sharein(Xd_0__inst_mult_6_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_43_sumout ),
	.cout(Xd_0__inst_mult_7_44 ),
	.shareout(Xd_0__inst_mult_7_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_6_119 (
// Equation(s):
// Xd_0__inst_mult_6_376  = SUM(( !Xd_0__inst_mult_6_572  $ (((!din_a[81]) # (!din_b[82]))) ) + ( Xd_0__inst_mult_6_374  ) + ( Xd_0__inst_mult_6_373  ))
// Xd_0__inst_mult_6_377  = CARRY(( !Xd_0__inst_mult_6_572  $ (((!din_a[81]) # (!din_b[82]))) ) + ( Xd_0__inst_mult_6_374  ) + ( Xd_0__inst_mult_6_373  ))
// Xd_0__inst_mult_6_378  = SHARE((din_a[81] & (din_b[82] & Xd_0__inst_mult_6_572 )))

	.dataa(!din_a[81]),
	.datab(!din_b[82]),
	.datac(!Xd_0__inst_mult_6_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_373 ),
	.sharein(Xd_0__inst_mult_6_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_376 ),
	.cout(Xd_0__inst_mult_6_377 ),
	.shareout(Xd_0__inst_mult_6_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_47 (
// Equation(s):
// Xd_0__inst_mult_6_47_sumout  = SUM(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_7_45  ) + ( Xd_0__inst_mult_7_44  ))
// Xd_0__inst_mult_6_48  = CARRY(( (din_a[82] & din_b[81]) ) + ( Xd_0__inst_mult_7_45  ) + ( Xd_0__inst_mult_7_44  ))
// Xd_0__inst_mult_6_49  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[81]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_44 ),
	.sharein(Xd_0__inst_mult_7_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_47_sumout ),
	.cout(Xd_0__inst_mult_6_48 ),
	.shareout(Xd_0__inst_mult_6_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_7_120 (
// Equation(s):
// Xd_0__inst_mult_7_380  = SUM(( !Xd_0__inst_mult_7_568  $ (((!din_a[93]) # (!din_b[94]))) ) + ( Xd_0__inst_mult_7_378  ) + ( Xd_0__inst_mult_7_377  ))
// Xd_0__inst_mult_7_381  = CARRY(( !Xd_0__inst_mult_7_568  $ (((!din_a[93]) # (!din_b[94]))) ) + ( Xd_0__inst_mult_7_378  ) + ( Xd_0__inst_mult_7_377  ))
// Xd_0__inst_mult_7_382  = SHARE((din_a[93] & (din_b[94] & Xd_0__inst_mult_7_568 )))

	.dataa(!din_a[93]),
	.datab(!din_b[94]),
	.datac(!Xd_0__inst_mult_7_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_377 ),
	.sharein(Xd_0__inst_mult_7_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_380 ),
	.cout(Xd_0__inst_mult_7_381 ),
	.shareout(Xd_0__inst_mult_7_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_47 (
// Equation(s):
// Xd_0__inst_mult_7_47_sumout  = SUM(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_6_49  ) + ( Xd_0__inst_mult_6_48  ))
// Xd_0__inst_mult_7_48  = CARRY(( (din_a[94] & din_b[93]) ) + ( Xd_0__inst_mult_6_49  ) + ( Xd_0__inst_mult_6_48  ))
// Xd_0__inst_mult_7_49  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[93]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_48 ),
	.sharein(Xd_0__inst_mult_6_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_47_sumout ),
	.cout(Xd_0__inst_mult_7_48 ),
	.shareout(Xd_0__inst_mult_7_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_120 (
// Equation(s):
// Xd_0__inst_mult_6_380  = SUM(( GND ) + ( Xd_0__inst_mult_6_378  ) + ( Xd_0__inst_mult_6_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_377 ),
	.sharein(Xd_0__inst_mult_6_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_51 (
// Equation(s):
// Xd_0__inst_mult_6_51_sumout  = SUM(( (din_a[82] & din_b[82]) ) + ( Xd_0__inst_mult_7_49  ) + ( Xd_0__inst_mult_7_48  ))
// Xd_0__inst_mult_6_52  = CARRY(( (din_a[82] & din_b[82]) ) + ( Xd_0__inst_mult_7_49  ) + ( Xd_0__inst_mult_7_48  ))
// Xd_0__inst_mult_6_53  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_48 ),
	.sharein(Xd_0__inst_mult_7_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_51_sumout ),
	.cout(Xd_0__inst_mult_6_52 ),
	.shareout(Xd_0__inst_mult_6_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_121 (
// Equation(s):
// Xd_0__inst_mult_7_384  = SUM(( GND ) + ( Xd_0__inst_mult_7_382  ) + ( Xd_0__inst_mult_7_381  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_381 ),
	.sharein(Xd_0__inst_mult_7_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_384 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_51 (
// Equation(s):
// Xd_0__inst_mult_7_51_sumout  = SUM(( (din_a[94] & din_b[94]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_52  = CARRY(( (din_a[94] & din_b[94]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_53  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_51_sumout ),
	.cout(Xd_0__inst_mult_7_52 ),
	.shareout(Xd_0__inst_mult_7_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_95 (
// Equation(s):
// Xd_0__inst_mult_3_292  = SUM(( (din_a[45] & din_b[40]) ) + ( Xd_0__inst_mult_3_410  ) + ( Xd_0__inst_mult_3_409  ))
// Xd_0__inst_mult_3_293  = CARRY(( (din_a[45] & din_b[40]) ) + ( Xd_0__inst_mult_3_410  ) + ( Xd_0__inst_mult_3_409  ))
// Xd_0__inst_mult_3_294  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[40]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_409 ),
	.sharein(Xd_0__inst_mult_3_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_292 ),
	.cout(Xd_0__inst_mult_3_293 ),
	.shareout(Xd_0__inst_mult_3_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_96 (
// Equation(s):
// Xd_0__inst_mult_3_296  = SUM(( !Xd_0__inst_mult_3_412  $ (!Xd_0__inst_mult_3_408  $ (((din_b[38] & din_a[46])))) ) + ( Xd_0__inst_mult_3_366  ) + ( Xd_0__inst_mult_3_365  ))
// Xd_0__inst_mult_3_297  = CARRY(( !Xd_0__inst_mult_3_412  $ (!Xd_0__inst_mult_3_408  $ (((din_b[38] & din_a[46])))) ) + ( Xd_0__inst_mult_3_366  ) + ( Xd_0__inst_mult_3_365  ))
// Xd_0__inst_mult_3_298  = SHARE((!Xd_0__inst_mult_3_412  & (Xd_0__inst_mult_3_408  & (din_b[38] & din_a[46]))) # (Xd_0__inst_mult_3_412  & (((din_b[38] & din_a[46])) # (Xd_0__inst_mult_3_408 ))))

	.dataa(!Xd_0__inst_mult_3_412 ),
	.datab(!Xd_0__inst_mult_3_408 ),
	.datac(!din_b[38]),
	.datad(!din_a[46]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_365 ),
	.sharein(Xd_0__inst_mult_3_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_296 ),
	.cout(Xd_0__inst_mult_3_297 ),
	.shareout(Xd_0__inst_mult_3_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_121 (
// Equation(s):
// Xd_0__inst_mult_6_384  = SUM(( (din_a[81] & din_b[76]) ) + ( Xd_0__inst_mult_6_502  ) + ( Xd_0__inst_mult_6_501  ))
// Xd_0__inst_mult_6_385  = CARRY(( (din_a[81] & din_b[76]) ) + ( Xd_0__inst_mult_6_502  ) + ( Xd_0__inst_mult_6_501  ))
// Xd_0__inst_mult_6_386  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[76]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_501 ),
	.sharein(Xd_0__inst_mult_6_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_384 ),
	.cout(Xd_0__inst_mult_6_385 ),
	.shareout(Xd_0__inst_mult_6_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_39 (
// Equation(s):
// Xd_0__inst_mult_3_39_sumout  = SUM(( (din_a[46] & din_b[42]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_40  = CARRY(( (din_a[46] & din_b[42]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_41  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_39_sumout ),
	.cout(Xd_0__inst_mult_3_40 ),
	.shareout(Xd_0__inst_mult_3_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_90 (
// Equation(s):
// Xd_0__inst_mult_0_272  = SUM(( (din_a[9] & din_b[4]) ) + ( Xd_0__inst_mult_0_386  ) + ( Xd_0__inst_mult_0_385  ))
// Xd_0__inst_mult_0_273  = CARRY(( (din_a[9] & din_b[4]) ) + ( Xd_0__inst_mult_0_386  ) + ( Xd_0__inst_mult_0_385  ))
// Xd_0__inst_mult_0_274  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[4]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_385 ),
	.sharein(Xd_0__inst_mult_0_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_272 ),
	.cout(Xd_0__inst_mult_0_273 ),
	.shareout(Xd_0__inst_mult_0_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_91 (
// Equation(s):
// Xd_0__inst_mult_0_276  = SUM(( !Xd_0__inst_mult_0_388  $ (!Xd_0__inst_mult_0_384  $ (((din_b[2] & din_a[10])))) ) + ( Xd_0__inst_mult_0_342  ) + ( Xd_0__inst_mult_0_341  ))
// Xd_0__inst_mult_0_277  = CARRY(( !Xd_0__inst_mult_0_388  $ (!Xd_0__inst_mult_0_384  $ (((din_b[2] & din_a[10])))) ) + ( Xd_0__inst_mult_0_342  ) + ( Xd_0__inst_mult_0_341  ))
// Xd_0__inst_mult_0_278  = SHARE((!Xd_0__inst_mult_0_388  & (Xd_0__inst_mult_0_384  & (din_b[2] & din_a[10]))) # (Xd_0__inst_mult_0_388  & (((din_b[2] & din_a[10])) # (Xd_0__inst_mult_0_384 ))))

	.dataa(!Xd_0__inst_mult_0_388 ),
	.datab(!Xd_0__inst_mult_0_384 ),
	.datac(!din_b[2]),
	.datad(!din_a[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_341 ),
	.sharein(Xd_0__inst_mult_0_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_276 ),
	.cout(Xd_0__inst_mult_0_277 ),
	.shareout(Xd_0__inst_mult_0_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_97 (
// Equation(s):
// Xd_0__inst_mult_3_300  = SUM(( (din_a[41] & din_b[45]) ) + ( Xd_0__inst_mult_3_418  ) + ( Xd_0__inst_mult_3_417  ))
// Xd_0__inst_mult_3_301  = CARRY(( (din_a[41] & din_b[45]) ) + ( Xd_0__inst_mult_3_418  ) + ( Xd_0__inst_mult_3_417  ))
// Xd_0__inst_mult_3_302  = SHARE((din_a[41] & din_b[46]))

	.dataa(!din_a[41]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_417 ),
	.sharein(Xd_0__inst_mult_3_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_300 ),
	.cout(Xd_0__inst_mult_3_301 ),
	.shareout(Xd_0__inst_mult_3_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_122 (
// Equation(s):
// Xd_0__inst_mult_7_388  = SUM(( (!din_a[93] & (((din_a[92] & din_b[88])))) # (din_a[93] & (!din_b[87] $ (((!din_a[92]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_490  ) + ( Xd_0__inst_mult_7_489  ))
// Xd_0__inst_mult_7_389  = CARRY(( (!din_a[93] & (((din_a[92] & din_b[88])))) # (din_a[93] & (!din_b[87] $ (((!din_a[92]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_490  ) + ( Xd_0__inst_mult_7_489  ))
// Xd_0__inst_mult_7_390  = SHARE((din_a[93] & (din_b[87] & (din_a[92] & din_b[88]))))

	.dataa(!din_a[93]),
	.datab(!din_b[87]),
	.datac(!din_a[92]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_489 ),
	.sharein(Xd_0__inst_mult_7_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_388 ),
	.cout(Xd_0__inst_mult_7_389 ),
	.shareout(Xd_0__inst_mult_7_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_123 (
// Equation(s):
// Xd_0__inst_mult_7_392  = SUM(( GND ) + ( Xd_0__inst_mult_7_486  ) + ( Xd_0__inst_mult_7_485  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_485 ),
	.sharein(Xd_0__inst_mult_7_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_392 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_4_90 (
// Equation(s):
// Xd_0__inst_mult_4_261  = CARRY(( Xd_0__inst_mult_4_384  ) + ( Xd_0__inst_mult_4_390  ) + ( Xd_0__inst_mult_4_389  ))
// Xd_0__inst_mult_4_262  = SHARE((din_a[49] & din_b[50]))

	.dataa(!Xd_0__inst_mult_4_384 ),
	.datab(!din_a[49]),
	.datac(!din_b[50]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_389 ),
	.sharein(Xd_0__inst_mult_4_390 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_261 ),
	.shareout(Xd_0__inst_mult_4_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_5_90 (
// Equation(s):
// Xd_0__inst_mult_5_261  = CARRY(( Xd_0__inst_mult_5_380  ) + ( Xd_0__inst_mult_5_386  ) + ( Xd_0__inst_mult_5_385  ))
// Xd_0__inst_mult_5_262  = SHARE((din_a[61] & din_b[62]))

	.dataa(!Xd_0__inst_mult_5_380 ),
	.datab(!din_a[61]),
	.datac(!din_b[62]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_385 ),
	.sharein(Xd_0__inst_mult_5_386 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_261 ),
	.shareout(Xd_0__inst_mult_5_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_2_90 (
// Equation(s):
// Xd_0__inst_mult_2_261  = CARRY(( Xd_0__inst_mult_2_380  ) + ( Xd_0__inst_mult_2_386  ) + ( Xd_0__inst_mult_2_385  ))
// Xd_0__inst_mult_2_262  = SHARE((din_a[25] & din_b[26]))

	.dataa(!Xd_0__inst_mult_2_380 ),
	.datab(!din_a[25]),
	.datac(!din_b[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_385 ),
	.sharein(Xd_0__inst_mult_2_386 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_261 ),
	.shareout(Xd_0__inst_mult_2_262 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_3_98 (
// Equation(s):
// Xd_0__inst_mult_3_305  = CARRY(( Xd_0__inst_mult_3_420  ) + ( Xd_0__inst_mult_3_426  ) + ( Xd_0__inst_mult_3_425  ))
// Xd_0__inst_mult_3_306  = SHARE((din_a[37] & din_b[38]))

	.dataa(!Xd_0__inst_mult_3_420 ),
	.datab(!din_a[37]),
	.datac(!din_b[38]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_425 ),
	.sharein(Xd_0__inst_mult_3_426 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_305 ),
	.shareout(Xd_0__inst_mult_3_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_0_92 (
// Equation(s):
// Xd_0__inst_mult_0_281  = CARRY(( Xd_0__inst_mult_0_392  ) + ( Xd_0__inst_mult_0_398  ) + ( Xd_0__inst_mult_0_397  ))
// Xd_0__inst_mult_0_282  = SHARE((din_a[1] & din_b[2]))

	.dataa(!Xd_0__inst_mult_0_392 ),
	.datab(!din_a[1]),
	.datac(!din_b[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_397 ),
	.sharein(Xd_0__inst_mult_0_398 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_281 ),
	.shareout(Xd_0__inst_mult_0_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300005555),
	.shared_arith("on")
) Xd_0__inst_mult_1_88 (
// Equation(s):
// Xd_0__inst_mult_1_265  = CARRY(( Xd_0__inst_mult_1_173  ) + ( Xd_0__inst_mult_1_171  ) + ( Xd_0__inst_mult_1_170  ))
// Xd_0__inst_mult_1_266  = SHARE((din_a[13] & din_b[14]))

	.dataa(!Xd_0__inst_mult_1_173 ),
	.datab(!din_a[13]),
	.datac(!din_b[14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_170 ),
	.sharein(Xd_0__inst_mult_1_171 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_265 ),
	.shareout(Xd_0__inst_mult_1_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_122 (
// Equation(s):
// Xd_0__inst_mult_6_388  = SUM(( (!din_a[74] & (((din_a[75] & din_b[72])))) # (din_a[74] & (!din_b[73] $ (((!din_a[75]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_258  ) + ( Xd_0__inst_mult_6_257  ))
// Xd_0__inst_mult_6_389  = CARRY(( (!din_a[74] & (((din_a[75] & din_b[72])))) # (din_a[74] & (!din_b[73] $ (((!din_a[75]) # (!din_b[72]))))) ) + ( Xd_0__inst_mult_6_258  ) + ( Xd_0__inst_mult_6_257  ))
// Xd_0__inst_mult_6_390  = SHARE((din_a[74] & (din_b[73] & (din_a[75] & din_b[72]))))

	.dataa(!din_a[74]),
	.datab(!din_b[73]),
	.datac(!din_a[75]),
	.datad(!din_b[72]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_257 ),
	.sharein(Xd_0__inst_mult_6_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_388 ),
	.cout(Xd_0__inst_mult_6_389 ),
	.shareout(Xd_0__inst_mult_6_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_123 (
// Equation(s):
// Xd_0__inst_mult_6_393  = CARRY(( GND ) + ( Xd_0__inst_mult_5_65  ) + ( Xd_0__inst_mult_5_64  ))
// Xd_0__inst_mult_6_394  = SHARE(Xd_0__inst_mult_6_388 )

	.dataa(!Xd_0__inst_mult_6_388 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_64 ),
	.sharein(Xd_0__inst_mult_5_65 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_393 ),
	.shareout(Xd_0__inst_mult_6_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_124 (
// Equation(s):
// Xd_0__inst_mult_7_396  = SUM(( (!din_a[86] & (((din_a[87] & din_b[84])))) # (din_a[86] & (!din_b[85] $ (((!din_a[87]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_266  ) + ( Xd_0__inst_mult_7_265  ))
// Xd_0__inst_mult_7_397  = CARRY(( (!din_a[86] & (((din_a[87] & din_b[84])))) # (din_a[86] & (!din_b[85] $ (((!din_a[87]) # (!din_b[84]))))) ) + ( Xd_0__inst_mult_7_266  ) + ( Xd_0__inst_mult_7_265  ))
// Xd_0__inst_mult_7_398  = SHARE((din_a[86] & (din_b[85] & (din_a[87] & din_b[84]))))

	.dataa(!din_a[86]),
	.datab(!din_b[85]),
	.datac(!din_a[87]),
	.datad(!din_b[84]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_265 ),
	.sharein(Xd_0__inst_mult_7_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_396 ),
	.cout(Xd_0__inst_mult_7_397 ),
	.shareout(Xd_0__inst_mult_7_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_125 (
// Equation(s):
// Xd_0__inst_mult_7_401  = CARRY(( GND ) + ( Xd_0__inst_mult_3_53  ) + ( Xd_0__inst_mult_3_52  ))
// Xd_0__inst_mult_7_402  = SHARE(Xd_0__inst_mult_7_396 )

	.dataa(!Xd_0__inst_mult_7_396 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_52 ),
	.sharein(Xd_0__inst_mult_3_53 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_401 ),
	.shareout(Xd_0__inst_mult_7_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_91 (
// Equation(s):
// Xd_0__inst_mult_4_264  = SUM(( (din_a[52] & din_b[48]) ) + ( Xd_0__inst_mult_4_386  ) + ( Xd_0__inst_mult_4_385  ))
// Xd_0__inst_mult_4_265  = CARRY(( (din_a[52] & din_b[48]) ) + ( Xd_0__inst_mult_4_386  ) + ( Xd_0__inst_mult_4_385  ))
// Xd_0__inst_mult_4_266  = SHARE((din_a[52] & din_b[49]))

	.dataa(!din_a[52]),
	.datab(!din_b[48]),
	.datac(!din_b[49]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_385 ),
	.sharein(Xd_0__inst_mult_4_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_264 ),
	.cout(Xd_0__inst_mult_4_265 ),
	.shareout(Xd_0__inst_mult_4_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_92 (
// Equation(s):
// Xd_0__inst_mult_4_268  = SUM(( (din_a[49] & din_b[51]) ) + ( Xd_0__inst_mult_4_394  ) + ( Xd_0__inst_mult_4_393  ))
// Xd_0__inst_mult_4_269  = CARRY(( (din_a[49] & din_b[51]) ) + ( Xd_0__inst_mult_4_394  ) + ( Xd_0__inst_mult_4_393  ))
// Xd_0__inst_mult_4_270  = SHARE((din_b[51] & din_a[50]))

	.dataa(!din_a[49]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_393 ),
	.sharein(Xd_0__inst_mult_4_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_268 ),
	.cout(Xd_0__inst_mult_4_269 ),
	.shareout(Xd_0__inst_mult_4_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_91 (
// Equation(s):
// Xd_0__inst_mult_5_264  = SUM(( (din_a[64] & din_b[60]) ) + ( Xd_0__inst_mult_5_382  ) + ( Xd_0__inst_mult_5_381  ))
// Xd_0__inst_mult_5_265  = CARRY(( (din_a[64] & din_b[60]) ) + ( Xd_0__inst_mult_5_382  ) + ( Xd_0__inst_mult_5_381  ))
// Xd_0__inst_mult_5_266  = SHARE((din_a[64] & din_b[61]))

	.dataa(!din_a[64]),
	.datab(!din_b[60]),
	.datac(!din_b[61]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_381 ),
	.sharein(Xd_0__inst_mult_5_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_264 ),
	.cout(Xd_0__inst_mult_5_265 ),
	.shareout(Xd_0__inst_mult_5_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_92 (
// Equation(s):
// Xd_0__inst_mult_5_268  = SUM(( (din_a[61] & din_b[63]) ) + ( Xd_0__inst_mult_5_390  ) + ( Xd_0__inst_mult_5_389  ))
// Xd_0__inst_mult_5_269  = CARRY(( (din_a[61] & din_b[63]) ) + ( Xd_0__inst_mult_5_390  ) + ( Xd_0__inst_mult_5_389  ))
// Xd_0__inst_mult_5_270  = SHARE((din_b[63] & din_a[62]))

	.dataa(!din_a[61]),
	.datab(!din_b[63]),
	.datac(!din_a[62]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_389 ),
	.sharein(Xd_0__inst_mult_5_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_268 ),
	.cout(Xd_0__inst_mult_5_269 ),
	.shareout(Xd_0__inst_mult_5_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_91 (
// Equation(s):
// Xd_0__inst_mult_2_264  = SUM(( (din_a[28] & din_b[24]) ) + ( Xd_0__inst_mult_2_382  ) + ( Xd_0__inst_mult_2_381  ))
// Xd_0__inst_mult_2_265  = CARRY(( (din_a[28] & din_b[24]) ) + ( Xd_0__inst_mult_2_382  ) + ( Xd_0__inst_mult_2_381  ))
// Xd_0__inst_mult_2_266  = SHARE((din_a[28] & din_b[25]))

	.dataa(!din_a[28]),
	.datab(!din_b[24]),
	.datac(!din_b[25]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_381 ),
	.sharein(Xd_0__inst_mult_2_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_264 ),
	.cout(Xd_0__inst_mult_2_265 ),
	.shareout(Xd_0__inst_mult_2_266 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_92 (
// Equation(s):
// Xd_0__inst_mult_2_268  = SUM(( (din_a[25] & din_b[27]) ) + ( Xd_0__inst_mult_2_390  ) + ( Xd_0__inst_mult_2_389  ))
// Xd_0__inst_mult_2_269  = CARRY(( (din_a[25] & din_b[27]) ) + ( Xd_0__inst_mult_2_390  ) + ( Xd_0__inst_mult_2_389  ))
// Xd_0__inst_mult_2_270  = SHARE((din_b[27] & din_a[26]))

	.dataa(!din_a[25]),
	.datab(!din_b[27]),
	.datac(!din_a[26]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_389 ),
	.sharein(Xd_0__inst_mult_2_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_268 ),
	.cout(Xd_0__inst_mult_2_269 ),
	.shareout(Xd_0__inst_mult_2_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_99 (
// Equation(s):
// Xd_0__inst_mult_3_308  = SUM(( (din_a[40] & din_b[36]) ) + ( Xd_0__inst_mult_3_422  ) + ( Xd_0__inst_mult_3_421  ))
// Xd_0__inst_mult_3_309  = CARRY(( (din_a[40] & din_b[36]) ) + ( Xd_0__inst_mult_3_422  ) + ( Xd_0__inst_mult_3_421  ))
// Xd_0__inst_mult_3_310  = SHARE((din_a[40] & din_b[37]))

	.dataa(!din_a[40]),
	.datab(!din_b[36]),
	.datac(!din_b[37]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_421 ),
	.sharein(Xd_0__inst_mult_3_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_308 ),
	.cout(Xd_0__inst_mult_3_309 ),
	.shareout(Xd_0__inst_mult_3_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_100 (
// Equation(s):
// Xd_0__inst_mult_3_312  = SUM(( (din_a[37] & din_b[39]) ) + ( Xd_0__inst_mult_3_430  ) + ( Xd_0__inst_mult_3_429  ))
// Xd_0__inst_mult_3_313  = CARRY(( (din_a[37] & din_b[39]) ) + ( Xd_0__inst_mult_3_430  ) + ( Xd_0__inst_mult_3_429  ))
// Xd_0__inst_mult_3_314  = SHARE((din_b[39] & din_a[38]))

	.dataa(!din_a[37]),
	.datab(!din_b[39]),
	.datac(!din_a[38]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_429 ),
	.sharein(Xd_0__inst_mult_3_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_312 ),
	.cout(Xd_0__inst_mult_3_313 ),
	.shareout(Xd_0__inst_mult_3_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_93 (
// Equation(s):
// Xd_0__inst_mult_0_284  = SUM(( (din_a[4] & din_b[0]) ) + ( Xd_0__inst_mult_0_394  ) + ( Xd_0__inst_mult_0_393  ))
// Xd_0__inst_mult_0_285  = CARRY(( (din_a[4] & din_b[0]) ) + ( Xd_0__inst_mult_0_394  ) + ( Xd_0__inst_mult_0_393  ))
// Xd_0__inst_mult_0_286  = SHARE((din_a[4] & din_b[1]))

	.dataa(!din_a[4]),
	.datab(!din_b[0]),
	.datac(!din_b[1]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_393 ),
	.sharein(Xd_0__inst_mult_0_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_284 ),
	.cout(Xd_0__inst_mult_0_285 ),
	.shareout(Xd_0__inst_mult_0_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_94 (
// Equation(s):
// Xd_0__inst_mult_0_288  = SUM(( (din_a[1] & din_b[3]) ) + ( Xd_0__inst_mult_0_402  ) + ( Xd_0__inst_mult_0_401  ))
// Xd_0__inst_mult_0_289  = CARRY(( (din_a[1] & din_b[3]) ) + ( Xd_0__inst_mult_0_402  ) + ( Xd_0__inst_mult_0_401  ))
// Xd_0__inst_mult_0_290  = SHARE((din_b[3] & din_a[2]))

	.dataa(!din_a[1]),
	.datab(!din_b[3]),
	.datac(!din_a[2]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_401 ),
	.sharein(Xd_0__inst_mult_0_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_288 ),
	.cout(Xd_0__inst_mult_0_289 ),
	.shareout(Xd_0__inst_mult_0_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_89 (
// Equation(s):
// Xd_0__inst_mult_1_268  = SUM(( (din_a[16] & din_b[12]) ) + ( Xd_0__inst_mult_1_175  ) + ( Xd_0__inst_mult_1_174  ))
// Xd_0__inst_mult_1_269  = CARRY(( (din_a[16] & din_b[12]) ) + ( Xd_0__inst_mult_1_175  ) + ( Xd_0__inst_mult_1_174  ))
// Xd_0__inst_mult_1_270  = SHARE((din_a[16] & din_b[13]))

	.dataa(!din_a[16]),
	.datab(!din_b[12]),
	.datac(!din_b[13]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_174 ),
	.sharein(Xd_0__inst_mult_1_175 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_268 ),
	.cout(Xd_0__inst_mult_1_269 ),
	.shareout(Xd_0__inst_mult_1_270 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_90 (
// Equation(s):
// Xd_0__inst_mult_1_272  = SUM(( (din_a[13] & din_b[15]) ) + ( Xd_0__inst_mult_1_386  ) + ( Xd_0__inst_mult_1_385  ))
// Xd_0__inst_mult_1_273  = CARRY(( (din_a[13] & din_b[15]) ) + ( Xd_0__inst_mult_1_386  ) + ( Xd_0__inst_mult_1_385  ))
// Xd_0__inst_mult_1_274  = SHARE((din_b[15] & din_a[14]))

	.dataa(!din_a[13]),
	.datab(!din_b[15]),
	.datac(!din_a[14]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_385 ),
	.sharein(Xd_0__inst_mult_1_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_272 ),
	.cout(Xd_0__inst_mult_1_273 ),
	.shareout(Xd_0__inst_mult_1_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_124 (
// Equation(s):
// Xd_0__inst_mult_6_397  = CARRY(( (din_a[75] & din_b[73]) ) + ( Xd_0__inst_mult_6_550  ) + ( Xd_0__inst_mult_6_549  ))
// Xd_0__inst_mult_6_398  = SHARE((din_a[74] & din_b[74]))

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(!din_a[74]),
	.datad(!din_b[74]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_549 ),
	.sharein(Xd_0__inst_mult_6_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_397 ),
	.shareout(Xd_0__inst_mult_6_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_126 (
// Equation(s):
// Xd_0__inst_mult_7_405  = CARRY(( (din_a[87] & din_b[85]) ) + ( Xd_0__inst_mult_7_574  ) + ( Xd_0__inst_mult_7_573  ))
// Xd_0__inst_mult_7_406  = SHARE((din_a[86] & din_b[86]))

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(!din_a[86]),
	.datad(!din_b[86]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_573 ),
	.sharein(Xd_0__inst_mult_7_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_405 ),
	.shareout(Xd_0__inst_mult_7_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_93 (
// Equation(s):
// Xd_0__inst_mult_4_272  = SUM(( !Xd_0__inst_mult_4_396  $ (!Xd_0__inst_mult_4_400  $ (((din_b[52] & din_a[49])))) ) + ( Xd_0__inst_mult_4_258  ) + ( Xd_0__inst_mult_4_257  ))
// Xd_0__inst_mult_4_273  = CARRY(( !Xd_0__inst_mult_4_396  $ (!Xd_0__inst_mult_4_400  $ (((din_b[52] & din_a[49])))) ) + ( Xd_0__inst_mult_4_258  ) + ( Xd_0__inst_mult_4_257  ))
// Xd_0__inst_mult_4_274  = SHARE((!Xd_0__inst_mult_4_396  & (Xd_0__inst_mult_4_400  & (din_b[52] & din_a[49]))) # (Xd_0__inst_mult_4_396  & (((din_b[52] & din_a[49])) # (Xd_0__inst_mult_4_400 ))))

	.dataa(!Xd_0__inst_mult_4_396 ),
	.datab(!Xd_0__inst_mult_4_400 ),
	.datac(!din_b[52]),
	.datad(!din_a[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_257 ),
	.sharein(Xd_0__inst_mult_4_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_272 ),
	.cout(Xd_0__inst_mult_4_273 ),
	.shareout(Xd_0__inst_mult_4_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_94 (
// Equation(s):
// Xd_0__inst_mult_4_276  = SUM(( (din_a[48] & din_b[53]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_277  = CARRY(( (din_a[48] & din_b[53]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_278  = SHARE((din_a[48] & din_b[54]))

	.dataa(!din_a[48]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_276 ),
	.cout(Xd_0__inst_mult_4_277 ),
	.shareout(Xd_0__inst_mult_4_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_35 (
// Equation(s):
// Xd_0__inst_mult_5_35_sumout  = SUM(( (din_a[69] & din_b[60]) ) + ( Xd_0__inst_mult_0_61  ) + ( Xd_0__inst_mult_0_60  ))
// Xd_0__inst_mult_5_36  = CARRY(( (din_a[69] & din_b[60]) ) + ( Xd_0__inst_mult_0_61  ) + ( Xd_0__inst_mult_0_60  ))
// Xd_0__inst_mult_5_37  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_60 ),
	.sharein(Xd_0__inst_mult_0_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_35_sumout ),
	.cout(Xd_0__inst_mult_5_36 ),
	.shareout(Xd_0__inst_mult_5_37 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_93 (
// Equation(s):
// Xd_0__inst_mult_5_272  = SUM(( !Xd_0__inst_mult_5_392  $ (!Xd_0__inst_mult_5_396  $ (((din_b[64] & din_a[61])))) ) + ( Xd_0__inst_mult_5_258  ) + ( Xd_0__inst_mult_5_257  ))
// Xd_0__inst_mult_5_273  = CARRY(( !Xd_0__inst_mult_5_392  $ (!Xd_0__inst_mult_5_396  $ (((din_b[64] & din_a[61])))) ) + ( Xd_0__inst_mult_5_258  ) + ( Xd_0__inst_mult_5_257  ))
// Xd_0__inst_mult_5_274  = SHARE((!Xd_0__inst_mult_5_392  & (Xd_0__inst_mult_5_396  & (din_b[64] & din_a[61]))) # (Xd_0__inst_mult_5_392  & (((din_b[64] & din_a[61])) # (Xd_0__inst_mult_5_396 ))))

	.dataa(!Xd_0__inst_mult_5_392 ),
	.datab(!Xd_0__inst_mult_5_396 ),
	.datac(!din_b[64]),
	.datad(!din_a[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_257 ),
	.sharein(Xd_0__inst_mult_5_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_272 ),
	.cout(Xd_0__inst_mult_5_273 ),
	.shareout(Xd_0__inst_mult_5_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_94 (
// Equation(s):
// Xd_0__inst_mult_5_276  = SUM(( (din_a[60] & din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_277  = CARRY(( (din_a[60] & din_b[65]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_278  = SHARE((din_a[60] & din_b[66]))

	.dataa(!din_a[60]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_276 ),
	.cout(Xd_0__inst_mult_5_277 ),
	.shareout(Xd_0__inst_mult_5_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_47 (
// Equation(s):
// Xd_0__inst_mult_1_47_sumout  = SUM(( (din_a[22] & din_b[20]) ) + ( Xd_0__inst_mult_4_53  ) + ( Xd_0__inst_mult_4_52  ))
// Xd_0__inst_mult_1_48  = CARRY(( (din_a[22] & din_b[20]) ) + ( Xd_0__inst_mult_4_53  ) + ( Xd_0__inst_mult_4_52  ))
// Xd_0__inst_mult_1_49  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_52 ),
	.sharein(Xd_0__inst_mult_4_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_47_sumout ),
	.cout(Xd_0__inst_mult_1_48 ),
	.shareout(Xd_0__inst_mult_1_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_93 (
// Equation(s):
// Xd_0__inst_mult_2_272  = SUM(( !Xd_0__inst_mult_2_392  $ (!Xd_0__inst_mult_2_396  $ (((din_b[28] & din_a[25])))) ) + ( Xd_0__inst_mult_2_258  ) + ( Xd_0__inst_mult_2_257  ))
// Xd_0__inst_mult_2_273  = CARRY(( !Xd_0__inst_mult_2_392  $ (!Xd_0__inst_mult_2_396  $ (((din_b[28] & din_a[25])))) ) + ( Xd_0__inst_mult_2_258  ) + ( Xd_0__inst_mult_2_257  ))
// Xd_0__inst_mult_2_274  = SHARE((!Xd_0__inst_mult_2_392  & (Xd_0__inst_mult_2_396  & (din_b[28] & din_a[25]))) # (Xd_0__inst_mult_2_392  & (((din_b[28] & din_a[25])) # (Xd_0__inst_mult_2_396 ))))

	.dataa(!Xd_0__inst_mult_2_392 ),
	.datab(!Xd_0__inst_mult_2_396 ),
	.datac(!din_b[28]),
	.datad(!din_a[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_257 ),
	.sharein(Xd_0__inst_mult_2_258 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_272 ),
	.cout(Xd_0__inst_mult_2_273 ),
	.shareout(Xd_0__inst_mult_2_274 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_94 (
// Equation(s):
// Xd_0__inst_mult_2_276  = SUM(( (din_a[24] & din_b[29]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_277  = CARRY(( (din_a[24] & din_b[29]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_278  = SHARE((din_a[24] & din_b[30]))

	.dataa(!din_a[24]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_276 ),
	.cout(Xd_0__inst_mult_2_277 ),
	.shareout(Xd_0__inst_mult_2_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_39 (
// Equation(s):
// Xd_0__inst_mult_5_39_sumout  = SUM(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_3_49  ) + ( Xd_0__inst_mult_3_48  ))
// Xd_0__inst_mult_5_40  = CARRY(( (din_a[70] & din_b[69]) ) + ( Xd_0__inst_mult_3_49  ) + ( Xd_0__inst_mult_3_48  ))
// Xd_0__inst_mult_5_41  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[69]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_48 ),
	.sharein(Xd_0__inst_mult_3_49 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_39_sumout ),
	.cout(Xd_0__inst_mult_5_40 ),
	.shareout(Xd_0__inst_mult_5_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_101 (
// Equation(s):
// Xd_0__inst_mult_3_316  = SUM(( !Xd_0__inst_mult_3_432  $ (!Xd_0__inst_mult_3_436  $ (((din_b[40] & din_a[37])))) ) + ( Xd_0__inst_mult_3_290  ) + ( Xd_0__inst_mult_3_289  ))
// Xd_0__inst_mult_3_317  = CARRY(( !Xd_0__inst_mult_3_432  $ (!Xd_0__inst_mult_3_436  $ (((din_b[40] & din_a[37])))) ) + ( Xd_0__inst_mult_3_290  ) + ( Xd_0__inst_mult_3_289  ))
// Xd_0__inst_mult_3_318  = SHARE((!Xd_0__inst_mult_3_432  & (Xd_0__inst_mult_3_436  & (din_b[40] & din_a[37]))) # (Xd_0__inst_mult_3_432  & (((din_b[40] & din_a[37])) # (Xd_0__inst_mult_3_436 ))))

	.dataa(!Xd_0__inst_mult_3_432 ),
	.datab(!Xd_0__inst_mult_3_436 ),
	.datac(!din_b[40]),
	.datad(!din_a[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_289 ),
	.sharein(Xd_0__inst_mult_3_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_316 ),
	.cout(Xd_0__inst_mult_3_317 ),
	.shareout(Xd_0__inst_mult_3_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_102 (
// Equation(s):
// Xd_0__inst_mult_3_320  = SUM(( (din_a[36] & din_b[41]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_321  = CARRY(( (din_a[36] & din_b[41]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_322  = SHARE((din_a[36] & din_b[42]))

	.dataa(!din_a[36]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_320 ),
	.cout(Xd_0__inst_mult_3_321 ),
	.shareout(Xd_0__inst_mult_3_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_39 (
// Equation(s):
// Xd_0__inst_mult_0_39_sumout  = SUM(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_1_61  ) + ( Xd_0__inst_mult_1_60  ))
// Xd_0__inst_mult_0_40  = CARRY(( (din_a[10] & din_b[9]) ) + ( Xd_0__inst_mult_1_61  ) + ( Xd_0__inst_mult_1_60  ))
// Xd_0__inst_mult_0_41  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[9]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_60 ),
	.sharein(Xd_0__inst_mult_1_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_39_sumout ),
	.cout(Xd_0__inst_mult_0_40 ),
	.shareout(Xd_0__inst_mult_0_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_95 (
// Equation(s):
// Xd_0__inst_mult_0_292  = SUM(( !Xd_0__inst_mult_0_404  $ (!Xd_0__inst_mult_0_408  $ (((din_b[4] & din_a[1])))) ) + ( Xd_0__inst_mult_0_270  ) + ( Xd_0__inst_mult_0_269  ))
// Xd_0__inst_mult_0_293  = CARRY(( !Xd_0__inst_mult_0_404  $ (!Xd_0__inst_mult_0_408  $ (((din_b[4] & din_a[1])))) ) + ( Xd_0__inst_mult_0_270  ) + ( Xd_0__inst_mult_0_269  ))
// Xd_0__inst_mult_0_294  = SHARE((!Xd_0__inst_mult_0_404  & (Xd_0__inst_mult_0_408  & (din_b[4] & din_a[1]))) # (Xd_0__inst_mult_0_404  & (((din_b[4] & din_a[1])) # (Xd_0__inst_mult_0_408 ))))

	.dataa(!Xd_0__inst_mult_0_404 ),
	.datab(!Xd_0__inst_mult_0_408 ),
	.datac(!din_b[4]),
	.datad(!din_a[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_269 ),
	.sharein(Xd_0__inst_mult_0_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_292 ),
	.cout(Xd_0__inst_mult_0_293 ),
	.shareout(Xd_0__inst_mult_0_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_96 (
// Equation(s):
// Xd_0__inst_mult_0_296  = SUM(( (din_a[0] & din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_297  = CARRY(( (din_a[0] & din_b[5]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_298  = SHARE((din_a[0] & din_b[6]))

	.dataa(!din_a[0]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_296 ),
	.cout(Xd_0__inst_mult_0_297 ),
	.shareout(Xd_0__inst_mult_0_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_43 (
// Equation(s):
// Xd_0__inst_mult_5_43_sumout  = SUM(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_4_57  ) + ( Xd_0__inst_mult_4_56  ))
// Xd_0__inst_mult_5_44  = CARRY(( (din_a[70] & din_b[70]) ) + ( Xd_0__inst_mult_4_57  ) + ( Xd_0__inst_mult_4_56  ))
// Xd_0__inst_mult_5_45  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_56 ),
	.sharein(Xd_0__inst_mult_4_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_43_sumout ),
	.cout(Xd_0__inst_mult_5_44 ),
	.shareout(Xd_0__inst_mult_5_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_91 (
// Equation(s):
// Xd_0__inst_mult_1_276  = SUM(( !Xd_0__inst_mult_1_388  $ (!Xd_0__inst_mult_1_392  $ (((din_b[16] & din_a[13])))) ) + ( Xd_0__inst_mult_1_262  ) + ( Xd_0__inst_mult_1_261  ))
// Xd_0__inst_mult_1_277  = CARRY(( !Xd_0__inst_mult_1_388  $ (!Xd_0__inst_mult_1_392  $ (((din_b[16] & din_a[13])))) ) + ( Xd_0__inst_mult_1_262  ) + ( Xd_0__inst_mult_1_261  ))
// Xd_0__inst_mult_1_278  = SHARE((!Xd_0__inst_mult_1_388  & (Xd_0__inst_mult_1_392  & (din_b[16] & din_a[13]))) # (Xd_0__inst_mult_1_388  & (((din_b[16] & din_a[13])) # (Xd_0__inst_mult_1_392 ))))

	.dataa(!Xd_0__inst_mult_1_388 ),
	.datab(!Xd_0__inst_mult_1_392 ),
	.datac(!din_b[16]),
	.datad(!din_a[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_261 ),
	.sharein(Xd_0__inst_mult_1_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_276 ),
	.cout(Xd_0__inst_mult_1_277 ),
	.shareout(Xd_0__inst_mult_1_278 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_92 (
// Equation(s):
// Xd_0__inst_mult_1_280  = SUM(( (din_a[12] & din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_281  = CARRY(( (din_a[12] & din_b[17]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_282  = SHARE((din_a[12] & din_b[18]))

	.dataa(!din_a[12]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_280 ),
	.cout(Xd_0__inst_mult_1_281 ),
	.shareout(Xd_0__inst_mult_1_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_43 (
// Equation(s):
// Xd_0__inst_mult_0_43_sumout  = SUM(( (din_a[10] & din_b[10]) ) + ( Xd_0__inst_mult_3_57  ) + ( Xd_0__inst_mult_3_56  ))
// Xd_0__inst_mult_0_44  = CARRY(( (din_a[10] & din_b[10]) ) + ( Xd_0__inst_mult_3_57  ) + ( Xd_0__inst_mult_3_56  ))
// Xd_0__inst_mult_0_45  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_56 ),
	.sharein(Xd_0__inst_mult_3_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_43_sumout ),
	.cout(Xd_0__inst_mult_0_44 ),
	.shareout(Xd_0__inst_mult_0_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_125 (
// Equation(s):
// Xd_0__inst_mult_6_400  = SUM(( (din_a[77] & din_b[72]) ) + ( Xd_0__inst_mult_6_282  ) + ( Xd_0__inst_mult_6_281  ))
// Xd_0__inst_mult_6_401  = CARRY(( (din_a[77] & din_b[72]) ) + ( Xd_0__inst_mult_6_282  ) + ( Xd_0__inst_mult_6_281  ))
// Xd_0__inst_mult_6_402  = SHARE((din_b[72] & din_a[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[72]),
	.datac(!din_a[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_281 ),
	.sharein(Xd_0__inst_mult_6_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_400 ),
	.cout(Xd_0__inst_mult_6_401 ),
	.shareout(Xd_0__inst_mult_6_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_126 (
// Equation(s):
// Xd_0__inst_mult_6_404  = SUM(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_6_286  ) + ( Xd_0__inst_mult_6_285  ))
// Xd_0__inst_mult_6_405  = CARRY(( (din_a[75] & din_b[74]) ) + ( Xd_0__inst_mult_6_286  ) + ( Xd_0__inst_mult_6_285  ))
// Xd_0__inst_mult_6_406  = SHARE((din_b[74] & din_a[76]))

	.dataa(!din_a[75]),
	.datab(!din_b[74]),
	.datac(!din_a[76]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_285 ),
	.sharein(Xd_0__inst_mult_6_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_404 ),
	.cout(Xd_0__inst_mult_6_405 ),
	.shareout(Xd_0__inst_mult_6_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_47 (
// Equation(s):
// Xd_0__inst_mult_0_47_sumout  = SUM(( (din_a[9] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_48  = CARRY(( (din_a[9] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_49  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_47_sumout ),
	.cout(Xd_0__inst_mult_0_48 ),
	.shareout(Xd_0__inst_mult_0_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_127 (
// Equation(s):
// Xd_0__inst_mult_7_408  = SUM(( (din_a[89] & din_b[84]) ) + ( Xd_0__inst_mult_7_290  ) + ( Xd_0__inst_mult_7_289  ))
// Xd_0__inst_mult_7_409  = CARRY(( (din_a[89] & din_b[84]) ) + ( Xd_0__inst_mult_7_290  ) + ( Xd_0__inst_mult_7_289  ))
// Xd_0__inst_mult_7_410  = SHARE((din_b[84] & din_a[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[84]),
	.datac(!din_a[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_289 ),
	.sharein(Xd_0__inst_mult_7_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_408 ),
	.cout(Xd_0__inst_mult_7_409 ),
	.shareout(Xd_0__inst_mult_7_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_128 (
// Equation(s):
// Xd_0__inst_mult_7_412  = SUM(( (din_a[87] & din_b[86]) ) + ( Xd_0__inst_mult_7_294  ) + ( Xd_0__inst_mult_7_293  ))
// Xd_0__inst_mult_7_413  = CARRY(( (din_a[87] & din_b[86]) ) + ( Xd_0__inst_mult_7_294  ) + ( Xd_0__inst_mult_7_293  ))
// Xd_0__inst_mult_7_414  = SHARE((din_b[86] & din_a[88]))

	.dataa(!din_a[87]),
	.datab(!din_b[86]),
	.datac(!din_a[88]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_293 ),
	.sharein(Xd_0__inst_mult_7_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_412 ),
	.cout(Xd_0__inst_mult_7_413 ),
	.shareout(Xd_0__inst_mult_7_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_47 (
// Equation(s):
// Xd_0__inst_mult_5_47_sumout  = SUM(( (din_a[70] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_48  = CARRY(( (din_a[70] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_49  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_47_sumout ),
	.cout(Xd_0__inst_mult_5_48 ),
	.shareout(Xd_0__inst_mult_5_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_95 (
// Equation(s):
// Xd_0__inst_mult_4_280  = SUM(( !Xd_0__inst_mult_4_404  $ (!Xd_0__inst_mult_4_408 ) ) + ( Xd_0__inst_mult_4_274  ) + ( Xd_0__inst_mult_4_273  ))
// Xd_0__inst_mult_4_281  = CARRY(( !Xd_0__inst_mult_4_404  $ (!Xd_0__inst_mult_4_408 ) ) + ( Xd_0__inst_mult_4_274  ) + ( Xd_0__inst_mult_4_273  ))
// Xd_0__inst_mult_4_282  = SHARE((Xd_0__inst_mult_4_404  & Xd_0__inst_mult_4_408 ))

	.dataa(!Xd_0__inst_mult_4_404 ),
	.datab(!Xd_0__inst_mult_4_408 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_273 ),
	.sharein(Xd_0__inst_mult_4_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_280 ),
	.cout(Xd_0__inst_mult_4_281 ),
	.shareout(Xd_0__inst_mult_4_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_96 (
// Equation(s):
// Xd_0__inst_mult_4_284  = SUM(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_4_278  ) + ( Xd_0__inst_mult_4_277  ))
// Xd_0__inst_mult_4_285  = CARRY(( (din_a[49] & din_b[53]) ) + ( Xd_0__inst_mult_4_278  ) + ( Xd_0__inst_mult_4_277  ))
// Xd_0__inst_mult_4_286  = SHARE((din_a[48] & din_b[55]))

	.dataa(!din_a[49]),
	.datab(!din_b[53]),
	.datac(!din_a[48]),
	.datad(!din_b[55]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_277 ),
	.sharein(Xd_0__inst_mult_4_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_284 ),
	.cout(Xd_0__inst_mult_4_285 ),
	.shareout(Xd_0__inst_mult_4_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_95 (
// Equation(s):
// Xd_0__inst_mult_5_280  = SUM(( !Xd_0__inst_mult_5_400  $ (!Xd_0__inst_mult_5_404 ) ) + ( Xd_0__inst_mult_5_274  ) + ( Xd_0__inst_mult_5_273  ))
// Xd_0__inst_mult_5_281  = CARRY(( !Xd_0__inst_mult_5_400  $ (!Xd_0__inst_mult_5_404 ) ) + ( Xd_0__inst_mult_5_274  ) + ( Xd_0__inst_mult_5_273  ))
// Xd_0__inst_mult_5_282  = SHARE((Xd_0__inst_mult_5_400  & Xd_0__inst_mult_5_404 ))

	.dataa(!Xd_0__inst_mult_5_400 ),
	.datab(!Xd_0__inst_mult_5_404 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_273 ),
	.sharein(Xd_0__inst_mult_5_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_280 ),
	.cout(Xd_0__inst_mult_5_281 ),
	.shareout(Xd_0__inst_mult_5_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_96 (
// Equation(s):
// Xd_0__inst_mult_5_284  = SUM(( (din_a[61] & din_b[65]) ) + ( Xd_0__inst_mult_5_278  ) + ( Xd_0__inst_mult_5_277  ))
// Xd_0__inst_mult_5_285  = CARRY(( (din_a[61] & din_b[65]) ) + ( Xd_0__inst_mult_5_278  ) + ( Xd_0__inst_mult_5_277  ))
// Xd_0__inst_mult_5_286  = SHARE((din_a[60] & din_b[67]))

	.dataa(!din_a[61]),
	.datab(!din_b[65]),
	.datac(!din_a[60]),
	.datad(!din_b[67]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_277 ),
	.sharein(Xd_0__inst_mult_5_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_284 ),
	.cout(Xd_0__inst_mult_5_285 ),
	.shareout(Xd_0__inst_mult_5_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_95 (
// Equation(s):
// Xd_0__inst_mult_2_280  = SUM(( !Xd_0__inst_mult_2_400  $ (!Xd_0__inst_mult_2_404 ) ) + ( Xd_0__inst_mult_2_274  ) + ( Xd_0__inst_mult_2_273  ))
// Xd_0__inst_mult_2_281  = CARRY(( !Xd_0__inst_mult_2_400  $ (!Xd_0__inst_mult_2_404 ) ) + ( Xd_0__inst_mult_2_274  ) + ( Xd_0__inst_mult_2_273  ))
// Xd_0__inst_mult_2_282  = SHARE((Xd_0__inst_mult_2_400  & Xd_0__inst_mult_2_404 ))

	.dataa(!Xd_0__inst_mult_2_400 ),
	.datab(!Xd_0__inst_mult_2_404 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_273 ),
	.sharein(Xd_0__inst_mult_2_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_280 ),
	.cout(Xd_0__inst_mult_2_281 ),
	.shareout(Xd_0__inst_mult_2_282 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_96 (
// Equation(s):
// Xd_0__inst_mult_2_284  = SUM(( (din_a[25] & din_b[29]) ) + ( Xd_0__inst_mult_2_278  ) + ( Xd_0__inst_mult_2_277  ))
// Xd_0__inst_mult_2_285  = CARRY(( (din_a[25] & din_b[29]) ) + ( Xd_0__inst_mult_2_278  ) + ( Xd_0__inst_mult_2_277  ))
// Xd_0__inst_mult_2_286  = SHARE((din_a[24] & din_b[31]))

	.dataa(!din_a[25]),
	.datab(!din_b[29]),
	.datac(!din_a[24]),
	.datad(!din_b[31]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_277 ),
	.sharein(Xd_0__inst_mult_2_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_284 ),
	.cout(Xd_0__inst_mult_2_285 ),
	.shareout(Xd_0__inst_mult_2_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_103 (
// Equation(s):
// Xd_0__inst_mult_3_324  = SUM(( !Xd_0__inst_mult_3_440  $ (!Xd_0__inst_mult_3_444 ) ) + ( Xd_0__inst_mult_3_318  ) + ( Xd_0__inst_mult_3_317  ))
// Xd_0__inst_mult_3_325  = CARRY(( !Xd_0__inst_mult_3_440  $ (!Xd_0__inst_mult_3_444 ) ) + ( Xd_0__inst_mult_3_318  ) + ( Xd_0__inst_mult_3_317  ))
// Xd_0__inst_mult_3_326  = SHARE((Xd_0__inst_mult_3_440  & Xd_0__inst_mult_3_444 ))

	.dataa(!Xd_0__inst_mult_3_440 ),
	.datab(!Xd_0__inst_mult_3_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_317 ),
	.sharein(Xd_0__inst_mult_3_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_324 ),
	.cout(Xd_0__inst_mult_3_325 ),
	.shareout(Xd_0__inst_mult_3_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_104 (
// Equation(s):
// Xd_0__inst_mult_3_328  = SUM(( (din_a[37] & din_b[41]) ) + ( Xd_0__inst_mult_3_322  ) + ( Xd_0__inst_mult_3_321  ))
// Xd_0__inst_mult_3_329  = CARRY(( (din_a[37] & din_b[41]) ) + ( Xd_0__inst_mult_3_322  ) + ( Xd_0__inst_mult_3_321  ))
// Xd_0__inst_mult_3_330  = SHARE((din_a[36] & din_b[43]))

	.dataa(!din_a[37]),
	.datab(!din_b[41]),
	.datac(!din_a[36]),
	.datad(!din_b[43]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_321 ),
	.sharein(Xd_0__inst_mult_3_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_328 ),
	.cout(Xd_0__inst_mult_3_329 ),
	.shareout(Xd_0__inst_mult_3_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_97 (
// Equation(s):
// Xd_0__inst_mult_0_300  = SUM(( !Xd_0__inst_mult_0_412  $ (!Xd_0__inst_mult_0_416 ) ) + ( Xd_0__inst_mult_0_294  ) + ( Xd_0__inst_mult_0_293  ))
// Xd_0__inst_mult_0_301  = CARRY(( !Xd_0__inst_mult_0_412  $ (!Xd_0__inst_mult_0_416 ) ) + ( Xd_0__inst_mult_0_294  ) + ( Xd_0__inst_mult_0_293  ))
// Xd_0__inst_mult_0_302  = SHARE((Xd_0__inst_mult_0_412  & Xd_0__inst_mult_0_416 ))

	.dataa(!Xd_0__inst_mult_0_412 ),
	.datab(!Xd_0__inst_mult_0_416 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_293 ),
	.sharein(Xd_0__inst_mult_0_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_300 ),
	.cout(Xd_0__inst_mult_0_301 ),
	.shareout(Xd_0__inst_mult_0_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_98 (
// Equation(s):
// Xd_0__inst_mult_0_304  = SUM(( (din_a[1] & din_b[5]) ) + ( Xd_0__inst_mult_0_298  ) + ( Xd_0__inst_mult_0_297  ))
// Xd_0__inst_mult_0_305  = CARRY(( (din_a[1] & din_b[5]) ) + ( Xd_0__inst_mult_0_298  ) + ( Xd_0__inst_mult_0_297  ))
// Xd_0__inst_mult_0_306  = SHARE((din_a[0] & din_b[7]))

	.dataa(!din_a[1]),
	.datab(!din_b[5]),
	.datac(!din_a[0]),
	.datad(!din_b[7]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_297 ),
	.sharein(Xd_0__inst_mult_0_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_304 ),
	.cout(Xd_0__inst_mult_0_305 ),
	.shareout(Xd_0__inst_mult_0_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_93 (
// Equation(s):
// Xd_0__inst_mult_1_284  = SUM(( !Xd_0__inst_mult_1_396  $ (!Xd_0__inst_mult_1_400 ) ) + ( Xd_0__inst_mult_1_278  ) + ( Xd_0__inst_mult_1_277  ))
// Xd_0__inst_mult_1_285  = CARRY(( !Xd_0__inst_mult_1_396  $ (!Xd_0__inst_mult_1_400 ) ) + ( Xd_0__inst_mult_1_278  ) + ( Xd_0__inst_mult_1_277  ))
// Xd_0__inst_mult_1_286  = SHARE((Xd_0__inst_mult_1_396  & Xd_0__inst_mult_1_400 ))

	.dataa(!Xd_0__inst_mult_1_396 ),
	.datab(!Xd_0__inst_mult_1_400 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_277 ),
	.sharein(Xd_0__inst_mult_1_278 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_284 ),
	.cout(Xd_0__inst_mult_1_285 ),
	.shareout(Xd_0__inst_mult_1_286 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_94 (
// Equation(s):
// Xd_0__inst_mult_1_288  = SUM(( (din_a[13] & din_b[17]) ) + ( Xd_0__inst_mult_1_282  ) + ( Xd_0__inst_mult_1_281  ))
// Xd_0__inst_mult_1_289  = CARRY(( (din_a[13] & din_b[17]) ) + ( Xd_0__inst_mult_1_282  ) + ( Xd_0__inst_mult_1_281  ))
// Xd_0__inst_mult_1_290  = SHARE((din_a[12] & din_b[19]))

	.dataa(!din_a[13]),
	.datab(!din_b[17]),
	.datac(!din_a[12]),
	.datad(!din_b[19]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_281 ),
	.sharein(Xd_0__inst_mult_1_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_288 ),
	.cout(Xd_0__inst_mult_1_289 ),
	.shareout(Xd_0__inst_mult_1_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_127 (
// Equation(s):
// Xd_0__inst_mult_6_408  = SUM(( (din_a[77] & din_b[73]) ) + ( Xd_0__inst_mult_6_402  ) + ( Xd_0__inst_mult_6_401  ))
// Xd_0__inst_mult_6_409  = CARRY(( (din_a[77] & din_b[73]) ) + ( Xd_0__inst_mult_6_402  ) + ( Xd_0__inst_mult_6_401  ))
// Xd_0__inst_mult_6_410  = SHARE((din_b[73] & din_a[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[73]),
	.datac(!din_a[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_401 ),
	.sharein(Xd_0__inst_mult_6_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_408 ),
	.cout(Xd_0__inst_mult_6_409 ),
	.shareout(Xd_0__inst_mult_6_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_128 (
// Equation(s):
// Xd_0__inst_mult_6_412  = SUM(( (!din_a[75] & (((din_a[74] & din_b[76])))) # (din_a[75] & (!din_b[75] $ (((!din_a[74]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_406  ) + ( Xd_0__inst_mult_6_405  ))
// Xd_0__inst_mult_6_413  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[76])))) # (din_a[75] & (!din_b[75] $ (((!din_a[74]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_406  ) + ( Xd_0__inst_mult_6_405  ))
// Xd_0__inst_mult_6_414  = SHARE((din_a[75] & (din_b[75] & (din_a[74] & din_b[76]))))

	.dataa(!din_a[75]),
	.datab(!din_b[75]),
	.datac(!din_a[74]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_405 ),
	.sharein(Xd_0__inst_mult_6_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_412 ),
	.cout(Xd_0__inst_mult_6_413 ),
	.shareout(Xd_0__inst_mult_6_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_129 (
// Equation(s):
// Xd_0__inst_mult_7_416  = SUM(( (din_a[89] & din_b[85]) ) + ( Xd_0__inst_mult_7_410  ) + ( Xd_0__inst_mult_7_409  ))
// Xd_0__inst_mult_7_417  = CARRY(( (din_a[89] & din_b[85]) ) + ( Xd_0__inst_mult_7_410  ) + ( Xd_0__inst_mult_7_409  ))
// Xd_0__inst_mult_7_418  = SHARE((din_b[85] & din_a[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[85]),
	.datac(!din_a[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_409 ),
	.sharein(Xd_0__inst_mult_7_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_416 ),
	.cout(Xd_0__inst_mult_7_417 ),
	.shareout(Xd_0__inst_mult_7_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_130 (
// Equation(s):
// Xd_0__inst_mult_7_420  = SUM(( (!din_a[87] & (((din_a[86] & din_b[88])))) # (din_a[87] & (!din_b[87] $ (((!din_a[86]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_414  ) + ( Xd_0__inst_mult_7_413  ))
// Xd_0__inst_mult_7_421  = CARRY(( (!din_a[87] & (((din_a[86] & din_b[88])))) # (din_a[87] & (!din_b[87] $ (((!din_a[86]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_414  ) + ( Xd_0__inst_mult_7_413  ))
// Xd_0__inst_mult_7_422  = SHARE((din_a[87] & (din_b[87] & (din_a[86] & din_b[88]))))

	.dataa(!din_a[87]),
	.datab(!din_b[87]),
	.datac(!din_a[86]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_413 ),
	.sharein(Xd_0__inst_mult_7_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_420 ),
	.cout(Xd_0__inst_mult_7_421 ),
	.shareout(Xd_0__inst_mult_7_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_97 (
// Equation(s):
// Xd_0__inst_mult_4_288  = SUM(( !Xd_0__inst_mult_4_412  $ (!Xd_0__inst_mult_4_416  $ (Xd_0__inst_mult_4_59_sumout )) ) + ( Xd_0__inst_mult_4_282  ) + ( Xd_0__inst_mult_4_281  ))
// Xd_0__inst_mult_4_289  = CARRY(( !Xd_0__inst_mult_4_412  $ (!Xd_0__inst_mult_4_416  $ (Xd_0__inst_mult_4_59_sumout )) ) + ( Xd_0__inst_mult_4_282  ) + ( Xd_0__inst_mult_4_281  ))
// Xd_0__inst_mult_4_290  = SHARE((!Xd_0__inst_mult_4_412  & (Xd_0__inst_mult_4_416  & Xd_0__inst_mult_4_59_sumout )) # (Xd_0__inst_mult_4_412  & ((Xd_0__inst_mult_4_59_sumout ) # (Xd_0__inst_mult_4_416 ))))

	.dataa(!Xd_0__inst_mult_4_412 ),
	.datab(!Xd_0__inst_mult_4_416 ),
	.datac(!Xd_0__inst_mult_4_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_281 ),
	.sharein(Xd_0__inst_mult_4_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_288 ),
	.cout(Xd_0__inst_mult_4_289 ),
	.shareout(Xd_0__inst_mult_4_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_98 (
// Equation(s):
// Xd_0__inst_mult_4_292  = SUM(( (!din_a[49] & (((din_a[50] & din_b[53])))) # (din_a[49] & (!din_b[54] $ (((!din_a[50]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_286  ) + ( Xd_0__inst_mult_4_285  ))
// Xd_0__inst_mult_4_293  = CARRY(( (!din_a[49] & (((din_a[50] & din_b[53])))) # (din_a[49] & (!din_b[54] $ (((!din_a[50]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_286  ) + ( Xd_0__inst_mult_4_285  ))
// Xd_0__inst_mult_4_294  = SHARE((din_a[49] & (din_b[54] & (din_a[50] & din_b[53]))))

	.dataa(!din_a[49]),
	.datab(!din_b[54]),
	.datac(!din_a[50]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_285 ),
	.sharein(Xd_0__inst_mult_4_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_292 ),
	.cout(Xd_0__inst_mult_4_293 ),
	.shareout(Xd_0__inst_mult_4_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_97 (
// Equation(s):
// Xd_0__inst_mult_5_288  = SUM(( !Xd_0__inst_mult_5_408  $ (!Xd_0__inst_mult_5_412  $ (Xd_0__inst_mult_5_63_sumout )) ) + ( Xd_0__inst_mult_5_282  ) + ( Xd_0__inst_mult_5_281  ))
// Xd_0__inst_mult_5_289  = CARRY(( !Xd_0__inst_mult_5_408  $ (!Xd_0__inst_mult_5_412  $ (Xd_0__inst_mult_5_63_sumout )) ) + ( Xd_0__inst_mult_5_282  ) + ( Xd_0__inst_mult_5_281  ))
// Xd_0__inst_mult_5_290  = SHARE((!Xd_0__inst_mult_5_408  & (Xd_0__inst_mult_5_412  & Xd_0__inst_mult_5_63_sumout )) # (Xd_0__inst_mult_5_408  & ((Xd_0__inst_mult_5_63_sumout ) # (Xd_0__inst_mult_5_412 ))))

	.dataa(!Xd_0__inst_mult_5_408 ),
	.datab(!Xd_0__inst_mult_5_412 ),
	.datac(!Xd_0__inst_mult_5_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_281 ),
	.sharein(Xd_0__inst_mult_5_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_288 ),
	.cout(Xd_0__inst_mult_5_289 ),
	.shareout(Xd_0__inst_mult_5_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_98 (
// Equation(s):
// Xd_0__inst_mult_5_292  = SUM(( (!din_a[61] & (((din_a[62] & din_b[65])))) # (din_a[61] & (!din_b[66] $ (((!din_a[62]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_286  ) + ( Xd_0__inst_mult_5_285  ))
// Xd_0__inst_mult_5_293  = CARRY(( (!din_a[61] & (((din_a[62] & din_b[65])))) # (din_a[61] & (!din_b[66] $ (((!din_a[62]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_286  ) + ( Xd_0__inst_mult_5_285  ))
// Xd_0__inst_mult_5_294  = SHARE((din_a[61] & (din_b[66] & (din_a[62] & din_b[65]))))

	.dataa(!din_a[61]),
	.datab(!din_b[66]),
	.datac(!din_a[62]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_285 ),
	.sharein(Xd_0__inst_mult_5_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_292 ),
	.cout(Xd_0__inst_mult_5_293 ),
	.shareout(Xd_0__inst_mult_5_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_97 (
// Equation(s):
// Xd_0__inst_mult_2_288  = SUM(( !Xd_0__inst_mult_2_408  $ (!Xd_0__inst_mult_2_412  $ (Xd_0__inst_mult_2_59_sumout )) ) + ( Xd_0__inst_mult_2_282  ) + ( Xd_0__inst_mult_2_281  ))
// Xd_0__inst_mult_2_289  = CARRY(( !Xd_0__inst_mult_2_408  $ (!Xd_0__inst_mult_2_412  $ (Xd_0__inst_mult_2_59_sumout )) ) + ( Xd_0__inst_mult_2_282  ) + ( Xd_0__inst_mult_2_281  ))
// Xd_0__inst_mult_2_290  = SHARE((!Xd_0__inst_mult_2_408  & (Xd_0__inst_mult_2_412  & Xd_0__inst_mult_2_59_sumout )) # (Xd_0__inst_mult_2_408  & ((Xd_0__inst_mult_2_59_sumout ) # (Xd_0__inst_mult_2_412 ))))

	.dataa(!Xd_0__inst_mult_2_408 ),
	.datab(!Xd_0__inst_mult_2_412 ),
	.datac(!Xd_0__inst_mult_2_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_281 ),
	.sharein(Xd_0__inst_mult_2_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_288 ),
	.cout(Xd_0__inst_mult_2_289 ),
	.shareout(Xd_0__inst_mult_2_290 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_98 (
// Equation(s):
// Xd_0__inst_mult_2_292  = SUM(( (!din_a[25] & (((din_a[26] & din_b[29])))) # (din_a[25] & (!din_b[30] $ (((!din_a[26]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_286  ) + ( Xd_0__inst_mult_2_285  ))
// Xd_0__inst_mult_2_293  = CARRY(( (!din_a[25] & (((din_a[26] & din_b[29])))) # (din_a[25] & (!din_b[30] $ (((!din_a[26]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_286  ) + ( Xd_0__inst_mult_2_285  ))
// Xd_0__inst_mult_2_294  = SHARE((din_a[25] & (din_b[30] & (din_a[26] & din_b[29]))))

	.dataa(!din_a[25]),
	.datab(!din_b[30]),
	.datac(!din_a[26]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_285 ),
	.sharein(Xd_0__inst_mult_2_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_292 ),
	.cout(Xd_0__inst_mult_2_293 ),
	.shareout(Xd_0__inst_mult_2_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_105 (
// Equation(s):
// Xd_0__inst_mult_3_332  = SUM(( !Xd_0__inst_mult_3_448  $ (!Xd_0__inst_mult_3_452  $ (Xd_0__inst_mult_3_59_sumout )) ) + ( Xd_0__inst_mult_3_326  ) + ( Xd_0__inst_mult_3_325  ))
// Xd_0__inst_mult_3_333  = CARRY(( !Xd_0__inst_mult_3_448  $ (!Xd_0__inst_mult_3_452  $ (Xd_0__inst_mult_3_59_sumout )) ) + ( Xd_0__inst_mult_3_326  ) + ( Xd_0__inst_mult_3_325  ))
// Xd_0__inst_mult_3_334  = SHARE((!Xd_0__inst_mult_3_448  & (Xd_0__inst_mult_3_452  & Xd_0__inst_mult_3_59_sumout )) # (Xd_0__inst_mult_3_448  & ((Xd_0__inst_mult_3_59_sumout ) # (Xd_0__inst_mult_3_452 ))))

	.dataa(!Xd_0__inst_mult_3_448 ),
	.datab(!Xd_0__inst_mult_3_452 ),
	.datac(!Xd_0__inst_mult_3_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_325 ),
	.sharein(Xd_0__inst_mult_3_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_332 ),
	.cout(Xd_0__inst_mult_3_333 ),
	.shareout(Xd_0__inst_mult_3_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_106 (
// Equation(s):
// Xd_0__inst_mult_3_336  = SUM(( (!din_a[37] & (((din_a[38] & din_b[41])))) # (din_a[37] & (!din_b[42] $ (((!din_a[38]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_330  ) + ( Xd_0__inst_mult_3_329  ))
// Xd_0__inst_mult_3_337  = CARRY(( (!din_a[37] & (((din_a[38] & din_b[41])))) # (din_a[37] & (!din_b[42] $ (((!din_a[38]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_330  ) + ( Xd_0__inst_mult_3_329  ))
// Xd_0__inst_mult_3_338  = SHARE((din_a[37] & (din_b[42] & (din_a[38] & din_b[41]))))

	.dataa(!din_a[37]),
	.datab(!din_b[42]),
	.datac(!din_a[38]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_329 ),
	.sharein(Xd_0__inst_mult_3_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_336 ),
	.cout(Xd_0__inst_mult_3_337 ),
	.shareout(Xd_0__inst_mult_3_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_99 (
// Equation(s):
// Xd_0__inst_mult_0_308  = SUM(( !Xd_0__inst_mult_0_420  $ (!Xd_0__inst_mult_0_424  $ (Xd_0__inst_mult_0_63_sumout )) ) + ( Xd_0__inst_mult_0_302  ) + ( Xd_0__inst_mult_0_301  ))
// Xd_0__inst_mult_0_309  = CARRY(( !Xd_0__inst_mult_0_420  $ (!Xd_0__inst_mult_0_424  $ (Xd_0__inst_mult_0_63_sumout )) ) + ( Xd_0__inst_mult_0_302  ) + ( Xd_0__inst_mult_0_301  ))
// Xd_0__inst_mult_0_310  = SHARE((!Xd_0__inst_mult_0_420  & (Xd_0__inst_mult_0_424  & Xd_0__inst_mult_0_63_sumout )) # (Xd_0__inst_mult_0_420  & ((Xd_0__inst_mult_0_63_sumout ) # (Xd_0__inst_mult_0_424 ))))

	.dataa(!Xd_0__inst_mult_0_420 ),
	.datab(!Xd_0__inst_mult_0_424 ),
	.datac(!Xd_0__inst_mult_0_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_301 ),
	.sharein(Xd_0__inst_mult_0_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_308 ),
	.cout(Xd_0__inst_mult_0_309 ),
	.shareout(Xd_0__inst_mult_0_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_100 (
// Equation(s):
// Xd_0__inst_mult_0_312  = SUM(( (!din_a[1] & (((din_a[2] & din_b[5])))) # (din_a[1] & (!din_b[6] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_306  ) + ( Xd_0__inst_mult_0_305  ))
// Xd_0__inst_mult_0_313  = CARRY(( (!din_a[1] & (((din_a[2] & din_b[5])))) # (din_a[1] & (!din_b[6] $ (((!din_a[2]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_306  ) + ( Xd_0__inst_mult_0_305  ))
// Xd_0__inst_mult_0_314  = SHARE((din_a[1] & (din_b[6] & (din_a[2] & din_b[5]))))

	.dataa(!din_a[1]),
	.datab(!din_b[6]),
	.datac(!din_a[2]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_305 ),
	.sharein(Xd_0__inst_mult_0_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_312 ),
	.cout(Xd_0__inst_mult_0_313 ),
	.shareout(Xd_0__inst_mult_0_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_95 (
// Equation(s):
// Xd_0__inst_mult_1_292  = SUM(( !Xd_0__inst_mult_1_404  $ (!Xd_0__inst_mult_1_408  $ (Xd_0__inst_mult_2_384 )) ) + ( Xd_0__inst_mult_1_286  ) + ( Xd_0__inst_mult_1_285  ))
// Xd_0__inst_mult_1_293  = CARRY(( !Xd_0__inst_mult_1_404  $ (!Xd_0__inst_mult_1_408  $ (Xd_0__inst_mult_2_384 )) ) + ( Xd_0__inst_mult_1_286  ) + ( Xd_0__inst_mult_1_285  ))
// Xd_0__inst_mult_1_294  = SHARE((!Xd_0__inst_mult_1_404  & (Xd_0__inst_mult_1_408  & Xd_0__inst_mult_2_384 )) # (Xd_0__inst_mult_1_404  & ((Xd_0__inst_mult_2_384 ) # (Xd_0__inst_mult_1_408 ))))

	.dataa(!Xd_0__inst_mult_1_404 ),
	.datab(!Xd_0__inst_mult_1_408 ),
	.datac(!Xd_0__inst_mult_2_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_285 ),
	.sharein(Xd_0__inst_mult_1_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_292 ),
	.cout(Xd_0__inst_mult_1_293 ),
	.shareout(Xd_0__inst_mult_1_294 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_96 (
// Equation(s):
// Xd_0__inst_mult_1_296  = SUM(( (!din_a[13] & (((din_a[14] & din_b[17])))) # (din_a[13] & (!din_b[18] $ (((!din_a[14]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_290  ) + ( Xd_0__inst_mult_1_289  ))
// Xd_0__inst_mult_1_297  = CARRY(( (!din_a[13] & (((din_a[14] & din_b[17])))) # (din_a[13] & (!din_b[18] $ (((!din_a[14]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_290  ) + ( Xd_0__inst_mult_1_289  ))
// Xd_0__inst_mult_1_298  = SHARE((din_a[13] & (din_b[18] & (din_a[14] & din_b[17]))))

	.dataa(!din_a[13]),
	.datab(!din_b[18]),
	.datac(!din_a[14]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_289 ),
	.sharein(Xd_0__inst_mult_1_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_296 ),
	.cout(Xd_0__inst_mult_1_297 ),
	.shareout(Xd_0__inst_mult_1_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_129 (
// Equation(s):
// Xd_0__inst_mult_6_416  = SUM(( (din_a[77] & din_b[74]) ) + ( Xd_0__inst_mult_6_410  ) + ( Xd_0__inst_mult_6_409  ))
// Xd_0__inst_mult_6_417  = CARRY(( (din_a[77] & din_b[74]) ) + ( Xd_0__inst_mult_6_410  ) + ( Xd_0__inst_mult_6_409  ))
// Xd_0__inst_mult_6_418  = SHARE((din_a[79] & din_b[73]))

	.dataa(!din_a[77]),
	.datab(!din_b[74]),
	.datac(!din_a[79]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_409 ),
	.sharein(Xd_0__inst_mult_6_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_416 ),
	.cout(Xd_0__inst_mult_6_417 ),
	.shareout(Xd_0__inst_mult_6_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_130 (
// Equation(s):
// Xd_0__inst_mult_6_420  = SUM(( (!din_a[76] & (((din_a[75] & din_b[76])))) # (din_a[76] & (!din_b[75] $ (((!din_a[75]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_414  ) + ( Xd_0__inst_mult_6_413  ))
// Xd_0__inst_mult_6_421  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[76])))) # (din_a[76] & (!din_b[75] $ (((!din_a[75]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_414  ) + ( Xd_0__inst_mult_6_413  ))
// Xd_0__inst_mult_6_422  = SHARE((din_a[76] & (din_b[75] & (din_a[75] & din_b[76]))))

	.dataa(!din_a[76]),
	.datab(!din_b[75]),
	.datac(!din_a[75]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_413 ),
	.sharein(Xd_0__inst_mult_6_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_420 ),
	.cout(Xd_0__inst_mult_6_421 ),
	.shareout(Xd_0__inst_mult_6_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_55 (
// Equation(s):
// Xd_0__inst_mult_6_55_sumout  = SUM(( (din_a[79] & din_b[72]) ) + ( Xd_0__inst_mult_7_53  ) + ( Xd_0__inst_mult_7_52  ))
// Xd_0__inst_mult_6_56  = CARRY(( (din_a[79] & din_b[72]) ) + ( Xd_0__inst_mult_7_53  ) + ( Xd_0__inst_mult_7_52  ))
// Xd_0__inst_mult_6_57  = SHARE(GND)

	.dataa(!din_a[79]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_52 ),
	.sharein(Xd_0__inst_mult_7_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_55_sumout ),
	.cout(Xd_0__inst_mult_6_56 ),
	.shareout(Xd_0__inst_mult_6_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_131 (
// Equation(s):
// Xd_0__inst_mult_7_424  = SUM(( (din_a[89] & din_b[86]) ) + ( Xd_0__inst_mult_7_418  ) + ( Xd_0__inst_mult_7_417  ))
// Xd_0__inst_mult_7_425  = CARRY(( (din_a[89] & din_b[86]) ) + ( Xd_0__inst_mult_7_418  ) + ( Xd_0__inst_mult_7_417  ))
// Xd_0__inst_mult_7_426  = SHARE((din_a[91] & din_b[85]))

	.dataa(!din_a[89]),
	.datab(!din_b[86]),
	.datac(!din_a[91]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_417 ),
	.sharein(Xd_0__inst_mult_7_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_424 ),
	.cout(Xd_0__inst_mult_7_425 ),
	.shareout(Xd_0__inst_mult_7_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_132 (
// Equation(s):
// Xd_0__inst_mult_7_428  = SUM(( (!din_a[88] & (((din_a[87] & din_b[88])))) # (din_a[88] & (!din_b[87] $ (((!din_a[87]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_422  ) + ( Xd_0__inst_mult_7_421  ))
// Xd_0__inst_mult_7_429  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[88])))) # (din_a[88] & (!din_b[87] $ (((!din_a[87]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_422  ) + ( Xd_0__inst_mult_7_421  ))
// Xd_0__inst_mult_7_430  = SHARE((din_a[88] & (din_b[87] & (din_a[87] & din_b[88]))))

	.dataa(!din_a[88]),
	.datab(!din_b[87]),
	.datac(!din_a[87]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_421 ),
	.sharein(Xd_0__inst_mult_7_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_428 ),
	.cout(Xd_0__inst_mult_7_429 ),
	.shareout(Xd_0__inst_mult_7_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_55 (
// Equation(s):
// Xd_0__inst_mult_7_55_sumout  = SUM(( (din_a[91] & din_b[84]) ) + ( Xd_0__inst_mult_6_37  ) + ( Xd_0__inst_mult_6_36  ))
// Xd_0__inst_mult_7_56  = CARRY(( (din_a[91] & din_b[84]) ) + ( Xd_0__inst_mult_6_37  ) + ( Xd_0__inst_mult_6_36  ))
// Xd_0__inst_mult_7_57  = SHARE(GND)

	.dataa(!din_a[91]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_36 ),
	.sharein(Xd_0__inst_mult_6_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_55_sumout ),
	.cout(Xd_0__inst_mult_7_56 ),
	.shareout(Xd_0__inst_mult_7_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_99 (
// Equation(s):
// Xd_0__inst_mult_4_296  = SUM(( !Xd_0__inst_mult_4_420  $ (!Xd_0__inst_mult_4_424  $ (Xd_0__inst_mult_4_63_sumout )) ) + ( Xd_0__inst_mult_4_290  ) + ( Xd_0__inst_mult_4_289  ))
// Xd_0__inst_mult_4_297  = CARRY(( !Xd_0__inst_mult_4_420  $ (!Xd_0__inst_mult_4_424  $ (Xd_0__inst_mult_4_63_sumout )) ) + ( Xd_0__inst_mult_4_290  ) + ( Xd_0__inst_mult_4_289  ))
// Xd_0__inst_mult_4_298  = SHARE((!Xd_0__inst_mult_4_420  & (Xd_0__inst_mult_4_424  & Xd_0__inst_mult_4_63_sumout )) # (Xd_0__inst_mult_4_420  & ((Xd_0__inst_mult_4_63_sumout ) # (Xd_0__inst_mult_4_424 ))))

	.dataa(!Xd_0__inst_mult_4_420 ),
	.datab(!Xd_0__inst_mult_4_424 ),
	.datac(!Xd_0__inst_mult_4_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_289 ),
	.sharein(Xd_0__inst_mult_4_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_296 ),
	.cout(Xd_0__inst_mult_4_297 ),
	.shareout(Xd_0__inst_mult_4_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_100 (
// Equation(s):
// Xd_0__inst_mult_4_300  = SUM(( !Xd_0__inst_mult_4_428  $ (((!din_a[49]) # (!din_b[55]))) ) + ( Xd_0__inst_mult_4_434  ) + ( Xd_0__inst_mult_4_433  ))
// Xd_0__inst_mult_4_301  = CARRY(( !Xd_0__inst_mult_4_428  $ (((!din_a[49]) # (!din_b[55]))) ) + ( Xd_0__inst_mult_4_434  ) + ( Xd_0__inst_mult_4_433  ))
// Xd_0__inst_mult_4_302  = SHARE((din_a[49] & (din_b[55] & Xd_0__inst_mult_4_428 )))

	.dataa(!din_a[49]),
	.datab(!din_b[55]),
	.datac(!Xd_0__inst_mult_4_428 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_433 ),
	.sharein(Xd_0__inst_mult_4_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_300 ),
	.cout(Xd_0__inst_mult_4_301 ),
	.shareout(Xd_0__inst_mult_4_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_99 (
// Equation(s):
// Xd_0__inst_mult_5_296  = SUM(( !Xd_0__inst_mult_5_416  $ (!Xd_0__inst_mult_5_420  $ (Xd_0__inst_mult_5_67_sumout )) ) + ( Xd_0__inst_mult_5_290  ) + ( Xd_0__inst_mult_5_289  ))
// Xd_0__inst_mult_5_297  = CARRY(( !Xd_0__inst_mult_5_416  $ (!Xd_0__inst_mult_5_420  $ (Xd_0__inst_mult_5_67_sumout )) ) + ( Xd_0__inst_mult_5_290  ) + ( Xd_0__inst_mult_5_289  ))
// Xd_0__inst_mult_5_298  = SHARE((!Xd_0__inst_mult_5_416  & (Xd_0__inst_mult_5_420  & Xd_0__inst_mult_5_67_sumout )) # (Xd_0__inst_mult_5_416  & ((Xd_0__inst_mult_5_67_sumout ) # (Xd_0__inst_mult_5_420 ))))

	.dataa(!Xd_0__inst_mult_5_416 ),
	.datab(!Xd_0__inst_mult_5_420 ),
	.datac(!Xd_0__inst_mult_5_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_289 ),
	.sharein(Xd_0__inst_mult_5_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_296 ),
	.cout(Xd_0__inst_mult_5_297 ),
	.shareout(Xd_0__inst_mult_5_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_100 (
// Equation(s):
// Xd_0__inst_mult_5_300  = SUM(( !Xd_0__inst_mult_5_424  $ (((!din_a[61]) # (!din_b[67]))) ) + ( Xd_0__inst_mult_5_430  ) + ( Xd_0__inst_mult_5_429  ))
// Xd_0__inst_mult_5_301  = CARRY(( !Xd_0__inst_mult_5_424  $ (((!din_a[61]) # (!din_b[67]))) ) + ( Xd_0__inst_mult_5_430  ) + ( Xd_0__inst_mult_5_429  ))
// Xd_0__inst_mult_5_302  = SHARE((din_a[61] & (din_b[67] & Xd_0__inst_mult_5_424 )))

	.dataa(!din_a[61]),
	.datab(!din_b[67]),
	.datac(!Xd_0__inst_mult_5_424 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_429 ),
	.sharein(Xd_0__inst_mult_5_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_300 ),
	.cout(Xd_0__inst_mult_5_301 ),
	.shareout(Xd_0__inst_mult_5_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_99 (
// Equation(s):
// Xd_0__inst_mult_2_296  = SUM(( !Xd_0__inst_mult_2_416  $ (!Xd_0__inst_mult_2_420  $ (Xd_0__inst_mult_2_63_sumout )) ) + ( Xd_0__inst_mult_2_290  ) + ( Xd_0__inst_mult_2_289  ))
// Xd_0__inst_mult_2_297  = CARRY(( !Xd_0__inst_mult_2_416  $ (!Xd_0__inst_mult_2_420  $ (Xd_0__inst_mult_2_63_sumout )) ) + ( Xd_0__inst_mult_2_290  ) + ( Xd_0__inst_mult_2_289  ))
// Xd_0__inst_mult_2_298  = SHARE((!Xd_0__inst_mult_2_416  & (Xd_0__inst_mult_2_420  & Xd_0__inst_mult_2_63_sumout )) # (Xd_0__inst_mult_2_416  & ((Xd_0__inst_mult_2_63_sumout ) # (Xd_0__inst_mult_2_420 ))))

	.dataa(!Xd_0__inst_mult_2_416 ),
	.datab(!Xd_0__inst_mult_2_420 ),
	.datac(!Xd_0__inst_mult_2_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_289 ),
	.sharein(Xd_0__inst_mult_2_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_296 ),
	.cout(Xd_0__inst_mult_2_297 ),
	.shareout(Xd_0__inst_mult_2_298 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_100 (
// Equation(s):
// Xd_0__inst_mult_2_300  = SUM(( !Xd_0__inst_mult_2_424  $ (((!din_a[25]) # (!din_b[31]))) ) + ( Xd_0__inst_mult_2_430  ) + ( Xd_0__inst_mult_2_429  ))
// Xd_0__inst_mult_2_301  = CARRY(( !Xd_0__inst_mult_2_424  $ (((!din_a[25]) # (!din_b[31]))) ) + ( Xd_0__inst_mult_2_430  ) + ( Xd_0__inst_mult_2_429  ))
// Xd_0__inst_mult_2_302  = SHARE((din_a[25] & (din_b[31] & Xd_0__inst_mult_2_424 )))

	.dataa(!din_a[25]),
	.datab(!din_b[31]),
	.datac(!Xd_0__inst_mult_2_424 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_429 ),
	.sharein(Xd_0__inst_mult_2_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_300 ),
	.cout(Xd_0__inst_mult_2_301 ),
	.shareout(Xd_0__inst_mult_2_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_107 (
// Equation(s):
// Xd_0__inst_mult_3_340  = SUM(( !Xd_0__inst_mult_3_456  $ (!Xd_0__inst_mult_3_460  $ (Xd_0__inst_mult_3_63_sumout )) ) + ( Xd_0__inst_mult_3_334  ) + ( Xd_0__inst_mult_3_333  ))
// Xd_0__inst_mult_3_341  = CARRY(( !Xd_0__inst_mult_3_456  $ (!Xd_0__inst_mult_3_460  $ (Xd_0__inst_mult_3_63_sumout )) ) + ( Xd_0__inst_mult_3_334  ) + ( Xd_0__inst_mult_3_333  ))
// Xd_0__inst_mult_3_342  = SHARE((!Xd_0__inst_mult_3_456  & (Xd_0__inst_mult_3_460  & Xd_0__inst_mult_3_63_sumout )) # (Xd_0__inst_mult_3_456  & ((Xd_0__inst_mult_3_63_sumout ) # (Xd_0__inst_mult_3_460 ))))

	.dataa(!Xd_0__inst_mult_3_456 ),
	.datab(!Xd_0__inst_mult_3_460 ),
	.datac(!Xd_0__inst_mult_3_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_333 ),
	.sharein(Xd_0__inst_mult_3_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_340 ),
	.cout(Xd_0__inst_mult_3_341 ),
	.shareout(Xd_0__inst_mult_3_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_108 (
// Equation(s):
// Xd_0__inst_mult_3_344  = SUM(( !Xd_0__inst_mult_3_464  $ (((!din_a[37]) # (!din_b[43]))) ) + ( Xd_0__inst_mult_3_470  ) + ( Xd_0__inst_mult_3_469  ))
// Xd_0__inst_mult_3_345  = CARRY(( !Xd_0__inst_mult_3_464  $ (((!din_a[37]) # (!din_b[43]))) ) + ( Xd_0__inst_mult_3_470  ) + ( Xd_0__inst_mult_3_469  ))
// Xd_0__inst_mult_3_346  = SHARE((din_a[37] & (din_b[43] & Xd_0__inst_mult_3_464 )))

	.dataa(!din_a[37]),
	.datab(!din_b[43]),
	.datac(!Xd_0__inst_mult_3_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_469 ),
	.sharein(Xd_0__inst_mult_3_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_344 ),
	.cout(Xd_0__inst_mult_3_345 ),
	.shareout(Xd_0__inst_mult_3_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_101 (
// Equation(s):
// Xd_0__inst_mult_0_316  = SUM(( !Xd_0__inst_mult_0_428  $ (!Xd_0__inst_mult_0_432  $ (Xd_0__inst_mult_5_384 )) ) + ( Xd_0__inst_mult_0_310  ) + ( Xd_0__inst_mult_0_309  ))
// Xd_0__inst_mult_0_317  = CARRY(( !Xd_0__inst_mult_0_428  $ (!Xd_0__inst_mult_0_432  $ (Xd_0__inst_mult_5_384 )) ) + ( Xd_0__inst_mult_0_310  ) + ( Xd_0__inst_mult_0_309  ))
// Xd_0__inst_mult_0_318  = SHARE((!Xd_0__inst_mult_0_428  & (Xd_0__inst_mult_0_432  & Xd_0__inst_mult_5_384 )) # (Xd_0__inst_mult_0_428  & ((Xd_0__inst_mult_5_384 ) # (Xd_0__inst_mult_0_432 ))))

	.dataa(!Xd_0__inst_mult_0_428 ),
	.datab(!Xd_0__inst_mult_0_432 ),
	.datac(!Xd_0__inst_mult_5_384 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_309 ),
	.sharein(Xd_0__inst_mult_0_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_316 ),
	.cout(Xd_0__inst_mult_0_317 ),
	.shareout(Xd_0__inst_mult_0_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_102 (
// Equation(s):
// Xd_0__inst_mult_0_320  = SUM(( !Xd_0__inst_mult_0_436  $ (((!din_a[1]) # (!din_b[7]))) ) + ( Xd_0__inst_mult_0_442  ) + ( Xd_0__inst_mult_0_441  ))
// Xd_0__inst_mult_0_321  = CARRY(( !Xd_0__inst_mult_0_436  $ (((!din_a[1]) # (!din_b[7]))) ) + ( Xd_0__inst_mult_0_442  ) + ( Xd_0__inst_mult_0_441  ))
// Xd_0__inst_mult_0_322  = SHARE((din_a[1] & (din_b[7] & Xd_0__inst_mult_0_436 )))

	.dataa(!din_a[1]),
	.datab(!din_b[7]),
	.datac(!Xd_0__inst_mult_0_436 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_441 ),
	.sharein(Xd_0__inst_mult_0_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_320 ),
	.cout(Xd_0__inst_mult_0_321 ),
	.shareout(Xd_0__inst_mult_0_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_97 (
// Equation(s):
// Xd_0__inst_mult_1_300  = SUM(( !Xd_0__inst_mult_1_412  $ (!Xd_0__inst_mult_1_416  $ (Xd_0__inst_mult_1_63_sumout )) ) + ( Xd_0__inst_mult_1_294  ) + ( Xd_0__inst_mult_1_293  ))
// Xd_0__inst_mult_1_301  = CARRY(( !Xd_0__inst_mult_1_412  $ (!Xd_0__inst_mult_1_416  $ (Xd_0__inst_mult_1_63_sumout )) ) + ( Xd_0__inst_mult_1_294  ) + ( Xd_0__inst_mult_1_293  ))
// Xd_0__inst_mult_1_302  = SHARE((!Xd_0__inst_mult_1_412  & (Xd_0__inst_mult_1_416  & Xd_0__inst_mult_1_63_sumout )) # (Xd_0__inst_mult_1_412  & ((Xd_0__inst_mult_1_63_sumout ) # (Xd_0__inst_mult_1_416 ))))

	.dataa(!Xd_0__inst_mult_1_412 ),
	.datab(!Xd_0__inst_mult_1_416 ),
	.datac(!Xd_0__inst_mult_1_63_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_293 ),
	.sharein(Xd_0__inst_mult_1_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_300 ),
	.cout(Xd_0__inst_mult_1_301 ),
	.shareout(Xd_0__inst_mult_1_302 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_98 (
// Equation(s):
// Xd_0__inst_mult_1_304  = SUM(( !Xd_0__inst_mult_1_420  $ (((!din_a[13]) # (!din_b[19]))) ) + ( Xd_0__inst_mult_1_426  ) + ( Xd_0__inst_mult_1_425  ))
// Xd_0__inst_mult_1_305  = CARRY(( !Xd_0__inst_mult_1_420  $ (((!din_a[13]) # (!din_b[19]))) ) + ( Xd_0__inst_mult_1_426  ) + ( Xd_0__inst_mult_1_425  ))
// Xd_0__inst_mult_1_306  = SHARE((din_a[13] & (din_b[19] & Xd_0__inst_mult_1_420 )))

	.dataa(!din_a[13]),
	.datab(!din_b[19]),
	.datac(!Xd_0__inst_mult_1_420 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_425 ),
	.sharein(Xd_0__inst_mult_1_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_304 ),
	.cout(Xd_0__inst_mult_1_305 ),
	.shareout(Xd_0__inst_mult_1_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_131 (
// Equation(s):
// Xd_0__inst_mult_6_424  = SUM(( (din_a[78] & din_b[74]) ) + ( Xd_0__inst_mult_6_418  ) + ( Xd_0__inst_mult_6_417  ))
// Xd_0__inst_mult_6_425  = CARRY(( (din_a[78] & din_b[74]) ) + ( Xd_0__inst_mult_6_418  ) + ( Xd_0__inst_mult_6_417  ))
// Xd_0__inst_mult_6_426  = SHARE((din_a[80] & din_b[73]))

	.dataa(!din_a[78]),
	.datab(!din_b[74]),
	.datac(!din_a[80]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_417 ),
	.sharein(Xd_0__inst_mult_6_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_424 ),
	.cout(Xd_0__inst_mult_6_425 ),
	.shareout(Xd_0__inst_mult_6_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_132 (
// Equation(s):
// Xd_0__inst_mult_6_428  = SUM(( (!din_a[77] & (((din_a[76] & din_b[76])))) # (din_a[77] & (!din_b[75] $ (((!din_a[76]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_422  ) + ( Xd_0__inst_mult_6_421  ))
// Xd_0__inst_mult_6_429  = CARRY(( (!din_a[77] & (((din_a[76] & din_b[76])))) # (din_a[77] & (!din_b[75] $ (((!din_a[76]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_422  ) + ( Xd_0__inst_mult_6_421  ))
// Xd_0__inst_mult_6_430  = SHARE((din_a[77] & (din_b[75] & (din_a[76] & din_b[76]))))

	.dataa(!din_a[77]),
	.datab(!din_b[75]),
	.datac(!din_a[76]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_421 ),
	.sharein(Xd_0__inst_mult_6_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_428 ),
	.cout(Xd_0__inst_mult_6_429 ),
	.shareout(Xd_0__inst_mult_6_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_59 (
// Equation(s):
// Xd_0__inst_mult_6_59_sumout  = SUM(( (din_a[80] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_60  = CARRY(( (din_a[80] & din_b[72]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_61  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_6_59_sumout ),
	.cout(Xd_0__inst_mult_6_60 ),
	.shareout(Xd_0__inst_mult_6_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_133 (
// Equation(s):
// Xd_0__inst_mult_6_432  = SUM(( (!din_a[74] & (((din_a[75] & din_b[77])))) # (din_a[74] & (!din_b[78] $ (((!din_a[75]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_310  ) + ( Xd_0__inst_mult_6_309  ))
// Xd_0__inst_mult_6_433  = CARRY(( (!din_a[74] & (((din_a[75] & din_b[77])))) # (din_a[74] & (!din_b[78] $ (((!din_a[75]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_310  ) + ( Xd_0__inst_mult_6_309  ))
// Xd_0__inst_mult_6_434  = SHARE((din_a[74] & (din_b[78] & (din_a[75] & din_b[77]))))

	.dataa(!din_a[74]),
	.datab(!din_b[78]),
	.datac(!din_a[75]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_309 ),
	.sharein(Xd_0__inst_mult_6_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_432 ),
	.cout(Xd_0__inst_mult_6_433 ),
	.shareout(Xd_0__inst_mult_6_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_134 (
// Equation(s):
// Xd_0__inst_mult_6_437  = CARRY(( GND ) + ( Xd_0__inst_mult_4_41  ) + ( Xd_0__inst_mult_4_40  ))
// Xd_0__inst_mult_6_438  = SHARE((din_a[72] & din_b[80]))

	.dataa(!din_a[72]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_40 ),
	.sharein(Xd_0__inst_mult_4_41 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_437 ),
	.shareout(Xd_0__inst_mult_6_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_133 (
// Equation(s):
// Xd_0__inst_mult_7_432  = SUM(( (din_a[90] & din_b[86]) ) + ( Xd_0__inst_mult_7_426  ) + ( Xd_0__inst_mult_7_425  ))
// Xd_0__inst_mult_7_433  = CARRY(( (din_a[90] & din_b[86]) ) + ( Xd_0__inst_mult_7_426  ) + ( Xd_0__inst_mult_7_425  ))
// Xd_0__inst_mult_7_434  = SHARE((din_a[92] & din_b[85]))

	.dataa(!din_a[90]),
	.datab(!din_b[86]),
	.datac(!din_a[92]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_425 ),
	.sharein(Xd_0__inst_mult_7_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_432 ),
	.cout(Xd_0__inst_mult_7_433 ),
	.shareout(Xd_0__inst_mult_7_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_134 (
// Equation(s):
// Xd_0__inst_mult_7_436  = SUM(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_430  ) + ( Xd_0__inst_mult_7_429  ))
// Xd_0__inst_mult_7_437  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[88])))) # (din_a[89] & (!din_b[87] $ (((!din_a[88]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_430  ) + ( Xd_0__inst_mult_7_429  ))
// Xd_0__inst_mult_7_438  = SHARE((din_a[89] & (din_b[87] & (din_a[88] & din_b[88]))))

	.dataa(!din_a[89]),
	.datab(!din_b[87]),
	.datac(!din_a[88]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_429 ),
	.sharein(Xd_0__inst_mult_7_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_436 ),
	.cout(Xd_0__inst_mult_7_437 ),
	.shareout(Xd_0__inst_mult_7_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_59 (
// Equation(s):
// Xd_0__inst_mult_7_59_sumout  = SUM(( (din_a[92] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_60  = CARRY(( (din_a[92] & din_b[84]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_61  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_7_59_sumout ),
	.cout(Xd_0__inst_mult_7_60 ),
	.shareout(Xd_0__inst_mult_7_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_135 (
// Equation(s):
// Xd_0__inst_mult_7_440  = SUM(( (!din_a[86] & (((din_a[87] & din_b[89])))) # (din_a[86] & (!din_b[90] $ (((!din_a[87]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_318  ) + ( Xd_0__inst_mult_7_317  ))
// Xd_0__inst_mult_7_441  = CARRY(( (!din_a[86] & (((din_a[87] & din_b[89])))) # (din_a[86] & (!din_b[90] $ (((!din_a[87]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_318  ) + ( Xd_0__inst_mult_7_317  ))
// Xd_0__inst_mult_7_442  = SHARE((din_a[86] & (din_b[90] & (din_a[87] & din_b[89]))))

	.dataa(!din_a[86]),
	.datab(!din_b[90]),
	.datac(!din_a[87]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_317 ),
	.sharein(Xd_0__inst_mult_7_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_440 ),
	.cout(Xd_0__inst_mult_7_441 ),
	.shareout(Xd_0__inst_mult_7_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_136 (
// Equation(s):
// Xd_0__inst_mult_7_445  = CARRY(( GND ) + ( Xd_0__inst_mult_6_53  ) + ( Xd_0__inst_mult_6_52  ))
// Xd_0__inst_mult_7_446  = SHARE((din_a[84] & din_b[92]))

	.dataa(!din_a[84]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_52 ),
	.sharein(Xd_0__inst_mult_6_53 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_445 ),
	.shareout(Xd_0__inst_mult_7_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_101 (
// Equation(s):
// Xd_0__inst_mult_4_304  = SUM(( !Xd_0__inst_mult_4_436  $ (!Xd_0__inst_mult_4_440  $ (Xd_0__inst_mult_4_67_sumout )) ) + ( Xd_0__inst_mult_4_298  ) + ( Xd_0__inst_mult_4_297  ))
// Xd_0__inst_mult_4_305  = CARRY(( !Xd_0__inst_mult_4_436  $ (!Xd_0__inst_mult_4_440  $ (Xd_0__inst_mult_4_67_sumout )) ) + ( Xd_0__inst_mult_4_298  ) + ( Xd_0__inst_mult_4_297  ))
// Xd_0__inst_mult_4_306  = SHARE((!Xd_0__inst_mult_4_436  & (Xd_0__inst_mult_4_440  & Xd_0__inst_mult_4_67_sumout )) # (Xd_0__inst_mult_4_436  & ((Xd_0__inst_mult_4_67_sumout ) # (Xd_0__inst_mult_4_440 ))))

	.dataa(!Xd_0__inst_mult_4_436 ),
	.datab(!Xd_0__inst_mult_4_440 ),
	.datac(!Xd_0__inst_mult_4_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_297 ),
	.sharein(Xd_0__inst_mult_4_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_304 ),
	.cout(Xd_0__inst_mult_4_305 ),
	.shareout(Xd_0__inst_mult_4_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_102 (
// Equation(s):
// Xd_0__inst_mult_4_308  = SUM(( !Xd_0__inst_mult_4_444  $ (!Xd_0__inst_mult_4_448 ) ) + ( Xd_0__inst_mult_4_302  ) + ( Xd_0__inst_mult_4_301  ))
// Xd_0__inst_mult_4_309  = CARRY(( !Xd_0__inst_mult_4_444  $ (!Xd_0__inst_mult_4_448 ) ) + ( Xd_0__inst_mult_4_302  ) + ( Xd_0__inst_mult_4_301  ))
// Xd_0__inst_mult_4_310  = SHARE((Xd_0__inst_mult_4_444  & Xd_0__inst_mult_4_448 ))

	.dataa(!Xd_0__inst_mult_4_444 ),
	.datab(!Xd_0__inst_mult_4_448 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_301 ),
	.sharein(Xd_0__inst_mult_4_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_308 ),
	.cout(Xd_0__inst_mult_4_309 ),
	.shareout(Xd_0__inst_mult_4_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_101 (
// Equation(s):
// Xd_0__inst_mult_5_304  = SUM(( !Xd_0__inst_mult_5_432  $ (!Xd_0__inst_mult_5_436  $ (Xd_0__inst_mult_5_35_sumout )) ) + ( Xd_0__inst_mult_5_298  ) + ( Xd_0__inst_mult_5_297  ))
// Xd_0__inst_mult_5_305  = CARRY(( !Xd_0__inst_mult_5_432  $ (!Xd_0__inst_mult_5_436  $ (Xd_0__inst_mult_5_35_sumout )) ) + ( Xd_0__inst_mult_5_298  ) + ( Xd_0__inst_mult_5_297  ))
// Xd_0__inst_mult_5_306  = SHARE((!Xd_0__inst_mult_5_432  & (Xd_0__inst_mult_5_436  & Xd_0__inst_mult_5_35_sumout )) # (Xd_0__inst_mult_5_432  & ((Xd_0__inst_mult_5_35_sumout ) # (Xd_0__inst_mult_5_436 ))))

	.dataa(!Xd_0__inst_mult_5_432 ),
	.datab(!Xd_0__inst_mult_5_436 ),
	.datac(!Xd_0__inst_mult_5_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_297 ),
	.sharein(Xd_0__inst_mult_5_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_304 ),
	.cout(Xd_0__inst_mult_5_305 ),
	.shareout(Xd_0__inst_mult_5_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_102 (
// Equation(s):
// Xd_0__inst_mult_5_308  = SUM(( !Xd_0__inst_mult_5_440  $ (!Xd_0__inst_mult_5_444 ) ) + ( Xd_0__inst_mult_5_302  ) + ( Xd_0__inst_mult_5_301  ))
// Xd_0__inst_mult_5_309  = CARRY(( !Xd_0__inst_mult_5_440  $ (!Xd_0__inst_mult_5_444 ) ) + ( Xd_0__inst_mult_5_302  ) + ( Xd_0__inst_mult_5_301  ))
// Xd_0__inst_mult_5_310  = SHARE((Xd_0__inst_mult_5_440  & Xd_0__inst_mult_5_444 ))

	.dataa(!Xd_0__inst_mult_5_440 ),
	.datab(!Xd_0__inst_mult_5_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_301 ),
	.sharein(Xd_0__inst_mult_5_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_308 ),
	.cout(Xd_0__inst_mult_5_309 ),
	.shareout(Xd_0__inst_mult_5_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_101 (
// Equation(s):
// Xd_0__inst_mult_2_304  = SUM(( !Xd_0__inst_mult_2_432  $ (!Xd_0__inst_mult_2_436  $ (Xd_0__inst_mult_2_67_sumout )) ) + ( Xd_0__inst_mult_2_298  ) + ( Xd_0__inst_mult_2_297  ))
// Xd_0__inst_mult_2_305  = CARRY(( !Xd_0__inst_mult_2_432  $ (!Xd_0__inst_mult_2_436  $ (Xd_0__inst_mult_2_67_sumout )) ) + ( Xd_0__inst_mult_2_298  ) + ( Xd_0__inst_mult_2_297  ))
// Xd_0__inst_mult_2_306  = SHARE((!Xd_0__inst_mult_2_432  & (Xd_0__inst_mult_2_436  & Xd_0__inst_mult_2_67_sumout )) # (Xd_0__inst_mult_2_432  & ((Xd_0__inst_mult_2_67_sumout ) # (Xd_0__inst_mult_2_436 ))))

	.dataa(!Xd_0__inst_mult_2_432 ),
	.datab(!Xd_0__inst_mult_2_436 ),
	.datac(!Xd_0__inst_mult_2_67_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_297 ),
	.sharein(Xd_0__inst_mult_2_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_304 ),
	.cout(Xd_0__inst_mult_2_305 ),
	.shareout(Xd_0__inst_mult_2_306 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_102 (
// Equation(s):
// Xd_0__inst_mult_2_308  = SUM(( !Xd_0__inst_mult_2_440  $ (!Xd_0__inst_mult_2_444 ) ) + ( Xd_0__inst_mult_2_302  ) + ( Xd_0__inst_mult_2_301  ))
// Xd_0__inst_mult_2_309  = CARRY(( !Xd_0__inst_mult_2_440  $ (!Xd_0__inst_mult_2_444 ) ) + ( Xd_0__inst_mult_2_302  ) + ( Xd_0__inst_mult_2_301  ))
// Xd_0__inst_mult_2_310  = SHARE((Xd_0__inst_mult_2_440  & Xd_0__inst_mult_2_444 ))

	.dataa(!Xd_0__inst_mult_2_440 ),
	.datab(!Xd_0__inst_mult_2_444 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_301 ),
	.sharein(Xd_0__inst_mult_2_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_308 ),
	.cout(Xd_0__inst_mult_2_309 ),
	.shareout(Xd_0__inst_mult_2_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_109 (
// Equation(s):
// Xd_0__inst_mult_3_348  = SUM(( !Xd_0__inst_mult_3_472  $ (!Xd_0__inst_mult_3_476  $ (Xd_0__inst_mult_4_388 )) ) + ( Xd_0__inst_mult_3_342  ) + ( Xd_0__inst_mult_3_341  ))
// Xd_0__inst_mult_3_349  = CARRY(( !Xd_0__inst_mult_3_472  $ (!Xd_0__inst_mult_3_476  $ (Xd_0__inst_mult_4_388 )) ) + ( Xd_0__inst_mult_3_342  ) + ( Xd_0__inst_mult_3_341  ))
// Xd_0__inst_mult_3_350  = SHARE((!Xd_0__inst_mult_3_472  & (Xd_0__inst_mult_3_476  & Xd_0__inst_mult_4_388 )) # (Xd_0__inst_mult_3_472  & ((Xd_0__inst_mult_4_388 ) # (Xd_0__inst_mult_3_476 ))))

	.dataa(!Xd_0__inst_mult_3_472 ),
	.datab(!Xd_0__inst_mult_3_476 ),
	.datac(!Xd_0__inst_mult_4_388 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_341 ),
	.sharein(Xd_0__inst_mult_3_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_348 ),
	.cout(Xd_0__inst_mult_3_349 ),
	.shareout(Xd_0__inst_mult_3_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_110 (
// Equation(s):
// Xd_0__inst_mult_3_352  = SUM(( !Xd_0__inst_mult_3_480  $ (!Xd_0__inst_mult_3_484 ) ) + ( Xd_0__inst_mult_3_346  ) + ( Xd_0__inst_mult_3_345  ))
// Xd_0__inst_mult_3_353  = CARRY(( !Xd_0__inst_mult_3_480  $ (!Xd_0__inst_mult_3_484 ) ) + ( Xd_0__inst_mult_3_346  ) + ( Xd_0__inst_mult_3_345  ))
// Xd_0__inst_mult_3_354  = SHARE((Xd_0__inst_mult_3_480  & Xd_0__inst_mult_3_484 ))

	.dataa(!Xd_0__inst_mult_3_480 ),
	.datab(!Xd_0__inst_mult_3_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_345 ),
	.sharein(Xd_0__inst_mult_3_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_352 ),
	.cout(Xd_0__inst_mult_3_353 ),
	.shareout(Xd_0__inst_mult_3_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_103 (
// Equation(s):
// Xd_0__inst_mult_0_324  = SUM(( !Xd_0__inst_mult_0_444  $ (!Xd_0__inst_mult_0_448  $ (Xd_0__inst_mult_0_47_sumout )) ) + ( Xd_0__inst_mult_0_318  ) + ( Xd_0__inst_mult_0_317  ))
// Xd_0__inst_mult_0_325  = CARRY(( !Xd_0__inst_mult_0_444  $ (!Xd_0__inst_mult_0_448  $ (Xd_0__inst_mult_0_47_sumout )) ) + ( Xd_0__inst_mult_0_318  ) + ( Xd_0__inst_mult_0_317  ))
// Xd_0__inst_mult_0_326  = SHARE((!Xd_0__inst_mult_0_444  & (Xd_0__inst_mult_0_448  & Xd_0__inst_mult_0_47_sumout )) # (Xd_0__inst_mult_0_444  & ((Xd_0__inst_mult_0_47_sumout ) # (Xd_0__inst_mult_0_448 ))))

	.dataa(!Xd_0__inst_mult_0_444 ),
	.datab(!Xd_0__inst_mult_0_448 ),
	.datac(!Xd_0__inst_mult_0_47_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_317 ),
	.sharein(Xd_0__inst_mult_0_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_324 ),
	.cout(Xd_0__inst_mult_0_325 ),
	.shareout(Xd_0__inst_mult_0_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_104 (
// Equation(s):
// Xd_0__inst_mult_0_328  = SUM(( !Xd_0__inst_mult_0_452  $ (!Xd_0__inst_mult_0_456 ) ) + ( Xd_0__inst_mult_0_322  ) + ( Xd_0__inst_mult_0_321  ))
// Xd_0__inst_mult_0_329  = CARRY(( !Xd_0__inst_mult_0_452  $ (!Xd_0__inst_mult_0_456 ) ) + ( Xd_0__inst_mult_0_322  ) + ( Xd_0__inst_mult_0_321  ))
// Xd_0__inst_mult_0_330  = SHARE((Xd_0__inst_mult_0_452  & Xd_0__inst_mult_0_456 ))

	.dataa(!Xd_0__inst_mult_0_452 ),
	.datab(!Xd_0__inst_mult_0_456 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_321 ),
	.sharein(Xd_0__inst_mult_0_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_328 ),
	.cout(Xd_0__inst_mult_0_329 ),
	.shareout(Xd_0__inst_mult_0_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_99 (
// Equation(s):
// Xd_0__inst_mult_1_308  = SUM(( !Xd_0__inst_mult_1_428  $ (!Xd_0__inst_mult_1_432  $ (Xd_0__inst_mult_1_43_sumout )) ) + ( Xd_0__inst_mult_1_302  ) + ( Xd_0__inst_mult_1_301  ))
// Xd_0__inst_mult_1_309  = CARRY(( !Xd_0__inst_mult_1_428  $ (!Xd_0__inst_mult_1_432  $ (Xd_0__inst_mult_1_43_sumout )) ) + ( Xd_0__inst_mult_1_302  ) + ( Xd_0__inst_mult_1_301  ))
// Xd_0__inst_mult_1_310  = SHARE((!Xd_0__inst_mult_1_428  & (Xd_0__inst_mult_1_432  & Xd_0__inst_mult_1_43_sumout )) # (Xd_0__inst_mult_1_428  & ((Xd_0__inst_mult_1_43_sumout ) # (Xd_0__inst_mult_1_432 ))))

	.dataa(!Xd_0__inst_mult_1_428 ),
	.datab(!Xd_0__inst_mult_1_432 ),
	.datac(!Xd_0__inst_mult_1_43_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_301 ),
	.sharein(Xd_0__inst_mult_1_302 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_308 ),
	.cout(Xd_0__inst_mult_1_309 ),
	.shareout(Xd_0__inst_mult_1_310 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_100 (
// Equation(s):
// Xd_0__inst_mult_1_312  = SUM(( !Xd_0__inst_mult_1_436  $ (!Xd_0__inst_mult_1_440 ) ) + ( Xd_0__inst_mult_1_306  ) + ( Xd_0__inst_mult_1_305  ))
// Xd_0__inst_mult_1_313  = CARRY(( !Xd_0__inst_mult_1_436  $ (!Xd_0__inst_mult_1_440 ) ) + ( Xd_0__inst_mult_1_306  ) + ( Xd_0__inst_mult_1_305  ))
// Xd_0__inst_mult_1_314  = SHARE((Xd_0__inst_mult_1_436  & Xd_0__inst_mult_1_440 ))

	.dataa(!Xd_0__inst_mult_1_436 ),
	.datab(!Xd_0__inst_mult_1_440 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_305 ),
	.sharein(Xd_0__inst_mult_1_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_312 ),
	.cout(Xd_0__inst_mult_1_313 ),
	.shareout(Xd_0__inst_mult_1_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_135 (
// Equation(s):
// Xd_0__inst_mult_6_440  = SUM(( (din_a[79] & din_b[74]) ) + ( Xd_0__inst_mult_6_426  ) + ( Xd_0__inst_mult_6_425  ))
// Xd_0__inst_mult_6_441  = CARRY(( (din_a[79] & din_b[74]) ) + ( Xd_0__inst_mult_6_426  ) + ( Xd_0__inst_mult_6_425  ))
// Xd_0__inst_mult_6_442  = SHARE((din_a[81] & din_b[73]))

	.dataa(!din_a[79]),
	.datab(!din_b[74]),
	.datac(!din_a[81]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_425 ),
	.sharein(Xd_0__inst_mult_6_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_440 ),
	.cout(Xd_0__inst_mult_6_441 ),
	.shareout(Xd_0__inst_mult_6_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_136 (
// Equation(s):
// Xd_0__inst_mult_6_444  = SUM(( (!din_a[78] & (((din_a[77] & din_b[76])))) # (din_a[78] & (!din_b[75] $ (((!din_a[77]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_430  ) + ( Xd_0__inst_mult_6_429  ))
// Xd_0__inst_mult_6_445  = CARRY(( (!din_a[78] & (((din_a[77] & din_b[76])))) # (din_a[78] & (!din_b[75] $ (((!din_a[77]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_430  ) + ( Xd_0__inst_mult_6_429  ))
// Xd_0__inst_mult_6_446  = SHARE((din_a[78] & (din_b[75] & (din_a[77] & din_b[76]))))

	.dataa(!din_a[78]),
	.datab(!din_b[75]),
	.datac(!din_a[77]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_429 ),
	.sharein(Xd_0__inst_mult_6_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_444 ),
	.cout(Xd_0__inst_mult_6_445 ),
	.shareout(Xd_0__inst_mult_6_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_63 (
// Equation(s):
// Xd_0__inst_mult_6_63_sumout  = SUM(( (din_a[81] & din_b[72]) ) + ( Xd_0__inst_mult_7_61  ) + ( Xd_0__inst_mult_7_60  ))
// Xd_0__inst_mult_6_64  = CARRY(( (din_a[81] & din_b[72]) ) + ( Xd_0__inst_mult_7_61  ) + ( Xd_0__inst_mult_7_60  ))
// Xd_0__inst_mult_6_65  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_60 ),
	.sharein(Xd_0__inst_mult_7_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_63_sumout ),
	.cout(Xd_0__inst_mult_6_64 ),
	.shareout(Xd_0__inst_mult_6_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_137 (
// Equation(s):
// Xd_0__inst_mult_6_448  = SUM(( (!din_a[75] & (((din_a[76] & din_b[77])))) # (din_a[75] & (!din_b[78] $ (((!din_a[76]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_434  ) + ( Xd_0__inst_mult_6_433  ))
// Xd_0__inst_mult_6_449  = CARRY(( (!din_a[75] & (((din_a[76] & din_b[77])))) # (din_a[75] & (!din_b[78] $ (((!din_a[76]) # (!din_b[77]))))) ) + ( Xd_0__inst_mult_6_434  ) + ( Xd_0__inst_mult_6_433  ))
// Xd_0__inst_mult_6_450  = SHARE((din_a[75] & (din_b[78] & (din_a[76] & din_b[77]))))

	.dataa(!din_a[75]),
	.datab(!din_b[78]),
	.datac(!din_a[76]),
	.datad(!din_b[77]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_433 ),
	.sharein(Xd_0__inst_mult_6_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_448 ),
	.cout(Xd_0__inst_mult_6_449 ),
	.shareout(Xd_0__inst_mult_6_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_138 (
// Equation(s):
// Xd_0__inst_mult_6_452  = SUM(( (din_a[72] & din_b[81]) ) + ( Xd_0__inst_mult_6_578  ) + ( Xd_0__inst_mult_6_577  ))
// Xd_0__inst_mult_6_453  = CARRY(( (din_a[72] & din_b[81]) ) + ( Xd_0__inst_mult_6_578  ) + ( Xd_0__inst_mult_6_577  ))
// Xd_0__inst_mult_6_454  = SHARE((din_a[72] & din_b[82]))

	.dataa(!din_a[72]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_577 ),
	.sharein(Xd_0__inst_mult_6_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_452 ),
	.cout(Xd_0__inst_mult_6_453 ),
	.shareout(Xd_0__inst_mult_6_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_137 (
// Equation(s):
// Xd_0__inst_mult_7_448  = SUM(( (din_a[91] & din_b[86]) ) + ( Xd_0__inst_mult_7_434  ) + ( Xd_0__inst_mult_7_433  ))
// Xd_0__inst_mult_7_449  = CARRY(( (din_a[91] & din_b[86]) ) + ( Xd_0__inst_mult_7_434  ) + ( Xd_0__inst_mult_7_433  ))
// Xd_0__inst_mult_7_450  = SHARE((din_a[93] & din_b[85]))

	.dataa(!din_a[91]),
	.datab(!din_b[86]),
	.datac(!din_a[93]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_433 ),
	.sharein(Xd_0__inst_mult_7_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_448 ),
	.cout(Xd_0__inst_mult_7_449 ),
	.shareout(Xd_0__inst_mult_7_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_138 (
// Equation(s):
// Xd_0__inst_mult_7_452  = SUM(( (!din_a[90] & (((din_a[89] & din_b[88])))) # (din_a[90] & (!din_b[87] $ (((!din_a[89]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_438  ) + ( Xd_0__inst_mult_7_437  ))
// Xd_0__inst_mult_7_453  = CARRY(( (!din_a[90] & (((din_a[89] & din_b[88])))) # (din_a[90] & (!din_b[87] $ (((!din_a[89]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_438  ) + ( Xd_0__inst_mult_7_437  ))
// Xd_0__inst_mult_7_454  = SHARE((din_a[90] & (din_b[87] & (din_a[89] & din_b[88]))))

	.dataa(!din_a[90]),
	.datab(!din_b[87]),
	.datac(!din_a[89]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_437 ),
	.sharein(Xd_0__inst_mult_7_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_452 ),
	.cout(Xd_0__inst_mult_7_453 ),
	.shareout(Xd_0__inst_mult_7_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_63 (
// Equation(s):
// Xd_0__inst_mult_7_63_sumout  = SUM(( (din_a[93] & din_b[84]) ) + ( Xd_0__inst_mult_6_65  ) + ( Xd_0__inst_mult_6_64  ))
// Xd_0__inst_mult_7_64  = CARRY(( (din_a[93] & din_b[84]) ) + ( Xd_0__inst_mult_6_65  ) + ( Xd_0__inst_mult_6_64  ))
// Xd_0__inst_mult_7_65  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_64 ),
	.sharein(Xd_0__inst_mult_6_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_63_sumout ),
	.cout(Xd_0__inst_mult_7_64 ),
	.shareout(Xd_0__inst_mult_7_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_139 (
// Equation(s):
// Xd_0__inst_mult_7_456  = SUM(( (!din_a[87] & (((din_a[88] & din_b[89])))) # (din_a[87] & (!din_b[90] $ (((!din_a[88]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_442  ) + ( Xd_0__inst_mult_7_441  ))
// Xd_0__inst_mult_7_457  = CARRY(( (!din_a[87] & (((din_a[88] & din_b[89])))) # (din_a[87] & (!din_b[90] $ (((!din_a[88]) # (!din_b[89]))))) ) + ( Xd_0__inst_mult_7_442  ) + ( Xd_0__inst_mult_7_441  ))
// Xd_0__inst_mult_7_458  = SHARE((din_a[87] & (din_b[90] & (din_a[88] & din_b[89]))))

	.dataa(!din_a[87]),
	.datab(!din_b[90]),
	.datac(!din_a[88]),
	.datad(!din_b[89]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_441 ),
	.sharein(Xd_0__inst_mult_7_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_456 ),
	.cout(Xd_0__inst_mult_7_457 ),
	.shareout(Xd_0__inst_mult_7_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_140 (
// Equation(s):
// Xd_0__inst_mult_7_460  = SUM(( (din_a[84] & din_b[93]) ) + ( Xd_0__inst_mult_7_578  ) + ( Xd_0__inst_mult_7_577  ))
// Xd_0__inst_mult_7_461  = CARRY(( (din_a[84] & din_b[93]) ) + ( Xd_0__inst_mult_7_578  ) + ( Xd_0__inst_mult_7_577  ))
// Xd_0__inst_mult_7_462  = SHARE((din_a[84] & din_b[94]))

	.dataa(!din_a[84]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_577 ),
	.sharein(Xd_0__inst_mult_7_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_460 ),
	.cout(Xd_0__inst_mult_7_461 ),
	.shareout(Xd_0__inst_mult_7_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_103 (
// Equation(s):
// Xd_0__inst_mult_4_312  = SUM(( !Xd_0__inst_mult_4_452  $ (!Xd_0__inst_mult_4_456  $ (Xd_0__inst_mult_4_35_sumout )) ) + ( Xd_0__inst_mult_4_306  ) + ( Xd_0__inst_mult_4_305  ))
// Xd_0__inst_mult_4_313  = CARRY(( !Xd_0__inst_mult_4_452  $ (!Xd_0__inst_mult_4_456  $ (Xd_0__inst_mult_4_35_sumout )) ) + ( Xd_0__inst_mult_4_306  ) + ( Xd_0__inst_mult_4_305  ))
// Xd_0__inst_mult_4_314  = SHARE((!Xd_0__inst_mult_4_452  & (Xd_0__inst_mult_4_456  & Xd_0__inst_mult_4_35_sumout )) # (Xd_0__inst_mult_4_452  & ((Xd_0__inst_mult_4_35_sumout ) # (Xd_0__inst_mult_4_456 ))))

	.dataa(!Xd_0__inst_mult_4_452 ),
	.datab(!Xd_0__inst_mult_4_456 ),
	.datac(!Xd_0__inst_mult_4_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_305 ),
	.sharein(Xd_0__inst_mult_4_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_312 ),
	.cout(Xd_0__inst_mult_4_313 ),
	.shareout(Xd_0__inst_mult_4_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_104 (
// Equation(s):
// Xd_0__inst_mult_4_316  = SUM(( !Xd_0__inst_mult_4_460  $ (!Xd_0__inst_mult_4_464  $ (Xd_0__inst_mult_4_468 )) ) + ( Xd_0__inst_mult_4_310  ) + ( Xd_0__inst_mult_4_309  ))
// Xd_0__inst_mult_4_317  = CARRY(( !Xd_0__inst_mult_4_460  $ (!Xd_0__inst_mult_4_464  $ (Xd_0__inst_mult_4_468 )) ) + ( Xd_0__inst_mult_4_310  ) + ( Xd_0__inst_mult_4_309  ))
// Xd_0__inst_mult_4_318  = SHARE((!Xd_0__inst_mult_4_460  & (Xd_0__inst_mult_4_464  & Xd_0__inst_mult_4_468 )) # (Xd_0__inst_mult_4_460  & ((Xd_0__inst_mult_4_468 ) # (Xd_0__inst_mult_4_464 ))))

	.dataa(!Xd_0__inst_mult_4_460 ),
	.datab(!Xd_0__inst_mult_4_464 ),
	.datac(!Xd_0__inst_mult_4_468 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_309 ),
	.sharein(Xd_0__inst_mult_4_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_316 ),
	.cout(Xd_0__inst_mult_4_317 ),
	.shareout(Xd_0__inst_mult_4_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_103 (
// Equation(s):
// Xd_0__inst_mult_5_312  = SUM(( !Xd_0__inst_mult_5_448  $ (!Xd_0__inst_mult_5_452  $ (Xd_0__inst_mult_5_47_sumout )) ) + ( Xd_0__inst_mult_5_306  ) + ( Xd_0__inst_mult_5_305  ))
// Xd_0__inst_mult_5_313  = CARRY(( !Xd_0__inst_mult_5_448  $ (!Xd_0__inst_mult_5_452  $ (Xd_0__inst_mult_5_47_sumout )) ) + ( Xd_0__inst_mult_5_306  ) + ( Xd_0__inst_mult_5_305  ))
// Xd_0__inst_mult_5_314  = SHARE((!Xd_0__inst_mult_5_448  & (Xd_0__inst_mult_5_452  & Xd_0__inst_mult_5_47_sumout )) # (Xd_0__inst_mult_5_448  & ((Xd_0__inst_mult_5_47_sumout ) # (Xd_0__inst_mult_5_452 ))))

	.dataa(!Xd_0__inst_mult_5_448 ),
	.datab(!Xd_0__inst_mult_5_452 ),
	.datac(!Xd_0__inst_mult_5_47_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_305 ),
	.sharein(Xd_0__inst_mult_5_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_312 ),
	.cout(Xd_0__inst_mult_5_313 ),
	.shareout(Xd_0__inst_mult_5_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_104 (
// Equation(s):
// Xd_0__inst_mult_5_316  = SUM(( !Xd_0__inst_mult_5_456  $ (!Xd_0__inst_mult_5_460  $ (Xd_0__inst_mult_5_464 )) ) + ( Xd_0__inst_mult_5_310  ) + ( Xd_0__inst_mult_5_309  ))
// Xd_0__inst_mult_5_317  = CARRY(( !Xd_0__inst_mult_5_456  $ (!Xd_0__inst_mult_5_460  $ (Xd_0__inst_mult_5_464 )) ) + ( Xd_0__inst_mult_5_310  ) + ( Xd_0__inst_mult_5_309  ))
// Xd_0__inst_mult_5_318  = SHARE((!Xd_0__inst_mult_5_456  & (Xd_0__inst_mult_5_460  & Xd_0__inst_mult_5_464 )) # (Xd_0__inst_mult_5_456  & ((Xd_0__inst_mult_5_464 ) # (Xd_0__inst_mult_5_460 ))))

	.dataa(!Xd_0__inst_mult_5_456 ),
	.datab(!Xd_0__inst_mult_5_460 ),
	.datac(!Xd_0__inst_mult_5_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_309 ),
	.sharein(Xd_0__inst_mult_5_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_316 ),
	.cout(Xd_0__inst_mult_5_317 ),
	.shareout(Xd_0__inst_mult_5_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_103 (
// Equation(s):
// Xd_0__inst_mult_2_312  = SUM(( !Xd_0__inst_mult_2_448  $ (!Xd_0__inst_mult_2_452  $ (Xd_0__inst_mult_2_47_sumout )) ) + ( Xd_0__inst_mult_2_306  ) + ( Xd_0__inst_mult_2_305  ))
// Xd_0__inst_mult_2_313  = CARRY(( !Xd_0__inst_mult_2_448  $ (!Xd_0__inst_mult_2_452  $ (Xd_0__inst_mult_2_47_sumout )) ) + ( Xd_0__inst_mult_2_306  ) + ( Xd_0__inst_mult_2_305  ))
// Xd_0__inst_mult_2_314  = SHARE((!Xd_0__inst_mult_2_448  & (Xd_0__inst_mult_2_452  & Xd_0__inst_mult_2_47_sumout )) # (Xd_0__inst_mult_2_448  & ((Xd_0__inst_mult_2_47_sumout ) # (Xd_0__inst_mult_2_452 ))))

	.dataa(!Xd_0__inst_mult_2_448 ),
	.datab(!Xd_0__inst_mult_2_452 ),
	.datac(!Xd_0__inst_mult_2_47_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_305 ),
	.sharein(Xd_0__inst_mult_2_306 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_312 ),
	.cout(Xd_0__inst_mult_2_313 ),
	.shareout(Xd_0__inst_mult_2_314 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_104 (
// Equation(s):
// Xd_0__inst_mult_2_316  = SUM(( !Xd_0__inst_mult_2_456  $ (!Xd_0__inst_mult_2_460  $ (Xd_0__inst_mult_2_464 )) ) + ( Xd_0__inst_mult_2_310  ) + ( Xd_0__inst_mult_2_309  ))
// Xd_0__inst_mult_2_317  = CARRY(( !Xd_0__inst_mult_2_456  $ (!Xd_0__inst_mult_2_460  $ (Xd_0__inst_mult_2_464 )) ) + ( Xd_0__inst_mult_2_310  ) + ( Xd_0__inst_mult_2_309  ))
// Xd_0__inst_mult_2_318  = SHARE((!Xd_0__inst_mult_2_456  & (Xd_0__inst_mult_2_460  & Xd_0__inst_mult_2_464 )) # (Xd_0__inst_mult_2_456  & ((Xd_0__inst_mult_2_464 ) # (Xd_0__inst_mult_2_460 ))))

	.dataa(!Xd_0__inst_mult_2_456 ),
	.datab(!Xd_0__inst_mult_2_460 ),
	.datac(!Xd_0__inst_mult_2_464 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_309 ),
	.sharein(Xd_0__inst_mult_2_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_316 ),
	.cout(Xd_0__inst_mult_2_317 ),
	.shareout(Xd_0__inst_mult_2_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_111 (
// Equation(s):
// Xd_0__inst_mult_3_356  = SUM(( !Xd_0__inst_mult_3_488  $ (!Xd_0__inst_mult_3_492  $ (Xd_0__inst_mult_3_35_sumout )) ) + ( Xd_0__inst_mult_3_350  ) + ( Xd_0__inst_mult_3_349  ))
// Xd_0__inst_mult_3_357  = CARRY(( !Xd_0__inst_mult_3_488  $ (!Xd_0__inst_mult_3_492  $ (Xd_0__inst_mult_3_35_sumout )) ) + ( Xd_0__inst_mult_3_350  ) + ( Xd_0__inst_mult_3_349  ))
// Xd_0__inst_mult_3_358  = SHARE((!Xd_0__inst_mult_3_488  & (Xd_0__inst_mult_3_492  & Xd_0__inst_mult_3_35_sumout )) # (Xd_0__inst_mult_3_488  & ((Xd_0__inst_mult_3_35_sumout ) # (Xd_0__inst_mult_3_492 ))))

	.dataa(!Xd_0__inst_mult_3_488 ),
	.datab(!Xd_0__inst_mult_3_492 ),
	.datac(!Xd_0__inst_mult_3_35_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_349 ),
	.sharein(Xd_0__inst_mult_3_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_356 ),
	.cout(Xd_0__inst_mult_3_357 ),
	.shareout(Xd_0__inst_mult_3_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_112 (
// Equation(s):
// Xd_0__inst_mult_3_360  = SUM(( !Xd_0__inst_mult_3_496  $ (!Xd_0__inst_mult_3_500  $ (Xd_0__inst_mult_3_504 )) ) + ( Xd_0__inst_mult_3_354  ) + ( Xd_0__inst_mult_3_353  ))
// Xd_0__inst_mult_3_361  = CARRY(( !Xd_0__inst_mult_3_496  $ (!Xd_0__inst_mult_3_500  $ (Xd_0__inst_mult_3_504 )) ) + ( Xd_0__inst_mult_3_354  ) + ( Xd_0__inst_mult_3_353  ))
// Xd_0__inst_mult_3_362  = SHARE((!Xd_0__inst_mult_3_496  & (Xd_0__inst_mult_3_500  & Xd_0__inst_mult_3_504 )) # (Xd_0__inst_mult_3_496  & ((Xd_0__inst_mult_3_504 ) # (Xd_0__inst_mult_3_500 ))))

	.dataa(!Xd_0__inst_mult_3_496 ),
	.datab(!Xd_0__inst_mult_3_500 ),
	.datac(!Xd_0__inst_mult_3_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_353 ),
	.sharein(Xd_0__inst_mult_3_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_360 ),
	.cout(Xd_0__inst_mult_3_361 ),
	.shareout(Xd_0__inst_mult_3_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_105 (
// Equation(s):
// Xd_0__inst_mult_0_332  = SUM(( !Xd_0__inst_mult_0_460  $ (!Xd_0__inst_mult_0_464  $ (Xd_0__inst_mult_0_59_sumout )) ) + ( Xd_0__inst_mult_0_326  ) + ( Xd_0__inst_mult_0_325  ))
// Xd_0__inst_mult_0_333  = CARRY(( !Xd_0__inst_mult_0_460  $ (!Xd_0__inst_mult_0_464  $ (Xd_0__inst_mult_0_59_sumout )) ) + ( Xd_0__inst_mult_0_326  ) + ( Xd_0__inst_mult_0_325  ))
// Xd_0__inst_mult_0_334  = SHARE((!Xd_0__inst_mult_0_460  & (Xd_0__inst_mult_0_464  & Xd_0__inst_mult_0_59_sumout )) # (Xd_0__inst_mult_0_460  & ((Xd_0__inst_mult_0_59_sumout ) # (Xd_0__inst_mult_0_464 ))))

	.dataa(!Xd_0__inst_mult_0_460 ),
	.datab(!Xd_0__inst_mult_0_464 ),
	.datac(!Xd_0__inst_mult_0_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_325 ),
	.sharein(Xd_0__inst_mult_0_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_332 ),
	.cout(Xd_0__inst_mult_0_333 ),
	.shareout(Xd_0__inst_mult_0_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_106 (
// Equation(s):
// Xd_0__inst_mult_0_336  = SUM(( !Xd_0__inst_mult_0_468  $ (!Xd_0__inst_mult_0_472  $ (Xd_0__inst_mult_0_476 )) ) + ( Xd_0__inst_mult_0_330  ) + ( Xd_0__inst_mult_0_329  ))
// Xd_0__inst_mult_0_337  = CARRY(( !Xd_0__inst_mult_0_468  $ (!Xd_0__inst_mult_0_472  $ (Xd_0__inst_mult_0_476 )) ) + ( Xd_0__inst_mult_0_330  ) + ( Xd_0__inst_mult_0_329  ))
// Xd_0__inst_mult_0_338  = SHARE((!Xd_0__inst_mult_0_468  & (Xd_0__inst_mult_0_472  & Xd_0__inst_mult_0_476 )) # (Xd_0__inst_mult_0_468  & ((Xd_0__inst_mult_0_476 ) # (Xd_0__inst_mult_0_472 ))))

	.dataa(!Xd_0__inst_mult_0_468 ),
	.datab(!Xd_0__inst_mult_0_472 ),
	.datac(!Xd_0__inst_mult_0_476 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_329 ),
	.sharein(Xd_0__inst_mult_0_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_336 ),
	.cout(Xd_0__inst_mult_0_337 ),
	.shareout(Xd_0__inst_mult_0_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_101 (
// Equation(s):
// Xd_0__inst_mult_1_316  = SUM(( !Xd_0__inst_mult_1_444  $ (!Xd_0__inst_mult_1_448  $ (Xd_0__inst_mult_1_59_sumout )) ) + ( Xd_0__inst_mult_1_310  ) + ( Xd_0__inst_mult_1_309  ))
// Xd_0__inst_mult_1_317  = CARRY(( !Xd_0__inst_mult_1_444  $ (!Xd_0__inst_mult_1_448  $ (Xd_0__inst_mult_1_59_sumout )) ) + ( Xd_0__inst_mult_1_310  ) + ( Xd_0__inst_mult_1_309  ))
// Xd_0__inst_mult_1_318  = SHARE((!Xd_0__inst_mult_1_444  & (Xd_0__inst_mult_1_448  & Xd_0__inst_mult_1_59_sumout )) # (Xd_0__inst_mult_1_444  & ((Xd_0__inst_mult_1_59_sumout ) # (Xd_0__inst_mult_1_448 ))))

	.dataa(!Xd_0__inst_mult_1_444 ),
	.datab(!Xd_0__inst_mult_1_448 ),
	.datac(!Xd_0__inst_mult_1_59_sumout ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_309 ),
	.sharein(Xd_0__inst_mult_1_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_316 ),
	.cout(Xd_0__inst_mult_1_317 ),
	.shareout(Xd_0__inst_mult_1_318 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_102 (
// Equation(s):
// Xd_0__inst_mult_1_320  = SUM(( !Xd_0__inst_mult_1_452  $ (!Xd_0__inst_mult_1_456  $ (Xd_0__inst_mult_1_460 )) ) + ( Xd_0__inst_mult_1_314  ) + ( Xd_0__inst_mult_1_313  ))
// Xd_0__inst_mult_1_321  = CARRY(( !Xd_0__inst_mult_1_452  $ (!Xd_0__inst_mult_1_456  $ (Xd_0__inst_mult_1_460 )) ) + ( Xd_0__inst_mult_1_314  ) + ( Xd_0__inst_mult_1_313  ))
// Xd_0__inst_mult_1_322  = SHARE((!Xd_0__inst_mult_1_452  & (Xd_0__inst_mult_1_456  & Xd_0__inst_mult_1_460 )) # (Xd_0__inst_mult_1_452  & ((Xd_0__inst_mult_1_460 ) # (Xd_0__inst_mult_1_456 ))))

	.dataa(!Xd_0__inst_mult_1_452 ),
	.datab(!Xd_0__inst_mult_1_456 ),
	.datac(!Xd_0__inst_mult_1_460 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_313 ),
	.sharein(Xd_0__inst_mult_1_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_320 ),
	.cout(Xd_0__inst_mult_1_321 ),
	.shareout(Xd_0__inst_mult_1_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_139 (
// Equation(s):
// Xd_0__inst_mult_6_456  = SUM(( (din_a[80] & din_b[74]) ) + ( Xd_0__inst_mult_6_442  ) + ( Xd_0__inst_mult_6_441  ))
// Xd_0__inst_mult_6_457  = CARRY(( (din_a[80] & din_b[74]) ) + ( Xd_0__inst_mult_6_442  ) + ( Xd_0__inst_mult_6_441  ))
// Xd_0__inst_mult_6_458  = SHARE((din_a[82] & din_b[73]))

	.dataa(!din_a[80]),
	.datab(!din_b[74]),
	.datac(!din_a[82]),
	.datad(!din_b[73]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_441 ),
	.sharein(Xd_0__inst_mult_6_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_456 ),
	.cout(Xd_0__inst_mult_6_457 ),
	.shareout(Xd_0__inst_mult_6_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_140 (
// Equation(s):
// Xd_0__inst_mult_6_460  = SUM(( (!din_a[79] & (((din_a[78] & din_b[76])))) # (din_a[79] & (!din_b[75] $ (((!din_a[78]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_446  ) + ( Xd_0__inst_mult_6_445  ))
// Xd_0__inst_mult_6_461  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[76])))) # (din_a[79] & (!din_b[75] $ (((!din_a[78]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_446  ) + ( Xd_0__inst_mult_6_445  ))
// Xd_0__inst_mult_6_462  = SHARE((din_a[79] & (din_b[75] & (din_a[78] & din_b[76]))))

	.dataa(!din_a[79]),
	.datab(!din_b[75]),
	.datac(!din_a[78]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_445 ),
	.sharein(Xd_0__inst_mult_6_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_460 ),
	.cout(Xd_0__inst_mult_6_461 ),
	.shareout(Xd_0__inst_mult_6_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_67 (
// Equation(s):
// Xd_0__inst_mult_6_67_sumout  = SUM(( (din_a[82] & din_b[72]) ) + ( Xd_0__inst_mult_7_65  ) + ( Xd_0__inst_mult_7_64  ))
// Xd_0__inst_mult_6_68  = CARRY(( (din_a[82] & din_b[72]) ) + ( Xd_0__inst_mult_7_65  ) + ( Xd_0__inst_mult_7_64  ))
// Xd_0__inst_mult_6_69  = SHARE(GND)

	.dataa(!din_a[82]),
	.datab(!din_b[72]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_64 ),
	.sharein(Xd_0__inst_mult_7_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_67_sumout ),
	.cout(Xd_0__inst_mult_6_68 ),
	.shareout(Xd_0__inst_mult_6_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_141 (
// Equation(s):
// Xd_0__inst_mult_6_464  = SUM(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_6_450  ) + ( Xd_0__inst_mult_6_449  ))
// Xd_0__inst_mult_6_465  = CARRY(( (din_a[77] & din_b[77]) ) + ( Xd_0__inst_mult_6_450  ) + ( Xd_0__inst_mult_6_449  ))
// Xd_0__inst_mult_6_466  = SHARE((din_a[77] & din_b[78]))

	.dataa(!din_a[77]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_449 ),
	.sharein(Xd_0__inst_mult_6_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_464 ),
	.cout(Xd_0__inst_mult_6_465 ),
	.shareout(Xd_0__inst_mult_6_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_142 (
// Equation(s):
// Xd_0__inst_mult_6_468  = SUM(( (din_a[73] & din_b[81]) ) + ( Xd_0__inst_mult_6_454  ) + ( Xd_0__inst_mult_6_453  ))
// Xd_0__inst_mult_6_469  = CARRY(( (din_a[73] & din_b[81]) ) + ( Xd_0__inst_mult_6_454  ) + ( Xd_0__inst_mult_6_453  ))
// Xd_0__inst_mult_6_470  = SHARE((din_a[73] & din_b[82]))

	.dataa(!din_a[73]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_453 ),
	.sharein(Xd_0__inst_mult_6_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_468 ),
	.cout(Xd_0__inst_mult_6_469 ),
	.shareout(Xd_0__inst_mult_6_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_143 (
// Equation(s):
// Xd_0__inst_mult_6_472  = SUM(( (!din_a[75] & (((din_a[74] & din_b[80])))) # (din_a[75] & (!din_b[79] $ (((!din_a[74]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_582  ) + ( Xd_0__inst_mult_6_581  ))
// Xd_0__inst_mult_6_473  = CARRY(( (!din_a[75] & (((din_a[74] & din_b[80])))) # (din_a[75] & (!din_b[79] $ (((!din_a[74]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_582  ) + ( Xd_0__inst_mult_6_581  ))
// Xd_0__inst_mult_6_474  = SHARE((din_a[75] & (din_b[79] & (din_a[74] & din_b[80]))))

	.dataa(!din_a[75]),
	.datab(!din_b[79]),
	.datac(!din_a[74]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_581 ),
	.sharein(Xd_0__inst_mult_6_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_472 ),
	.cout(Xd_0__inst_mult_6_473 ),
	.shareout(Xd_0__inst_mult_6_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_141 (
// Equation(s):
// Xd_0__inst_mult_7_464  = SUM(( (din_a[92] & din_b[86]) ) + ( Xd_0__inst_mult_7_450  ) + ( Xd_0__inst_mult_7_449  ))
// Xd_0__inst_mult_7_465  = CARRY(( (din_a[92] & din_b[86]) ) + ( Xd_0__inst_mult_7_450  ) + ( Xd_0__inst_mult_7_449  ))
// Xd_0__inst_mult_7_466  = SHARE((din_a[94] & din_b[85]))

	.dataa(!din_a[92]),
	.datab(!din_b[86]),
	.datac(!din_a[94]),
	.datad(!din_b[85]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_449 ),
	.sharein(Xd_0__inst_mult_7_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_464 ),
	.cout(Xd_0__inst_mult_7_465 ),
	.shareout(Xd_0__inst_mult_7_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_142 (
// Equation(s):
// Xd_0__inst_mult_7_468  = SUM(( (!din_a[91] & (((din_a[90] & din_b[88])))) # (din_a[91] & (!din_b[87] $ (((!din_a[90]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_454  ) + ( Xd_0__inst_mult_7_453  ))
// Xd_0__inst_mult_7_469  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[88])))) # (din_a[91] & (!din_b[87] $ (((!din_a[90]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_454  ) + ( Xd_0__inst_mult_7_453  ))
// Xd_0__inst_mult_7_470  = SHARE((din_a[91] & (din_b[87] & (din_a[90] & din_b[88]))))

	.dataa(!din_a[91]),
	.datab(!din_b[87]),
	.datac(!din_a[90]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_453 ),
	.sharein(Xd_0__inst_mult_7_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_468 ),
	.cout(Xd_0__inst_mult_7_469 ),
	.shareout(Xd_0__inst_mult_7_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_67 (
// Equation(s):
// Xd_0__inst_mult_7_67_sumout  = SUM(( (din_a[94] & din_b[84]) ) + ( Xd_0__inst_mult_6_69  ) + ( Xd_0__inst_mult_6_68  ))
// Xd_0__inst_mult_7_68  = CARRY(( (din_a[94] & din_b[84]) ) + ( Xd_0__inst_mult_6_69  ) + ( Xd_0__inst_mult_6_68  ))
// Xd_0__inst_mult_7_69  = SHARE(GND)

	.dataa(!din_a[94]),
	.datab(!din_b[84]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_68 ),
	.sharein(Xd_0__inst_mult_6_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_67_sumout ),
	.cout(Xd_0__inst_mult_7_68 ),
	.shareout(Xd_0__inst_mult_7_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_143 (
// Equation(s):
// Xd_0__inst_mult_7_472  = SUM(( (din_a[89] & din_b[89]) ) + ( Xd_0__inst_mult_7_458  ) + ( Xd_0__inst_mult_7_457  ))
// Xd_0__inst_mult_7_473  = CARRY(( (din_a[89] & din_b[89]) ) + ( Xd_0__inst_mult_7_458  ) + ( Xd_0__inst_mult_7_457  ))
// Xd_0__inst_mult_7_474  = SHARE((din_a[89] & din_b[90]))

	.dataa(!din_a[89]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_457 ),
	.sharein(Xd_0__inst_mult_7_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_472 ),
	.cout(Xd_0__inst_mult_7_473 ),
	.shareout(Xd_0__inst_mult_7_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_144 (
// Equation(s):
// Xd_0__inst_mult_7_476  = SUM(( (din_a[85] & din_b[93]) ) + ( Xd_0__inst_mult_7_462  ) + ( Xd_0__inst_mult_7_461  ))
// Xd_0__inst_mult_7_477  = CARRY(( (din_a[85] & din_b[93]) ) + ( Xd_0__inst_mult_7_462  ) + ( Xd_0__inst_mult_7_461  ))
// Xd_0__inst_mult_7_478  = SHARE((din_a[85] & din_b[94]))

	.dataa(!din_a[85]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_461 ),
	.sharein(Xd_0__inst_mult_7_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_476 ),
	.cout(Xd_0__inst_mult_7_477 ),
	.shareout(Xd_0__inst_mult_7_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_145 (
// Equation(s):
// Xd_0__inst_mult_7_480  = SUM(( (!din_a[87] & (((din_a[86] & din_b[92])))) # (din_a[87] & (!din_b[91] $ (((!din_a[86]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_582  ) + ( Xd_0__inst_mult_7_581  ))
// Xd_0__inst_mult_7_481  = CARRY(( (!din_a[87] & (((din_a[86] & din_b[92])))) # (din_a[87] & (!din_b[91] $ (((!din_a[86]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_582  ) + ( Xd_0__inst_mult_7_581  ))
// Xd_0__inst_mult_7_482  = SHARE((din_a[87] & (din_b[91] & (din_a[86] & din_b[92]))))

	.dataa(!din_a[87]),
	.datab(!din_b[91]),
	.datac(!din_a[86]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_581 ),
	.sharein(Xd_0__inst_mult_7_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_480 ),
	.cout(Xd_0__inst_mult_7_481 ),
	.shareout(Xd_0__inst_mult_7_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_105 (
// Equation(s):
// Xd_0__inst_mult_4_320  = SUM(( !Xd_0__inst_mult_4_472  $ (!Xd_0__inst_mult_4_476 ) ) + ( Xd_0__inst_mult_4_314  ) + ( Xd_0__inst_mult_4_313  ))
// Xd_0__inst_mult_4_321  = CARRY(( !Xd_0__inst_mult_4_472  $ (!Xd_0__inst_mult_4_476 ) ) + ( Xd_0__inst_mult_4_314  ) + ( Xd_0__inst_mult_4_313  ))
// Xd_0__inst_mult_4_322  = SHARE((Xd_0__inst_mult_4_472  & Xd_0__inst_mult_4_476 ))

	.dataa(!Xd_0__inst_mult_4_472 ),
	.datab(!Xd_0__inst_mult_4_476 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_313 ),
	.sharein(Xd_0__inst_mult_4_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_320 ),
	.cout(Xd_0__inst_mult_4_321 ),
	.shareout(Xd_0__inst_mult_4_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_106 (
// Equation(s):
// Xd_0__inst_mult_4_324  = SUM(( !Xd_0__inst_mult_4_480  $ (!Xd_0__inst_mult_4_484  $ (Xd_0__inst_mult_4_488 )) ) + ( Xd_0__inst_mult_4_318  ) + ( Xd_0__inst_mult_4_317  ))
// Xd_0__inst_mult_4_325  = CARRY(( !Xd_0__inst_mult_4_480  $ (!Xd_0__inst_mult_4_484  $ (Xd_0__inst_mult_4_488 )) ) + ( Xd_0__inst_mult_4_318  ) + ( Xd_0__inst_mult_4_317  ))
// Xd_0__inst_mult_4_326  = SHARE((!Xd_0__inst_mult_4_480  & (Xd_0__inst_mult_4_484  & Xd_0__inst_mult_4_488 )) # (Xd_0__inst_mult_4_480  & ((Xd_0__inst_mult_4_488 ) # (Xd_0__inst_mult_4_484 ))))

	.dataa(!Xd_0__inst_mult_4_480 ),
	.datab(!Xd_0__inst_mult_4_484 ),
	.datac(!Xd_0__inst_mult_4_488 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_317 ),
	.sharein(Xd_0__inst_mult_4_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_324 ),
	.cout(Xd_0__inst_mult_4_325 ),
	.shareout(Xd_0__inst_mult_4_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_105 (
// Equation(s):
// Xd_0__inst_mult_5_320  = SUM(( !Xd_0__inst_mult_5_468  $ (!Xd_0__inst_mult_5_472 ) ) + ( Xd_0__inst_mult_5_314  ) + ( Xd_0__inst_mult_5_313  ))
// Xd_0__inst_mult_5_321  = CARRY(( !Xd_0__inst_mult_5_468  $ (!Xd_0__inst_mult_5_472 ) ) + ( Xd_0__inst_mult_5_314  ) + ( Xd_0__inst_mult_5_313  ))
// Xd_0__inst_mult_5_322  = SHARE((Xd_0__inst_mult_5_468  & Xd_0__inst_mult_5_472 ))

	.dataa(!Xd_0__inst_mult_5_468 ),
	.datab(!Xd_0__inst_mult_5_472 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_313 ),
	.sharein(Xd_0__inst_mult_5_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_320 ),
	.cout(Xd_0__inst_mult_5_321 ),
	.shareout(Xd_0__inst_mult_5_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_106 (
// Equation(s):
// Xd_0__inst_mult_5_324  = SUM(( !Xd_0__inst_mult_5_476  $ (!Xd_0__inst_mult_5_480  $ (Xd_0__inst_mult_5_484 )) ) + ( Xd_0__inst_mult_5_318  ) + ( Xd_0__inst_mult_5_317  ))
// Xd_0__inst_mult_5_325  = CARRY(( !Xd_0__inst_mult_5_476  $ (!Xd_0__inst_mult_5_480  $ (Xd_0__inst_mult_5_484 )) ) + ( Xd_0__inst_mult_5_318  ) + ( Xd_0__inst_mult_5_317  ))
// Xd_0__inst_mult_5_326  = SHARE((!Xd_0__inst_mult_5_476  & (Xd_0__inst_mult_5_480  & Xd_0__inst_mult_5_484 )) # (Xd_0__inst_mult_5_476  & ((Xd_0__inst_mult_5_484 ) # (Xd_0__inst_mult_5_480 ))))

	.dataa(!Xd_0__inst_mult_5_476 ),
	.datab(!Xd_0__inst_mult_5_480 ),
	.datac(!Xd_0__inst_mult_5_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_317 ),
	.sharein(Xd_0__inst_mult_5_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_324 ),
	.cout(Xd_0__inst_mult_5_325 ),
	.shareout(Xd_0__inst_mult_5_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_105 (
// Equation(s):
// Xd_0__inst_mult_2_320  = SUM(( !Xd_0__inst_mult_2_468  $ (!Xd_0__inst_mult_2_472 ) ) + ( Xd_0__inst_mult_2_314  ) + ( Xd_0__inst_mult_2_313  ))
// Xd_0__inst_mult_2_321  = CARRY(( !Xd_0__inst_mult_2_468  $ (!Xd_0__inst_mult_2_472 ) ) + ( Xd_0__inst_mult_2_314  ) + ( Xd_0__inst_mult_2_313  ))
// Xd_0__inst_mult_2_322  = SHARE((Xd_0__inst_mult_2_468  & Xd_0__inst_mult_2_472 ))

	.dataa(!Xd_0__inst_mult_2_468 ),
	.datab(!Xd_0__inst_mult_2_472 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_313 ),
	.sharein(Xd_0__inst_mult_2_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_320 ),
	.cout(Xd_0__inst_mult_2_321 ),
	.shareout(Xd_0__inst_mult_2_322 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_106 (
// Equation(s):
// Xd_0__inst_mult_2_324  = SUM(( !Xd_0__inst_mult_2_476  $ (!Xd_0__inst_mult_2_480  $ (Xd_0__inst_mult_2_484 )) ) + ( Xd_0__inst_mult_2_318  ) + ( Xd_0__inst_mult_2_317  ))
// Xd_0__inst_mult_2_325  = CARRY(( !Xd_0__inst_mult_2_476  $ (!Xd_0__inst_mult_2_480  $ (Xd_0__inst_mult_2_484 )) ) + ( Xd_0__inst_mult_2_318  ) + ( Xd_0__inst_mult_2_317  ))
// Xd_0__inst_mult_2_326  = SHARE((!Xd_0__inst_mult_2_476  & (Xd_0__inst_mult_2_480  & Xd_0__inst_mult_2_484 )) # (Xd_0__inst_mult_2_476  & ((Xd_0__inst_mult_2_484 ) # (Xd_0__inst_mult_2_480 ))))

	.dataa(!Xd_0__inst_mult_2_476 ),
	.datab(!Xd_0__inst_mult_2_480 ),
	.datac(!Xd_0__inst_mult_2_484 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_317 ),
	.sharein(Xd_0__inst_mult_2_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_324 ),
	.cout(Xd_0__inst_mult_2_325 ),
	.shareout(Xd_0__inst_mult_2_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_113 (
// Equation(s):
// Xd_0__inst_mult_3_364  = SUM(( !Xd_0__inst_mult_3_508  $ (!Xd_0__inst_mult_3_512 ) ) + ( Xd_0__inst_mult_3_358  ) + ( Xd_0__inst_mult_3_357  ))
// Xd_0__inst_mult_3_365  = CARRY(( !Xd_0__inst_mult_3_508  $ (!Xd_0__inst_mult_3_512 ) ) + ( Xd_0__inst_mult_3_358  ) + ( Xd_0__inst_mult_3_357  ))
// Xd_0__inst_mult_3_366  = SHARE((Xd_0__inst_mult_3_508  & Xd_0__inst_mult_3_512 ))

	.dataa(!Xd_0__inst_mult_3_508 ),
	.datab(!Xd_0__inst_mult_3_512 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_357 ),
	.sharein(Xd_0__inst_mult_3_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_364 ),
	.cout(Xd_0__inst_mult_3_365 ),
	.shareout(Xd_0__inst_mult_3_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_114 (
// Equation(s):
// Xd_0__inst_mult_3_368  = SUM(( !Xd_0__inst_mult_3_516  $ (!Xd_0__inst_mult_3_520  $ (Xd_0__inst_mult_3_524 )) ) + ( Xd_0__inst_mult_3_362  ) + ( Xd_0__inst_mult_3_361  ))
// Xd_0__inst_mult_3_369  = CARRY(( !Xd_0__inst_mult_3_516  $ (!Xd_0__inst_mult_3_520  $ (Xd_0__inst_mult_3_524 )) ) + ( Xd_0__inst_mult_3_362  ) + ( Xd_0__inst_mult_3_361  ))
// Xd_0__inst_mult_3_370  = SHARE((!Xd_0__inst_mult_3_516  & (Xd_0__inst_mult_3_520  & Xd_0__inst_mult_3_524 )) # (Xd_0__inst_mult_3_516  & ((Xd_0__inst_mult_3_524 ) # (Xd_0__inst_mult_3_520 ))))

	.dataa(!Xd_0__inst_mult_3_516 ),
	.datab(!Xd_0__inst_mult_3_520 ),
	.datac(!Xd_0__inst_mult_3_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_361 ),
	.sharein(Xd_0__inst_mult_3_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_368 ),
	.cout(Xd_0__inst_mult_3_369 ),
	.shareout(Xd_0__inst_mult_3_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_107 (
// Equation(s):
// Xd_0__inst_mult_0_340  = SUM(( !Xd_0__inst_mult_0_480  $ (!Xd_0__inst_mult_0_484 ) ) + ( Xd_0__inst_mult_0_334  ) + ( Xd_0__inst_mult_0_333  ))
// Xd_0__inst_mult_0_341  = CARRY(( !Xd_0__inst_mult_0_480  $ (!Xd_0__inst_mult_0_484 ) ) + ( Xd_0__inst_mult_0_334  ) + ( Xd_0__inst_mult_0_333  ))
// Xd_0__inst_mult_0_342  = SHARE((Xd_0__inst_mult_0_480  & Xd_0__inst_mult_0_484 ))

	.dataa(!Xd_0__inst_mult_0_480 ),
	.datab(!Xd_0__inst_mult_0_484 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_333 ),
	.sharein(Xd_0__inst_mult_0_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_340 ),
	.cout(Xd_0__inst_mult_0_341 ),
	.shareout(Xd_0__inst_mult_0_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_108 (
// Equation(s):
// Xd_0__inst_mult_0_344  = SUM(( !Xd_0__inst_mult_0_488  $ (!Xd_0__inst_mult_0_492  $ (Xd_0__inst_mult_0_496 )) ) + ( Xd_0__inst_mult_0_338  ) + ( Xd_0__inst_mult_0_337  ))
// Xd_0__inst_mult_0_345  = CARRY(( !Xd_0__inst_mult_0_488  $ (!Xd_0__inst_mult_0_492  $ (Xd_0__inst_mult_0_496 )) ) + ( Xd_0__inst_mult_0_338  ) + ( Xd_0__inst_mult_0_337  ))
// Xd_0__inst_mult_0_346  = SHARE((!Xd_0__inst_mult_0_488  & (Xd_0__inst_mult_0_492  & Xd_0__inst_mult_0_496 )) # (Xd_0__inst_mult_0_488  & ((Xd_0__inst_mult_0_496 ) # (Xd_0__inst_mult_0_492 ))))

	.dataa(!Xd_0__inst_mult_0_488 ),
	.datab(!Xd_0__inst_mult_0_492 ),
	.datac(!Xd_0__inst_mult_0_496 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_337 ),
	.sharein(Xd_0__inst_mult_0_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_344 ),
	.cout(Xd_0__inst_mult_0_345 ),
	.shareout(Xd_0__inst_mult_0_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_103 (
// Equation(s):
// Xd_0__inst_mult_1_324  = SUM(( !Xd_0__inst_mult_1_464  $ (!Xd_0__inst_mult_1_468 ) ) + ( Xd_0__inst_mult_1_318  ) + ( Xd_0__inst_mult_1_317  ))
// Xd_0__inst_mult_1_325  = CARRY(( !Xd_0__inst_mult_1_464  $ (!Xd_0__inst_mult_1_468 ) ) + ( Xd_0__inst_mult_1_318  ) + ( Xd_0__inst_mult_1_317  ))
// Xd_0__inst_mult_1_326  = SHARE((Xd_0__inst_mult_1_464  & Xd_0__inst_mult_1_468 ))

	.dataa(!Xd_0__inst_mult_1_464 ),
	.datab(!Xd_0__inst_mult_1_468 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_317 ),
	.sharein(Xd_0__inst_mult_1_318 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_324 ),
	.cout(Xd_0__inst_mult_1_325 ),
	.shareout(Xd_0__inst_mult_1_326 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_104 (
// Equation(s):
// Xd_0__inst_mult_1_328  = SUM(( !Xd_0__inst_mult_1_472  $ (!Xd_0__inst_mult_1_476  $ (Xd_0__inst_mult_1_480 )) ) + ( Xd_0__inst_mult_1_322  ) + ( Xd_0__inst_mult_1_321  ))
// Xd_0__inst_mult_1_329  = CARRY(( !Xd_0__inst_mult_1_472  $ (!Xd_0__inst_mult_1_476  $ (Xd_0__inst_mult_1_480 )) ) + ( Xd_0__inst_mult_1_322  ) + ( Xd_0__inst_mult_1_321  ))
// Xd_0__inst_mult_1_330  = SHARE((!Xd_0__inst_mult_1_472  & (Xd_0__inst_mult_1_476  & Xd_0__inst_mult_1_480 )) # (Xd_0__inst_mult_1_472  & ((Xd_0__inst_mult_1_480 ) # (Xd_0__inst_mult_1_476 ))))

	.dataa(!Xd_0__inst_mult_1_472 ),
	.datab(!Xd_0__inst_mult_1_476 ),
	.datac(!Xd_0__inst_mult_1_480 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_321 ),
	.sharein(Xd_0__inst_mult_1_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_328 ),
	.cout(Xd_0__inst_mult_1_329 ),
	.shareout(Xd_0__inst_mult_1_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_144 (
// Equation(s):
// Xd_0__inst_mult_6_476  = SUM(( (din_a[81] & din_b[74]) ) + ( Xd_0__inst_mult_6_458  ) + ( Xd_0__inst_mult_6_457  ))
// Xd_0__inst_mult_6_477  = CARRY(( (din_a[81] & din_b[74]) ) + ( Xd_0__inst_mult_6_458  ) + ( Xd_0__inst_mult_6_457  ))
// Xd_0__inst_mult_6_478  = SHARE(GND)

	.dataa(!din_a[81]),
	.datab(!din_b[74]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_457 ),
	.sharein(Xd_0__inst_mult_6_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_476 ),
	.cout(Xd_0__inst_mult_6_477 ),
	.shareout(Xd_0__inst_mult_6_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_145 (
// Equation(s):
// Xd_0__inst_mult_6_480  = SUM(( (!din_a[80] & (((din_a[79] & din_b[76])))) # (din_a[80] & (!din_b[75] $ (((!din_a[79]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_462  ) + ( Xd_0__inst_mult_6_461  ))
// Xd_0__inst_mult_6_481  = CARRY(( (!din_a[80] & (((din_a[79] & din_b[76])))) # (din_a[80] & (!din_b[75] $ (((!din_a[79]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_462  ) + ( Xd_0__inst_mult_6_461  ))
// Xd_0__inst_mult_6_482  = SHARE((din_a[80] & (din_b[75] & (din_a[79] & din_b[76]))))

	.dataa(!din_a[80]),
	.datab(!din_b[75]),
	.datac(!din_a[79]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_461 ),
	.sharein(Xd_0__inst_mult_6_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_480 ),
	.cout(Xd_0__inst_mult_6_481 ),
	.shareout(Xd_0__inst_mult_6_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_146 (
// Equation(s):
// Xd_0__inst_mult_6_484  = SUM(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_6_466  ) + ( Xd_0__inst_mult_6_465  ))
// Xd_0__inst_mult_6_485  = CARRY(( (din_a[78] & din_b[77]) ) + ( Xd_0__inst_mult_6_466  ) + ( Xd_0__inst_mult_6_465  ))
// Xd_0__inst_mult_6_486  = SHARE((din_a[78] & din_b[78]))

	.dataa(!din_a[78]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_465 ),
	.sharein(Xd_0__inst_mult_6_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_484 ),
	.cout(Xd_0__inst_mult_6_485 ),
	.shareout(Xd_0__inst_mult_6_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_147 (
// Equation(s):
// Xd_0__inst_mult_6_488  = SUM(( (din_a[74] & din_b[81]) ) + ( Xd_0__inst_mult_6_470  ) + ( Xd_0__inst_mult_6_469  ))
// Xd_0__inst_mult_6_489  = CARRY(( (din_a[74] & din_b[81]) ) + ( Xd_0__inst_mult_6_470  ) + ( Xd_0__inst_mult_6_469  ))
// Xd_0__inst_mult_6_490  = SHARE((din_a[74] & din_b[82]))

	.dataa(!din_a[74]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_469 ),
	.sharein(Xd_0__inst_mult_6_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_488 ),
	.cout(Xd_0__inst_mult_6_489 ),
	.shareout(Xd_0__inst_mult_6_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_148 (
// Equation(s):
// Xd_0__inst_mult_6_492  = SUM(( (!din_a[76] & (((din_a[75] & din_b[80])))) # (din_a[76] & (!din_b[79] $ (((!din_a[75]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_474  ) + ( Xd_0__inst_mult_6_473  ))
// Xd_0__inst_mult_6_493  = CARRY(( (!din_a[76] & (((din_a[75] & din_b[80])))) # (din_a[76] & (!din_b[79] $ (((!din_a[75]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_474  ) + ( Xd_0__inst_mult_6_473  ))
// Xd_0__inst_mult_6_494  = SHARE((din_a[76] & (din_b[79] & (din_a[75] & din_b[80]))))

	.dataa(!din_a[76]),
	.datab(!din_b[79]),
	.datac(!din_a[75]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_473 ),
	.sharein(Xd_0__inst_mult_6_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_492 ),
	.cout(Xd_0__inst_mult_6_493 ),
	.shareout(Xd_0__inst_mult_6_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_146 (
// Equation(s):
// Xd_0__inst_mult_7_484  = SUM(( (din_a[93] & din_b[86]) ) + ( Xd_0__inst_mult_7_466  ) + ( Xd_0__inst_mult_7_465  ))
// Xd_0__inst_mult_7_485  = CARRY(( (din_a[93] & din_b[86]) ) + ( Xd_0__inst_mult_7_466  ) + ( Xd_0__inst_mult_7_465  ))
// Xd_0__inst_mult_7_486  = SHARE(GND)

	.dataa(!din_a[93]),
	.datab(!din_b[86]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_465 ),
	.sharein(Xd_0__inst_mult_7_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_484 ),
	.cout(Xd_0__inst_mult_7_485 ),
	.shareout(Xd_0__inst_mult_7_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_147 (
// Equation(s):
// Xd_0__inst_mult_7_488  = SUM(( (!din_a[92] & (((din_a[91] & din_b[88])))) # (din_a[92] & (!din_b[87] $ (((!din_a[91]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_470  ) + ( Xd_0__inst_mult_7_469  ))
// Xd_0__inst_mult_7_489  = CARRY(( (!din_a[92] & (((din_a[91] & din_b[88])))) # (din_a[92] & (!din_b[87] $ (((!din_a[91]) # (!din_b[88]))))) ) + ( Xd_0__inst_mult_7_470  ) + ( Xd_0__inst_mult_7_469  ))
// Xd_0__inst_mult_7_490  = SHARE((din_a[92] & (din_b[87] & (din_a[91] & din_b[88]))))

	.dataa(!din_a[92]),
	.datab(!din_b[87]),
	.datac(!din_a[91]),
	.datad(!din_b[88]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_469 ),
	.sharein(Xd_0__inst_mult_7_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_488 ),
	.cout(Xd_0__inst_mult_7_489 ),
	.shareout(Xd_0__inst_mult_7_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_148 (
// Equation(s):
// Xd_0__inst_mult_7_492  = SUM(( (din_a[90] & din_b[89]) ) + ( Xd_0__inst_mult_7_474  ) + ( Xd_0__inst_mult_7_473  ))
// Xd_0__inst_mult_7_493  = CARRY(( (din_a[90] & din_b[89]) ) + ( Xd_0__inst_mult_7_474  ) + ( Xd_0__inst_mult_7_473  ))
// Xd_0__inst_mult_7_494  = SHARE((din_a[90] & din_b[90]))

	.dataa(!din_a[90]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_473 ),
	.sharein(Xd_0__inst_mult_7_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_492 ),
	.cout(Xd_0__inst_mult_7_493 ),
	.shareout(Xd_0__inst_mult_7_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_149 (
// Equation(s):
// Xd_0__inst_mult_7_496  = SUM(( (din_a[86] & din_b[93]) ) + ( Xd_0__inst_mult_7_478  ) + ( Xd_0__inst_mult_7_477  ))
// Xd_0__inst_mult_7_497  = CARRY(( (din_a[86] & din_b[93]) ) + ( Xd_0__inst_mult_7_478  ) + ( Xd_0__inst_mult_7_477  ))
// Xd_0__inst_mult_7_498  = SHARE((din_a[86] & din_b[94]))

	.dataa(!din_a[86]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_477 ),
	.sharein(Xd_0__inst_mult_7_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_496 ),
	.cout(Xd_0__inst_mult_7_497 ),
	.shareout(Xd_0__inst_mult_7_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_150 (
// Equation(s):
// Xd_0__inst_mult_7_500  = SUM(( (!din_a[88] & (((din_a[87] & din_b[92])))) # (din_a[88] & (!din_b[91] $ (((!din_a[87]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_482  ) + ( Xd_0__inst_mult_7_481  ))
// Xd_0__inst_mult_7_501  = CARRY(( (!din_a[88] & (((din_a[87] & din_b[92])))) # (din_a[88] & (!din_b[91] $ (((!din_a[87]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_482  ) + ( Xd_0__inst_mult_7_481  ))
// Xd_0__inst_mult_7_502  = SHARE((din_a[88] & (din_b[91] & (din_a[87] & din_b[92]))))

	.dataa(!din_a[88]),
	.datab(!din_b[91]),
	.datac(!din_a[87]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_481 ),
	.sharein(Xd_0__inst_mult_7_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_500 ),
	.cout(Xd_0__inst_mult_7_501 ),
	.shareout(Xd_0__inst_mult_7_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_107 (
// Equation(s):
// Xd_0__inst_mult_4_328  = SUM(( !Xd_0__inst_mult_4_492  $ (!Xd_0__inst_mult_4_496  $ (((din_b[50] & din_a[58])))) ) + ( Xd_0__inst_mult_4_322  ) + ( Xd_0__inst_mult_4_321  ))
// Xd_0__inst_mult_4_329  = CARRY(( !Xd_0__inst_mult_4_492  $ (!Xd_0__inst_mult_4_496  $ (((din_b[50] & din_a[58])))) ) + ( Xd_0__inst_mult_4_322  ) + ( Xd_0__inst_mult_4_321  ))
// Xd_0__inst_mult_4_330  = SHARE((!Xd_0__inst_mult_4_492  & (Xd_0__inst_mult_4_496  & (din_b[50] & din_a[58]))) # (Xd_0__inst_mult_4_492  & (((din_b[50] & din_a[58])) # (Xd_0__inst_mult_4_496 ))))

	.dataa(!Xd_0__inst_mult_4_492 ),
	.datab(!Xd_0__inst_mult_4_496 ),
	.datac(!din_b[50]),
	.datad(!din_a[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_321 ),
	.sharein(Xd_0__inst_mult_4_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_328 ),
	.cout(Xd_0__inst_mult_4_329 ),
	.shareout(Xd_0__inst_mult_4_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_108 (
// Equation(s):
// Xd_0__inst_mult_4_332  = SUM(( !Xd_0__inst_mult_4_500  $ (!Xd_0__inst_mult_4_504  $ (Xd_0__inst_mult_4_508 )) ) + ( Xd_0__inst_mult_4_326  ) + ( Xd_0__inst_mult_4_325  ))
// Xd_0__inst_mult_4_333  = CARRY(( !Xd_0__inst_mult_4_500  $ (!Xd_0__inst_mult_4_504  $ (Xd_0__inst_mult_4_508 )) ) + ( Xd_0__inst_mult_4_326  ) + ( Xd_0__inst_mult_4_325  ))
// Xd_0__inst_mult_4_334  = SHARE((!Xd_0__inst_mult_4_500  & (Xd_0__inst_mult_4_504  & Xd_0__inst_mult_4_508 )) # (Xd_0__inst_mult_4_500  & ((Xd_0__inst_mult_4_508 ) # (Xd_0__inst_mult_4_504 ))))

	.dataa(!Xd_0__inst_mult_4_500 ),
	.datab(!Xd_0__inst_mult_4_504 ),
	.datac(!Xd_0__inst_mult_4_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_325 ),
	.sharein(Xd_0__inst_mult_4_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_332 ),
	.cout(Xd_0__inst_mult_4_333 ),
	.shareout(Xd_0__inst_mult_4_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_107 (
// Equation(s):
// Xd_0__inst_mult_5_328  = SUM(( !Xd_0__inst_mult_5_488  $ (!Xd_0__inst_mult_5_492  $ (((din_b[62] & din_a[70])))) ) + ( Xd_0__inst_mult_5_322  ) + ( Xd_0__inst_mult_5_321  ))
// Xd_0__inst_mult_5_329  = CARRY(( !Xd_0__inst_mult_5_488  $ (!Xd_0__inst_mult_5_492  $ (((din_b[62] & din_a[70])))) ) + ( Xd_0__inst_mult_5_322  ) + ( Xd_0__inst_mult_5_321  ))
// Xd_0__inst_mult_5_330  = SHARE((!Xd_0__inst_mult_5_488  & (Xd_0__inst_mult_5_492  & (din_b[62] & din_a[70]))) # (Xd_0__inst_mult_5_488  & (((din_b[62] & din_a[70])) # (Xd_0__inst_mult_5_492 ))))

	.dataa(!Xd_0__inst_mult_5_488 ),
	.datab(!Xd_0__inst_mult_5_492 ),
	.datac(!din_b[62]),
	.datad(!din_a[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_321 ),
	.sharein(Xd_0__inst_mult_5_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_328 ),
	.cout(Xd_0__inst_mult_5_329 ),
	.shareout(Xd_0__inst_mult_5_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_108 (
// Equation(s):
// Xd_0__inst_mult_5_332  = SUM(( !Xd_0__inst_mult_5_496  $ (!Xd_0__inst_mult_5_500  $ (Xd_0__inst_mult_5_504 )) ) + ( Xd_0__inst_mult_5_326  ) + ( Xd_0__inst_mult_5_325  ))
// Xd_0__inst_mult_5_333  = CARRY(( !Xd_0__inst_mult_5_496  $ (!Xd_0__inst_mult_5_500  $ (Xd_0__inst_mult_5_504 )) ) + ( Xd_0__inst_mult_5_326  ) + ( Xd_0__inst_mult_5_325  ))
// Xd_0__inst_mult_5_334  = SHARE((!Xd_0__inst_mult_5_496  & (Xd_0__inst_mult_5_500  & Xd_0__inst_mult_5_504 )) # (Xd_0__inst_mult_5_496  & ((Xd_0__inst_mult_5_504 ) # (Xd_0__inst_mult_5_500 ))))

	.dataa(!Xd_0__inst_mult_5_496 ),
	.datab(!Xd_0__inst_mult_5_500 ),
	.datac(!Xd_0__inst_mult_5_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_325 ),
	.sharein(Xd_0__inst_mult_5_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_332 ),
	.cout(Xd_0__inst_mult_5_333 ),
	.shareout(Xd_0__inst_mult_5_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_107 (
// Equation(s):
// Xd_0__inst_mult_2_328  = SUM(( !Xd_0__inst_mult_2_488  $ (!Xd_0__inst_mult_2_492  $ (((din_b[26] & din_a[34])))) ) + ( Xd_0__inst_mult_2_322  ) + ( Xd_0__inst_mult_2_321  ))
// Xd_0__inst_mult_2_329  = CARRY(( !Xd_0__inst_mult_2_488  $ (!Xd_0__inst_mult_2_492  $ (((din_b[26] & din_a[34])))) ) + ( Xd_0__inst_mult_2_322  ) + ( Xd_0__inst_mult_2_321  ))
// Xd_0__inst_mult_2_330  = SHARE((!Xd_0__inst_mult_2_488  & (Xd_0__inst_mult_2_492  & (din_b[26] & din_a[34]))) # (Xd_0__inst_mult_2_488  & (((din_b[26] & din_a[34])) # (Xd_0__inst_mult_2_492 ))))

	.dataa(!Xd_0__inst_mult_2_488 ),
	.datab(!Xd_0__inst_mult_2_492 ),
	.datac(!din_b[26]),
	.datad(!din_a[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_321 ),
	.sharein(Xd_0__inst_mult_2_322 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_328 ),
	.cout(Xd_0__inst_mult_2_329 ),
	.shareout(Xd_0__inst_mult_2_330 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_108 (
// Equation(s):
// Xd_0__inst_mult_2_332  = SUM(( !Xd_0__inst_mult_2_496  $ (!Xd_0__inst_mult_2_500  $ (Xd_0__inst_mult_2_504 )) ) + ( Xd_0__inst_mult_2_326  ) + ( Xd_0__inst_mult_2_325  ))
// Xd_0__inst_mult_2_333  = CARRY(( !Xd_0__inst_mult_2_496  $ (!Xd_0__inst_mult_2_500  $ (Xd_0__inst_mult_2_504 )) ) + ( Xd_0__inst_mult_2_326  ) + ( Xd_0__inst_mult_2_325  ))
// Xd_0__inst_mult_2_334  = SHARE((!Xd_0__inst_mult_2_496  & (Xd_0__inst_mult_2_500  & Xd_0__inst_mult_2_504 )) # (Xd_0__inst_mult_2_496  & ((Xd_0__inst_mult_2_504 ) # (Xd_0__inst_mult_2_500 ))))

	.dataa(!Xd_0__inst_mult_2_496 ),
	.datab(!Xd_0__inst_mult_2_500 ),
	.datac(!Xd_0__inst_mult_2_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_325 ),
	.sharein(Xd_0__inst_mult_2_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_332 ),
	.cout(Xd_0__inst_mult_2_333 ),
	.shareout(Xd_0__inst_mult_2_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_115 (
// Equation(s):
// Xd_0__inst_mult_3_372  = SUM(( !Xd_0__inst_mult_3_528  $ (!Xd_0__inst_mult_3_532  $ (Xd_0__inst_mult_3_536 )) ) + ( Xd_0__inst_mult_3_370  ) + ( Xd_0__inst_mult_3_369  ))
// Xd_0__inst_mult_3_373  = CARRY(( !Xd_0__inst_mult_3_528  $ (!Xd_0__inst_mult_3_532  $ (Xd_0__inst_mult_3_536 )) ) + ( Xd_0__inst_mult_3_370  ) + ( Xd_0__inst_mult_3_369  ))
// Xd_0__inst_mult_3_374  = SHARE((!Xd_0__inst_mult_3_528  & (Xd_0__inst_mult_3_532  & Xd_0__inst_mult_3_536 )) # (Xd_0__inst_mult_3_528  & ((Xd_0__inst_mult_3_536 ) # (Xd_0__inst_mult_3_532 ))))

	.dataa(!Xd_0__inst_mult_3_528 ),
	.datab(!Xd_0__inst_mult_3_532 ),
	.datac(!Xd_0__inst_mult_3_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_369 ),
	.sharein(Xd_0__inst_mult_3_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_372 ),
	.cout(Xd_0__inst_mult_3_373 ),
	.shareout(Xd_0__inst_mult_3_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_109 (
// Equation(s):
// Xd_0__inst_mult_0_348  = SUM(( !Xd_0__inst_mult_0_500  $ (!Xd_0__inst_mult_0_504  $ (Xd_0__inst_mult_0_508 )) ) + ( Xd_0__inst_mult_0_346  ) + ( Xd_0__inst_mult_0_345  ))
// Xd_0__inst_mult_0_349  = CARRY(( !Xd_0__inst_mult_0_500  $ (!Xd_0__inst_mult_0_504  $ (Xd_0__inst_mult_0_508 )) ) + ( Xd_0__inst_mult_0_346  ) + ( Xd_0__inst_mult_0_345  ))
// Xd_0__inst_mult_0_350  = SHARE((!Xd_0__inst_mult_0_500  & (Xd_0__inst_mult_0_504  & Xd_0__inst_mult_0_508 )) # (Xd_0__inst_mult_0_500  & ((Xd_0__inst_mult_0_508 ) # (Xd_0__inst_mult_0_504 ))))

	.dataa(!Xd_0__inst_mult_0_500 ),
	.datab(!Xd_0__inst_mult_0_504 ),
	.datac(!Xd_0__inst_mult_0_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_345 ),
	.sharein(Xd_0__inst_mult_0_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_348 ),
	.cout(Xd_0__inst_mult_0_349 ),
	.shareout(Xd_0__inst_mult_0_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_105 (
// Equation(s):
// Xd_0__inst_mult_1_332  = SUM(( !Xd_0__inst_mult_1_484  $ (!Xd_0__inst_mult_1_488  $ (((din_b[14] & din_a[22])))) ) + ( Xd_0__inst_mult_1_326  ) + ( Xd_0__inst_mult_1_325  ))
// Xd_0__inst_mult_1_333  = CARRY(( !Xd_0__inst_mult_1_484  $ (!Xd_0__inst_mult_1_488  $ (((din_b[14] & din_a[22])))) ) + ( Xd_0__inst_mult_1_326  ) + ( Xd_0__inst_mult_1_325  ))
// Xd_0__inst_mult_1_334  = SHARE((!Xd_0__inst_mult_1_484  & (Xd_0__inst_mult_1_488  & (din_b[14] & din_a[22]))) # (Xd_0__inst_mult_1_484  & (((din_b[14] & din_a[22])) # (Xd_0__inst_mult_1_488 ))))

	.dataa(!Xd_0__inst_mult_1_484 ),
	.datab(!Xd_0__inst_mult_1_488 ),
	.datac(!din_b[14]),
	.datad(!din_a[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_325 ),
	.sharein(Xd_0__inst_mult_1_326 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_332 ),
	.cout(Xd_0__inst_mult_1_333 ),
	.shareout(Xd_0__inst_mult_1_334 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_106 (
// Equation(s):
// Xd_0__inst_mult_1_336  = SUM(( !Xd_0__inst_mult_1_492  $ (!Xd_0__inst_mult_1_496  $ (Xd_0__inst_mult_1_500 )) ) + ( Xd_0__inst_mult_1_330  ) + ( Xd_0__inst_mult_1_329  ))
// Xd_0__inst_mult_1_337  = CARRY(( !Xd_0__inst_mult_1_492  $ (!Xd_0__inst_mult_1_496  $ (Xd_0__inst_mult_1_500 )) ) + ( Xd_0__inst_mult_1_330  ) + ( Xd_0__inst_mult_1_329  ))
// Xd_0__inst_mult_1_338  = SHARE((!Xd_0__inst_mult_1_492  & (Xd_0__inst_mult_1_496  & Xd_0__inst_mult_1_500 )) # (Xd_0__inst_mult_1_492  & ((Xd_0__inst_mult_1_500 ) # (Xd_0__inst_mult_1_496 ))))

	.dataa(!Xd_0__inst_mult_1_492 ),
	.datab(!Xd_0__inst_mult_1_496 ),
	.datac(!Xd_0__inst_mult_1_500 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_329 ),
	.sharein(Xd_0__inst_mult_1_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_336 ),
	.cout(Xd_0__inst_mult_1_337 ),
	.shareout(Xd_0__inst_mult_1_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_149 (
// Equation(s):
// Xd_0__inst_mult_6_496  = SUM(( GND ) + ( Xd_0__inst_mult_6_478  ) + ( Xd_0__inst_mult_6_477  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_477 ),
	.sharein(Xd_0__inst_mult_6_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_496 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_150 (
// Equation(s):
// Xd_0__inst_mult_6_500  = SUM(( (!din_a[81] & (((din_a[80] & din_b[76])))) # (din_a[81] & (!din_b[75] $ (((!din_a[80]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_482  ) + ( Xd_0__inst_mult_6_481  ))
// Xd_0__inst_mult_6_501  = CARRY(( (!din_a[81] & (((din_a[80] & din_b[76])))) # (din_a[81] & (!din_b[75] $ (((!din_a[80]) # (!din_b[76]))))) ) + ( Xd_0__inst_mult_6_482  ) + ( Xd_0__inst_mult_6_481  ))
// Xd_0__inst_mult_6_502  = SHARE((din_a[81] & (din_b[75] & (din_a[80] & din_b[76]))))

	.dataa(!din_a[81]),
	.datab(!din_b[75]),
	.datac(!din_a[80]),
	.datad(!din_b[76]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_481 ),
	.sharein(Xd_0__inst_mult_6_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_500 ),
	.cout(Xd_0__inst_mult_6_501 ),
	.shareout(Xd_0__inst_mult_6_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_151 (
// Equation(s):
// Xd_0__inst_mult_6_504  = SUM(( (din_a[79] & din_b[77]) ) + ( Xd_0__inst_mult_6_486  ) + ( Xd_0__inst_mult_6_485  ))
// Xd_0__inst_mult_6_505  = CARRY(( (din_a[79] & din_b[77]) ) + ( Xd_0__inst_mult_6_486  ) + ( Xd_0__inst_mult_6_485  ))
// Xd_0__inst_mult_6_506  = SHARE((din_a[79] & din_b[78]))

	.dataa(!din_a[79]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_485 ),
	.sharein(Xd_0__inst_mult_6_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_504 ),
	.cout(Xd_0__inst_mult_6_505 ),
	.shareout(Xd_0__inst_mult_6_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_152 (
// Equation(s):
// Xd_0__inst_mult_6_508  = SUM(( (din_a[75] & din_b[81]) ) + ( Xd_0__inst_mult_6_490  ) + ( Xd_0__inst_mult_6_489  ))
// Xd_0__inst_mult_6_509  = CARRY(( (din_a[75] & din_b[81]) ) + ( Xd_0__inst_mult_6_490  ) + ( Xd_0__inst_mult_6_489  ))
// Xd_0__inst_mult_6_510  = SHARE((din_a[75] & din_b[82]))

	.dataa(!din_a[75]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_489 ),
	.sharein(Xd_0__inst_mult_6_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_508 ),
	.cout(Xd_0__inst_mult_6_509 ),
	.shareout(Xd_0__inst_mult_6_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_153 (
// Equation(s):
// Xd_0__inst_mult_6_512  = SUM(( (!din_a[77] & (((din_a[76] & din_b[80])))) # (din_a[77] & (!din_b[79] $ (((!din_a[76]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_494  ) + ( Xd_0__inst_mult_6_493  ))
// Xd_0__inst_mult_6_513  = CARRY(( (!din_a[77] & (((din_a[76] & din_b[80])))) # (din_a[77] & (!din_b[79] $ (((!din_a[76]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_494  ) + ( Xd_0__inst_mult_6_493  ))
// Xd_0__inst_mult_6_514  = SHARE((din_a[77] & (din_b[79] & (din_a[76] & din_b[80]))))

	.dataa(!din_a[77]),
	.datab(!din_b[79]),
	.datac(!din_a[76]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_493 ),
	.sharein(Xd_0__inst_mult_6_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_512 ),
	.cout(Xd_0__inst_mult_6_513 ),
	.shareout(Xd_0__inst_mult_6_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_151 (
// Equation(s):
// Xd_0__inst_mult_7_504  = SUM(( (din_a[91] & din_b[89]) ) + ( Xd_0__inst_mult_7_494  ) + ( Xd_0__inst_mult_7_493  ))
// Xd_0__inst_mult_7_505  = CARRY(( (din_a[91] & din_b[89]) ) + ( Xd_0__inst_mult_7_494  ) + ( Xd_0__inst_mult_7_493  ))
// Xd_0__inst_mult_7_506  = SHARE((din_a[91] & din_b[90]))

	.dataa(!din_a[91]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_493 ),
	.sharein(Xd_0__inst_mult_7_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_504 ),
	.cout(Xd_0__inst_mult_7_505 ),
	.shareout(Xd_0__inst_mult_7_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_152 (
// Equation(s):
// Xd_0__inst_mult_7_508  = SUM(( (din_a[87] & din_b[93]) ) + ( Xd_0__inst_mult_7_498  ) + ( Xd_0__inst_mult_7_497  ))
// Xd_0__inst_mult_7_509  = CARRY(( (din_a[87] & din_b[93]) ) + ( Xd_0__inst_mult_7_498  ) + ( Xd_0__inst_mult_7_497  ))
// Xd_0__inst_mult_7_510  = SHARE((din_a[87] & din_b[94]))

	.dataa(!din_a[87]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_497 ),
	.sharein(Xd_0__inst_mult_7_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_508 ),
	.cout(Xd_0__inst_mult_7_509 ),
	.shareout(Xd_0__inst_mult_7_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_153 (
// Equation(s):
// Xd_0__inst_mult_7_512  = SUM(( (!din_a[89] & (((din_a[88] & din_b[92])))) # (din_a[89] & (!din_b[91] $ (((!din_a[88]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_502  ) + ( Xd_0__inst_mult_7_501  ))
// Xd_0__inst_mult_7_513  = CARRY(( (!din_a[89] & (((din_a[88] & din_b[92])))) # (din_a[89] & (!din_b[91] $ (((!din_a[88]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_502  ) + ( Xd_0__inst_mult_7_501  ))
// Xd_0__inst_mult_7_514  = SHARE((din_a[89] & (din_b[91] & (din_a[88] & din_b[92]))))

	.dataa(!din_a[89]),
	.datab(!din_b[91]),
	.datac(!din_a[88]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_501 ),
	.sharein(Xd_0__inst_mult_7_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_512 ),
	.cout(Xd_0__inst_mult_7_513 ),
	.shareout(Xd_0__inst_mult_7_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_109 (
// Equation(s):
// Xd_0__inst_mult_4_336  = SUM(( !Xd_0__inst_mult_4_512  $ (((!din_b[51]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_330  ) + ( Xd_0__inst_mult_4_329  ))
// Xd_0__inst_mult_4_337  = CARRY(( !Xd_0__inst_mult_4_512  $ (((!din_b[51]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_330  ) + ( Xd_0__inst_mult_4_329  ))
// Xd_0__inst_mult_4_338  = SHARE((din_b[51] & (din_a[58] & Xd_0__inst_mult_4_512 )))

	.dataa(!din_b[51]),
	.datab(!din_a[58]),
	.datac(!Xd_0__inst_mult_4_512 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_329 ),
	.sharein(Xd_0__inst_mult_4_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_336 ),
	.cout(Xd_0__inst_mult_4_337 ),
	.shareout(Xd_0__inst_mult_4_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_110 (
// Equation(s):
// Xd_0__inst_mult_4_340  = SUM(( !Xd_0__inst_mult_4_516  $ (!Xd_0__inst_mult_4_520  $ (Xd_0__inst_mult_4_524 )) ) + ( Xd_0__inst_mult_4_334  ) + ( Xd_0__inst_mult_4_333  ))
// Xd_0__inst_mult_4_341  = CARRY(( !Xd_0__inst_mult_4_516  $ (!Xd_0__inst_mult_4_520  $ (Xd_0__inst_mult_4_524 )) ) + ( Xd_0__inst_mult_4_334  ) + ( Xd_0__inst_mult_4_333  ))
// Xd_0__inst_mult_4_342  = SHARE((!Xd_0__inst_mult_4_516  & (Xd_0__inst_mult_4_520  & Xd_0__inst_mult_4_524 )) # (Xd_0__inst_mult_4_516  & ((Xd_0__inst_mult_4_524 ) # (Xd_0__inst_mult_4_520 ))))

	.dataa(!Xd_0__inst_mult_4_516 ),
	.datab(!Xd_0__inst_mult_4_520 ),
	.datac(!Xd_0__inst_mult_4_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_333 ),
	.sharein(Xd_0__inst_mult_4_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_340 ),
	.cout(Xd_0__inst_mult_4_341 ),
	.shareout(Xd_0__inst_mult_4_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_109 (
// Equation(s):
// Xd_0__inst_mult_5_336  = SUM(( !Xd_0__inst_mult_5_508  $ (((!din_b[63]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_330  ) + ( Xd_0__inst_mult_5_329  ))
// Xd_0__inst_mult_5_337  = CARRY(( !Xd_0__inst_mult_5_508  $ (((!din_b[63]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_330  ) + ( Xd_0__inst_mult_5_329  ))
// Xd_0__inst_mult_5_338  = SHARE((din_b[63] & (din_a[70] & Xd_0__inst_mult_5_508 )))

	.dataa(!din_b[63]),
	.datab(!din_a[70]),
	.datac(!Xd_0__inst_mult_5_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_329 ),
	.sharein(Xd_0__inst_mult_5_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_336 ),
	.cout(Xd_0__inst_mult_5_337 ),
	.shareout(Xd_0__inst_mult_5_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_110 (
// Equation(s):
// Xd_0__inst_mult_5_340  = SUM(( !Xd_0__inst_mult_5_512  $ (!Xd_0__inst_mult_5_516  $ (Xd_0__inst_mult_5_520 )) ) + ( Xd_0__inst_mult_5_334  ) + ( Xd_0__inst_mult_5_333  ))
// Xd_0__inst_mult_5_341  = CARRY(( !Xd_0__inst_mult_5_512  $ (!Xd_0__inst_mult_5_516  $ (Xd_0__inst_mult_5_520 )) ) + ( Xd_0__inst_mult_5_334  ) + ( Xd_0__inst_mult_5_333  ))
// Xd_0__inst_mult_5_342  = SHARE((!Xd_0__inst_mult_5_512  & (Xd_0__inst_mult_5_516  & Xd_0__inst_mult_5_520 )) # (Xd_0__inst_mult_5_512  & ((Xd_0__inst_mult_5_520 ) # (Xd_0__inst_mult_5_516 ))))

	.dataa(!Xd_0__inst_mult_5_512 ),
	.datab(!Xd_0__inst_mult_5_516 ),
	.datac(!Xd_0__inst_mult_5_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_333 ),
	.sharein(Xd_0__inst_mult_5_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_340 ),
	.cout(Xd_0__inst_mult_5_341 ),
	.shareout(Xd_0__inst_mult_5_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_109 (
// Equation(s):
// Xd_0__inst_mult_2_336  = SUM(( !Xd_0__inst_mult_2_508  $ (((!din_b[27]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_330  ) + ( Xd_0__inst_mult_2_329  ))
// Xd_0__inst_mult_2_337  = CARRY(( !Xd_0__inst_mult_2_508  $ (((!din_b[27]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_330  ) + ( Xd_0__inst_mult_2_329  ))
// Xd_0__inst_mult_2_338  = SHARE((din_b[27] & (din_a[34] & Xd_0__inst_mult_2_508 )))

	.dataa(!din_b[27]),
	.datab(!din_a[34]),
	.datac(!Xd_0__inst_mult_2_508 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_329 ),
	.sharein(Xd_0__inst_mult_2_330 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_336 ),
	.cout(Xd_0__inst_mult_2_337 ),
	.shareout(Xd_0__inst_mult_2_338 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_110 (
// Equation(s):
// Xd_0__inst_mult_2_340  = SUM(( !Xd_0__inst_mult_2_512  $ (!Xd_0__inst_mult_2_516  $ (Xd_0__inst_mult_2_520 )) ) + ( Xd_0__inst_mult_2_334  ) + ( Xd_0__inst_mult_2_333  ))
// Xd_0__inst_mult_2_341  = CARRY(( !Xd_0__inst_mult_2_512  $ (!Xd_0__inst_mult_2_516  $ (Xd_0__inst_mult_2_520 )) ) + ( Xd_0__inst_mult_2_334  ) + ( Xd_0__inst_mult_2_333  ))
// Xd_0__inst_mult_2_342  = SHARE((!Xd_0__inst_mult_2_512  & (Xd_0__inst_mult_2_516  & Xd_0__inst_mult_2_520 )) # (Xd_0__inst_mult_2_512  & ((Xd_0__inst_mult_2_520 ) # (Xd_0__inst_mult_2_516 ))))

	.dataa(!Xd_0__inst_mult_2_512 ),
	.datab(!Xd_0__inst_mult_2_516 ),
	.datac(!Xd_0__inst_mult_2_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_333 ),
	.sharein(Xd_0__inst_mult_2_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_340 ),
	.cout(Xd_0__inst_mult_2_341 ),
	.shareout(Xd_0__inst_mult_2_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_116 (
// Equation(s):
// Xd_0__inst_mult_3_376  = SUM(( !Xd_0__inst_mult_3_540  $ (!Xd_0__inst_mult_3_416  $ (Xd_0__inst_mult_3_544 )) ) + ( Xd_0__inst_mult_3_374  ) + ( Xd_0__inst_mult_3_373  ))
// Xd_0__inst_mult_3_377  = CARRY(( !Xd_0__inst_mult_3_540  $ (!Xd_0__inst_mult_3_416  $ (Xd_0__inst_mult_3_544 )) ) + ( Xd_0__inst_mult_3_374  ) + ( Xd_0__inst_mult_3_373  ))
// Xd_0__inst_mult_3_378  = SHARE((!Xd_0__inst_mult_3_540  & (Xd_0__inst_mult_3_416  & Xd_0__inst_mult_3_544 )) # (Xd_0__inst_mult_3_540  & ((Xd_0__inst_mult_3_544 ) # (Xd_0__inst_mult_3_416 ))))

	.dataa(!Xd_0__inst_mult_3_540 ),
	.datab(!Xd_0__inst_mult_3_416 ),
	.datac(!Xd_0__inst_mult_3_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_373 ),
	.sharein(Xd_0__inst_mult_3_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_376 ),
	.cout(Xd_0__inst_mult_3_377 ),
	.shareout(Xd_0__inst_mult_3_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_110 (
// Equation(s):
// Xd_0__inst_mult_0_352  = SUM(( !Xd_0__inst_mult_0_512  $ (!Xd_0__inst_mult_0_516  $ (Xd_0__inst_mult_0_520 )) ) + ( Xd_0__inst_mult_0_350  ) + ( Xd_0__inst_mult_0_349  ))
// Xd_0__inst_mult_0_353  = CARRY(( !Xd_0__inst_mult_0_512  $ (!Xd_0__inst_mult_0_516  $ (Xd_0__inst_mult_0_520 )) ) + ( Xd_0__inst_mult_0_350  ) + ( Xd_0__inst_mult_0_349  ))
// Xd_0__inst_mult_0_354  = SHARE((!Xd_0__inst_mult_0_512  & (Xd_0__inst_mult_0_516  & Xd_0__inst_mult_0_520 )) # (Xd_0__inst_mult_0_512  & ((Xd_0__inst_mult_0_520 ) # (Xd_0__inst_mult_0_516 ))))

	.dataa(!Xd_0__inst_mult_0_512 ),
	.datab(!Xd_0__inst_mult_0_516 ),
	.datac(!Xd_0__inst_mult_0_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_349 ),
	.sharein(Xd_0__inst_mult_0_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_352 ),
	.cout(Xd_0__inst_mult_0_353 ),
	.shareout(Xd_0__inst_mult_0_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_107 (
// Equation(s):
// Xd_0__inst_mult_1_340  = SUM(( !Xd_0__inst_mult_1_504  $ (((!din_b[15]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_334  ) + ( Xd_0__inst_mult_1_333  ))
// Xd_0__inst_mult_1_341  = CARRY(( !Xd_0__inst_mult_1_504  $ (((!din_b[15]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_334  ) + ( Xd_0__inst_mult_1_333  ))
// Xd_0__inst_mult_1_342  = SHARE((din_b[15] & (din_a[22] & Xd_0__inst_mult_1_504 )))

	.dataa(!din_b[15]),
	.datab(!din_a[22]),
	.datac(!Xd_0__inst_mult_1_504 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_333 ),
	.sharein(Xd_0__inst_mult_1_334 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_340 ),
	.cout(Xd_0__inst_mult_1_341 ),
	.shareout(Xd_0__inst_mult_1_342 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_108 (
// Equation(s):
// Xd_0__inst_mult_1_344  = SUM(( !Xd_0__inst_mult_1_508  $ (!Xd_0__inst_mult_1_512  $ (Xd_0__inst_mult_1_516 )) ) + ( Xd_0__inst_mult_1_338  ) + ( Xd_0__inst_mult_1_337  ))
// Xd_0__inst_mult_1_345  = CARRY(( !Xd_0__inst_mult_1_508  $ (!Xd_0__inst_mult_1_512  $ (Xd_0__inst_mult_1_516 )) ) + ( Xd_0__inst_mult_1_338  ) + ( Xd_0__inst_mult_1_337  ))
// Xd_0__inst_mult_1_346  = SHARE((!Xd_0__inst_mult_1_508  & (Xd_0__inst_mult_1_512  & Xd_0__inst_mult_1_516 )) # (Xd_0__inst_mult_1_508  & ((Xd_0__inst_mult_1_516 ) # (Xd_0__inst_mult_1_512 ))))

	.dataa(!Xd_0__inst_mult_1_508 ),
	.datab(!Xd_0__inst_mult_1_512 ),
	.datac(!Xd_0__inst_mult_1_516 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_337 ),
	.sharein(Xd_0__inst_mult_1_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_344 ),
	.cout(Xd_0__inst_mult_1_345 ),
	.shareout(Xd_0__inst_mult_1_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_154 (
// Equation(s):
// Xd_0__inst_mult_6_516  = SUM(( (din_a[80] & din_b[77]) ) + ( Xd_0__inst_mult_6_506  ) + ( Xd_0__inst_mult_6_505  ))
// Xd_0__inst_mult_6_517  = CARRY(( (din_a[80] & din_b[77]) ) + ( Xd_0__inst_mult_6_506  ) + ( Xd_0__inst_mult_6_505  ))
// Xd_0__inst_mult_6_518  = SHARE((din_a[80] & din_b[78]))

	.dataa(!din_a[80]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_505 ),
	.sharein(Xd_0__inst_mult_6_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_516 ),
	.cout(Xd_0__inst_mult_6_517 ),
	.shareout(Xd_0__inst_mult_6_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_155 (
// Equation(s):
// Xd_0__inst_mult_6_520  = SUM(( (din_a[76] & din_b[81]) ) + ( Xd_0__inst_mult_6_510  ) + ( Xd_0__inst_mult_6_509  ))
// Xd_0__inst_mult_6_521  = CARRY(( (din_a[76] & din_b[81]) ) + ( Xd_0__inst_mult_6_510  ) + ( Xd_0__inst_mult_6_509  ))
// Xd_0__inst_mult_6_522  = SHARE((din_a[76] & din_b[82]))

	.dataa(!din_a[76]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_509 ),
	.sharein(Xd_0__inst_mult_6_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_520 ),
	.cout(Xd_0__inst_mult_6_521 ),
	.shareout(Xd_0__inst_mult_6_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_156 (
// Equation(s):
// Xd_0__inst_mult_6_524  = SUM(( (!din_a[78] & (((din_a[77] & din_b[80])))) # (din_a[78] & (!din_b[79] $ (((!din_a[77]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_514  ) + ( Xd_0__inst_mult_6_513  ))
// Xd_0__inst_mult_6_525  = CARRY(( (!din_a[78] & (((din_a[77] & din_b[80])))) # (din_a[78] & (!din_b[79] $ (((!din_a[77]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_514  ) + ( Xd_0__inst_mult_6_513  ))
// Xd_0__inst_mult_6_526  = SHARE((din_a[78] & (din_b[79] & (din_a[77] & din_b[80]))))

	.dataa(!din_a[78]),
	.datab(!din_b[79]),
	.datac(!din_a[77]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_513 ),
	.sharein(Xd_0__inst_mult_6_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_524 ),
	.cout(Xd_0__inst_mult_6_525 ),
	.shareout(Xd_0__inst_mult_6_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_154 (
// Equation(s):
// Xd_0__inst_mult_7_516  = SUM(( (din_a[92] & din_b[89]) ) + ( Xd_0__inst_mult_7_506  ) + ( Xd_0__inst_mult_7_505  ))
// Xd_0__inst_mult_7_517  = CARRY(( (din_a[92] & din_b[89]) ) + ( Xd_0__inst_mult_7_506  ) + ( Xd_0__inst_mult_7_505  ))
// Xd_0__inst_mult_7_518  = SHARE((din_a[92] & din_b[90]))

	.dataa(!din_a[92]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_505 ),
	.sharein(Xd_0__inst_mult_7_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_516 ),
	.cout(Xd_0__inst_mult_7_517 ),
	.shareout(Xd_0__inst_mult_7_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_155 (
// Equation(s):
// Xd_0__inst_mult_7_520  = SUM(( (din_a[88] & din_b[93]) ) + ( Xd_0__inst_mult_7_510  ) + ( Xd_0__inst_mult_7_509  ))
// Xd_0__inst_mult_7_521  = CARRY(( (din_a[88] & din_b[93]) ) + ( Xd_0__inst_mult_7_510  ) + ( Xd_0__inst_mult_7_509  ))
// Xd_0__inst_mult_7_522  = SHARE((din_a[88] & din_b[94]))

	.dataa(!din_a[88]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_509 ),
	.sharein(Xd_0__inst_mult_7_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_520 ),
	.cout(Xd_0__inst_mult_7_521 ),
	.shareout(Xd_0__inst_mult_7_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_156 (
// Equation(s):
// Xd_0__inst_mult_7_524  = SUM(( (!din_a[90] & (((din_a[89] & din_b[92])))) # (din_a[90] & (!din_b[91] $ (((!din_a[89]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_514  ) + ( Xd_0__inst_mult_7_513  ))
// Xd_0__inst_mult_7_525  = CARRY(( (!din_a[90] & (((din_a[89] & din_b[92])))) # (din_a[90] & (!din_b[91] $ (((!din_a[89]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_514  ) + ( Xd_0__inst_mult_7_513  ))
// Xd_0__inst_mult_7_526  = SHARE((din_a[90] & (din_b[91] & (din_a[89] & din_b[92]))))

	.dataa(!din_a[90]),
	.datab(!din_b[91]),
	.datac(!din_a[89]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_513 ),
	.sharein(Xd_0__inst_mult_7_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_524 ),
	.cout(Xd_0__inst_mult_7_525 ),
	.shareout(Xd_0__inst_mult_7_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_111 (
// Equation(s):
// Xd_0__inst_mult_4_344  = SUM(( !Xd_0__inst_mult_4_528  $ (((!din_b[52]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_338  ) + ( Xd_0__inst_mult_4_337  ))
// Xd_0__inst_mult_4_345  = CARRY(( !Xd_0__inst_mult_4_528  $ (((!din_b[52]) # (!din_a[58]))) ) + ( Xd_0__inst_mult_4_338  ) + ( Xd_0__inst_mult_4_337  ))
// Xd_0__inst_mult_4_346  = SHARE((din_b[52] & (din_a[58] & Xd_0__inst_mult_4_528 )))

	.dataa(!din_b[52]),
	.datab(!din_a[58]),
	.datac(!Xd_0__inst_mult_4_528 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_337 ),
	.sharein(Xd_0__inst_mult_4_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_344 ),
	.cout(Xd_0__inst_mult_4_345 ),
	.shareout(Xd_0__inst_mult_4_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_112 (
// Equation(s):
// Xd_0__inst_mult_4_348  = SUM(( !Xd_0__inst_mult_4_532  $ (!Xd_0__inst_mult_4_536  $ (Xd_0__inst_mult_4_540 )) ) + ( Xd_0__inst_mult_4_342  ) + ( Xd_0__inst_mult_4_341  ))
// Xd_0__inst_mult_4_349  = CARRY(( !Xd_0__inst_mult_4_532  $ (!Xd_0__inst_mult_4_536  $ (Xd_0__inst_mult_4_540 )) ) + ( Xd_0__inst_mult_4_342  ) + ( Xd_0__inst_mult_4_341  ))
// Xd_0__inst_mult_4_350  = SHARE((!Xd_0__inst_mult_4_532  & (Xd_0__inst_mult_4_536  & Xd_0__inst_mult_4_540 )) # (Xd_0__inst_mult_4_532  & ((Xd_0__inst_mult_4_540 ) # (Xd_0__inst_mult_4_536 ))))

	.dataa(!Xd_0__inst_mult_4_532 ),
	.datab(!Xd_0__inst_mult_4_536 ),
	.datac(!Xd_0__inst_mult_4_540 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_341 ),
	.sharein(Xd_0__inst_mult_4_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_348 ),
	.cout(Xd_0__inst_mult_4_349 ),
	.shareout(Xd_0__inst_mult_4_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_111 (
// Equation(s):
// Xd_0__inst_mult_5_344  = SUM(( !Xd_0__inst_mult_5_524  $ (((!din_b[64]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_338  ) + ( Xd_0__inst_mult_5_337  ))
// Xd_0__inst_mult_5_345  = CARRY(( !Xd_0__inst_mult_5_524  $ (((!din_b[64]) # (!din_a[70]))) ) + ( Xd_0__inst_mult_5_338  ) + ( Xd_0__inst_mult_5_337  ))
// Xd_0__inst_mult_5_346  = SHARE((din_b[64] & (din_a[70] & Xd_0__inst_mult_5_524 )))

	.dataa(!din_b[64]),
	.datab(!din_a[70]),
	.datac(!Xd_0__inst_mult_5_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_337 ),
	.sharein(Xd_0__inst_mult_5_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_344 ),
	.cout(Xd_0__inst_mult_5_345 ),
	.shareout(Xd_0__inst_mult_5_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_112 (
// Equation(s):
// Xd_0__inst_mult_5_348  = SUM(( !Xd_0__inst_mult_5_528  $ (!Xd_0__inst_mult_5_532  $ (Xd_0__inst_mult_5_536 )) ) + ( Xd_0__inst_mult_5_342  ) + ( Xd_0__inst_mult_5_341  ))
// Xd_0__inst_mult_5_349  = CARRY(( !Xd_0__inst_mult_5_528  $ (!Xd_0__inst_mult_5_532  $ (Xd_0__inst_mult_5_536 )) ) + ( Xd_0__inst_mult_5_342  ) + ( Xd_0__inst_mult_5_341  ))
// Xd_0__inst_mult_5_350  = SHARE((!Xd_0__inst_mult_5_528  & (Xd_0__inst_mult_5_532  & Xd_0__inst_mult_5_536 )) # (Xd_0__inst_mult_5_528  & ((Xd_0__inst_mult_5_536 ) # (Xd_0__inst_mult_5_532 ))))

	.dataa(!Xd_0__inst_mult_5_528 ),
	.datab(!Xd_0__inst_mult_5_532 ),
	.datac(!Xd_0__inst_mult_5_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_341 ),
	.sharein(Xd_0__inst_mult_5_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_348 ),
	.cout(Xd_0__inst_mult_5_349 ),
	.shareout(Xd_0__inst_mult_5_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_111 (
// Equation(s):
// Xd_0__inst_mult_2_344  = SUM(( !Xd_0__inst_mult_2_524  $ (((!din_b[28]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_338  ) + ( Xd_0__inst_mult_2_337  ))
// Xd_0__inst_mult_2_345  = CARRY(( !Xd_0__inst_mult_2_524  $ (((!din_b[28]) # (!din_a[34]))) ) + ( Xd_0__inst_mult_2_338  ) + ( Xd_0__inst_mult_2_337  ))
// Xd_0__inst_mult_2_346  = SHARE((din_b[28] & (din_a[34] & Xd_0__inst_mult_2_524 )))

	.dataa(!din_b[28]),
	.datab(!din_a[34]),
	.datac(!Xd_0__inst_mult_2_524 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_337 ),
	.sharein(Xd_0__inst_mult_2_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_344 ),
	.cout(Xd_0__inst_mult_2_345 ),
	.shareout(Xd_0__inst_mult_2_346 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_112 (
// Equation(s):
// Xd_0__inst_mult_2_348  = SUM(( !Xd_0__inst_mult_2_528  $ (!Xd_0__inst_mult_2_532  $ (Xd_0__inst_mult_2_536 )) ) + ( Xd_0__inst_mult_2_342  ) + ( Xd_0__inst_mult_2_341  ))
// Xd_0__inst_mult_2_349  = CARRY(( !Xd_0__inst_mult_2_528  $ (!Xd_0__inst_mult_2_532  $ (Xd_0__inst_mult_2_536 )) ) + ( Xd_0__inst_mult_2_342  ) + ( Xd_0__inst_mult_2_341  ))
// Xd_0__inst_mult_2_350  = SHARE((!Xd_0__inst_mult_2_528  & (Xd_0__inst_mult_2_532  & Xd_0__inst_mult_2_536 )) # (Xd_0__inst_mult_2_528  & ((Xd_0__inst_mult_2_536 ) # (Xd_0__inst_mult_2_532 ))))

	.dataa(!Xd_0__inst_mult_2_528 ),
	.datab(!Xd_0__inst_mult_2_532 ),
	.datac(!Xd_0__inst_mult_2_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_341 ),
	.sharein(Xd_0__inst_mult_2_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_348 ),
	.cout(Xd_0__inst_mult_2_349 ),
	.shareout(Xd_0__inst_mult_2_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_117 (
// Equation(s):
// Xd_0__inst_mult_3_380  = SUM(( !Xd_0__inst_mult_3_548  $ (!Xd_0__inst_mult_3_300  $ (Xd_0__inst_mult_3_552 )) ) + ( Xd_0__inst_mult_3_378  ) + ( Xd_0__inst_mult_3_377  ))
// Xd_0__inst_mult_3_381  = CARRY(( !Xd_0__inst_mult_3_548  $ (!Xd_0__inst_mult_3_300  $ (Xd_0__inst_mult_3_552 )) ) + ( Xd_0__inst_mult_3_378  ) + ( Xd_0__inst_mult_3_377  ))
// Xd_0__inst_mult_3_382  = SHARE((!Xd_0__inst_mult_3_548  & (Xd_0__inst_mult_3_300  & Xd_0__inst_mult_3_552 )) # (Xd_0__inst_mult_3_548  & ((Xd_0__inst_mult_3_552 ) # (Xd_0__inst_mult_3_300 ))))

	.dataa(!Xd_0__inst_mult_3_548 ),
	.datab(!Xd_0__inst_mult_3_300 ),
	.datac(!Xd_0__inst_mult_3_552 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_377 ),
	.sharein(Xd_0__inst_mult_3_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_380 ),
	.cout(Xd_0__inst_mult_3_381 ),
	.shareout(Xd_0__inst_mult_3_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_111 (
// Equation(s):
// Xd_0__inst_mult_0_356  = SUM(( !Xd_0__inst_mult_0_524  $ (!Xd_0__inst_mult_0_528  $ (Xd_0__inst_mult_0_532 )) ) + ( Xd_0__inst_mult_0_354  ) + ( Xd_0__inst_mult_0_353  ))
// Xd_0__inst_mult_0_357  = CARRY(( !Xd_0__inst_mult_0_524  $ (!Xd_0__inst_mult_0_528  $ (Xd_0__inst_mult_0_532 )) ) + ( Xd_0__inst_mult_0_354  ) + ( Xd_0__inst_mult_0_353  ))
// Xd_0__inst_mult_0_358  = SHARE((!Xd_0__inst_mult_0_524  & (Xd_0__inst_mult_0_528  & Xd_0__inst_mult_0_532 )) # (Xd_0__inst_mult_0_524  & ((Xd_0__inst_mult_0_532 ) # (Xd_0__inst_mult_0_528 ))))

	.dataa(!Xd_0__inst_mult_0_524 ),
	.datab(!Xd_0__inst_mult_0_528 ),
	.datac(!Xd_0__inst_mult_0_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_353 ),
	.sharein(Xd_0__inst_mult_0_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_356 ),
	.cout(Xd_0__inst_mult_0_357 ),
	.shareout(Xd_0__inst_mult_0_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_109 (
// Equation(s):
// Xd_0__inst_mult_1_348  = SUM(( !Xd_0__inst_mult_1_520  $ (((!din_b[16]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_342  ) + ( Xd_0__inst_mult_1_341  ))
// Xd_0__inst_mult_1_349  = CARRY(( !Xd_0__inst_mult_1_520  $ (((!din_b[16]) # (!din_a[22]))) ) + ( Xd_0__inst_mult_1_342  ) + ( Xd_0__inst_mult_1_341  ))
// Xd_0__inst_mult_1_350  = SHARE((din_b[16] & (din_a[22] & Xd_0__inst_mult_1_520 )))

	.dataa(!din_b[16]),
	.datab(!din_a[22]),
	.datac(!Xd_0__inst_mult_1_520 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_341 ),
	.sharein(Xd_0__inst_mult_1_342 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_348 ),
	.cout(Xd_0__inst_mult_1_349 ),
	.shareout(Xd_0__inst_mult_1_350 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_110 (
// Equation(s):
// Xd_0__inst_mult_1_352  = SUM(( !Xd_0__inst_mult_1_524  $ (!Xd_0__inst_mult_1_528  $ (Xd_0__inst_mult_1_532 )) ) + ( Xd_0__inst_mult_1_346  ) + ( Xd_0__inst_mult_1_345  ))
// Xd_0__inst_mult_1_353  = CARRY(( !Xd_0__inst_mult_1_524  $ (!Xd_0__inst_mult_1_528  $ (Xd_0__inst_mult_1_532 )) ) + ( Xd_0__inst_mult_1_346  ) + ( Xd_0__inst_mult_1_345  ))
// Xd_0__inst_mult_1_354  = SHARE((!Xd_0__inst_mult_1_524  & (Xd_0__inst_mult_1_528  & Xd_0__inst_mult_1_532 )) # (Xd_0__inst_mult_1_524  & ((Xd_0__inst_mult_1_532 ) # (Xd_0__inst_mult_1_528 ))))

	.dataa(!Xd_0__inst_mult_1_524 ),
	.datab(!Xd_0__inst_mult_1_528 ),
	.datac(!Xd_0__inst_mult_1_532 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_345 ),
	.sharein(Xd_0__inst_mult_1_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_352 ),
	.cout(Xd_0__inst_mult_1_353 ),
	.shareout(Xd_0__inst_mult_1_354 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_157 (
// Equation(s):
// Xd_0__inst_mult_6_528  = SUM(( (din_a[81] & din_b[77]) ) + ( Xd_0__inst_mult_6_518  ) + ( Xd_0__inst_mult_6_517  ))
// Xd_0__inst_mult_6_529  = CARRY(( (din_a[81] & din_b[77]) ) + ( Xd_0__inst_mult_6_518  ) + ( Xd_0__inst_mult_6_517  ))
// Xd_0__inst_mult_6_530  = SHARE((din_a[81] & din_b[78]))

	.dataa(!din_a[81]),
	.datab(!din_b[77]),
	.datac(!din_b[78]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_517 ),
	.sharein(Xd_0__inst_mult_6_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_528 ),
	.cout(Xd_0__inst_mult_6_529 ),
	.shareout(Xd_0__inst_mult_6_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_158 (
// Equation(s):
// Xd_0__inst_mult_6_532  = SUM(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_6_522  ) + ( Xd_0__inst_mult_6_521  ))
// Xd_0__inst_mult_6_533  = CARRY(( (din_a[77] & din_b[81]) ) + ( Xd_0__inst_mult_6_522  ) + ( Xd_0__inst_mult_6_521  ))
// Xd_0__inst_mult_6_534  = SHARE((din_a[77] & din_b[82]))

	.dataa(!din_a[77]),
	.datab(!din_b[81]),
	.datac(!din_b[82]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_521 ),
	.sharein(Xd_0__inst_mult_6_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_532 ),
	.cout(Xd_0__inst_mult_6_533 ),
	.shareout(Xd_0__inst_mult_6_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_159 (
// Equation(s):
// Xd_0__inst_mult_6_536  = SUM(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_526  ) + ( Xd_0__inst_mult_6_525  ))
// Xd_0__inst_mult_6_537  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[80])))) # (din_a[79] & (!din_b[79] $ (((!din_a[78]) # (!din_b[80]))))) ) + ( Xd_0__inst_mult_6_526  ) + ( Xd_0__inst_mult_6_525  ))
// Xd_0__inst_mult_6_538  = SHARE((din_a[79] & (din_b[79] & (din_a[78] & din_b[80]))))

	.dataa(!din_a[79]),
	.datab(!din_b[79]),
	.datac(!din_a[78]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_525 ),
	.sharein(Xd_0__inst_mult_6_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_536 ),
	.cout(Xd_0__inst_mult_6_537 ),
	.shareout(Xd_0__inst_mult_6_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_157 (
// Equation(s):
// Xd_0__inst_mult_7_528  = SUM(( (din_a[93] & din_b[89]) ) + ( Xd_0__inst_mult_7_518  ) + ( Xd_0__inst_mult_7_517  ))
// Xd_0__inst_mult_7_529  = CARRY(( (din_a[93] & din_b[89]) ) + ( Xd_0__inst_mult_7_518  ) + ( Xd_0__inst_mult_7_517  ))
// Xd_0__inst_mult_7_530  = SHARE((din_a[93] & din_b[90]))

	.dataa(!din_a[93]),
	.datab(!din_b[89]),
	.datac(!din_b[90]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_517 ),
	.sharein(Xd_0__inst_mult_7_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_528 ),
	.cout(Xd_0__inst_mult_7_529 ),
	.shareout(Xd_0__inst_mult_7_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_158 (
// Equation(s):
// Xd_0__inst_mult_7_532  = SUM(( (din_a[89] & din_b[93]) ) + ( Xd_0__inst_mult_7_522  ) + ( Xd_0__inst_mult_7_521  ))
// Xd_0__inst_mult_7_533  = CARRY(( (din_a[89] & din_b[93]) ) + ( Xd_0__inst_mult_7_522  ) + ( Xd_0__inst_mult_7_521  ))
// Xd_0__inst_mult_7_534  = SHARE((din_a[89] & din_b[94]))

	.dataa(!din_a[89]),
	.datab(!din_b[93]),
	.datac(!din_b[94]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_521 ),
	.sharein(Xd_0__inst_mult_7_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_532 ),
	.cout(Xd_0__inst_mult_7_533 ),
	.shareout(Xd_0__inst_mult_7_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_159 (
// Equation(s):
// Xd_0__inst_mult_7_536  = SUM(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_526  ) + ( Xd_0__inst_mult_7_525  ))
// Xd_0__inst_mult_7_537  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[92])))) # (din_a[91] & (!din_b[91] $ (((!din_a[90]) # (!din_b[92]))))) ) + ( Xd_0__inst_mult_7_526  ) + ( Xd_0__inst_mult_7_525  ))
// Xd_0__inst_mult_7_538  = SHARE((din_a[91] & (din_b[91] & (din_a[90] & din_b[92]))))

	.dataa(!din_a[91]),
	.datab(!din_b[91]),
	.datac(!din_a[90]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_525 ),
	.sharein(Xd_0__inst_mult_7_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_536 ),
	.cout(Xd_0__inst_mult_7_537 ),
	.shareout(Xd_0__inst_mult_7_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_113 (
// Equation(s):
// Xd_0__inst_mult_4_352  = SUM(( GND ) + ( Xd_0__inst_mult_4_346  ) + ( Xd_0__inst_mult_4_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_345 ),
	.sharein(Xd_0__inst_mult_4_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_4_114 (
// Equation(s):
// Xd_0__inst_mult_4_356  = SUM(( !Xd_0__inst_mult_4_544  $ (!Xd_0__inst_mult_4_548  $ (Xd_0__inst_mult_7_572 )) ) + ( Xd_0__inst_mult_4_350  ) + ( Xd_0__inst_mult_4_349  ))
// Xd_0__inst_mult_4_357  = CARRY(( !Xd_0__inst_mult_4_544  $ (!Xd_0__inst_mult_4_548  $ (Xd_0__inst_mult_7_572 )) ) + ( Xd_0__inst_mult_4_350  ) + ( Xd_0__inst_mult_4_349  ))
// Xd_0__inst_mult_4_358  = SHARE((!Xd_0__inst_mult_4_544  & (Xd_0__inst_mult_4_548  & Xd_0__inst_mult_7_572 )) # (Xd_0__inst_mult_4_544  & ((Xd_0__inst_mult_7_572 ) # (Xd_0__inst_mult_4_548 ))))

	.dataa(!Xd_0__inst_mult_4_544 ),
	.datab(!Xd_0__inst_mult_4_548 ),
	.datac(!Xd_0__inst_mult_7_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_349 ),
	.sharein(Xd_0__inst_mult_4_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_356 ),
	.cout(Xd_0__inst_mult_4_357 ),
	.shareout(Xd_0__inst_mult_4_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_113 (
// Equation(s):
// Xd_0__inst_mult_5_352  = SUM(( GND ) + ( Xd_0__inst_mult_5_346  ) + ( Xd_0__inst_mult_5_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_345 ),
	.sharein(Xd_0__inst_mult_5_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_5_114 (
// Equation(s):
// Xd_0__inst_mult_5_356  = SUM(( !Xd_0__inst_mult_5_540  $ (!Xd_0__inst_mult_5_544  $ (Xd_0__inst_mult_5_548 )) ) + ( Xd_0__inst_mult_5_350  ) + ( Xd_0__inst_mult_5_349  ))
// Xd_0__inst_mult_5_357  = CARRY(( !Xd_0__inst_mult_5_540  $ (!Xd_0__inst_mult_5_544  $ (Xd_0__inst_mult_5_548 )) ) + ( Xd_0__inst_mult_5_350  ) + ( Xd_0__inst_mult_5_349  ))
// Xd_0__inst_mult_5_358  = SHARE((!Xd_0__inst_mult_5_540  & (Xd_0__inst_mult_5_544  & Xd_0__inst_mult_5_548 )) # (Xd_0__inst_mult_5_540  & ((Xd_0__inst_mult_5_548 ) # (Xd_0__inst_mult_5_544 ))))

	.dataa(!Xd_0__inst_mult_5_540 ),
	.datab(!Xd_0__inst_mult_5_544 ),
	.datac(!Xd_0__inst_mult_5_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_349 ),
	.sharein(Xd_0__inst_mult_5_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_356 ),
	.cout(Xd_0__inst_mult_5_357 ),
	.shareout(Xd_0__inst_mult_5_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_113 (
// Equation(s):
// Xd_0__inst_mult_2_352  = SUM(( GND ) + ( Xd_0__inst_mult_2_346  ) + ( Xd_0__inst_mult_2_345  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_345 ),
	.sharein(Xd_0__inst_mult_2_346 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_352 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_2_114 (
// Equation(s):
// Xd_0__inst_mult_2_356  = SUM(( !Xd_0__inst_mult_2_540  $ (!Xd_0__inst_mult_2_544  $ (Xd_0__inst_mult_1_536 )) ) + ( Xd_0__inst_mult_2_350  ) + ( Xd_0__inst_mult_2_349  ))
// Xd_0__inst_mult_2_357  = CARRY(( !Xd_0__inst_mult_2_540  $ (!Xd_0__inst_mult_2_544  $ (Xd_0__inst_mult_1_536 )) ) + ( Xd_0__inst_mult_2_350  ) + ( Xd_0__inst_mult_2_349  ))
// Xd_0__inst_mult_2_358  = SHARE((!Xd_0__inst_mult_2_540  & (Xd_0__inst_mult_2_544  & Xd_0__inst_mult_1_536 )) # (Xd_0__inst_mult_2_540  & ((Xd_0__inst_mult_1_536 ) # (Xd_0__inst_mult_2_544 ))))

	.dataa(!Xd_0__inst_mult_2_540 ),
	.datab(!Xd_0__inst_mult_2_544 ),
	.datac(!Xd_0__inst_mult_1_536 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_349 ),
	.sharein(Xd_0__inst_mult_2_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_356 ),
	.cout(Xd_0__inst_mult_2_357 ),
	.shareout(Xd_0__inst_mult_2_358 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_3_118 (
// Equation(s):
// Xd_0__inst_mult_3_384  = SUM(( !Xd_0__inst_mult_3_556  $ (!Xd_0__inst_mult_3_272  $ (Xd_0__inst_mult_2_548 )) ) + ( Xd_0__inst_mult_3_382  ) + ( Xd_0__inst_mult_3_381  ))
// Xd_0__inst_mult_3_385  = CARRY(( !Xd_0__inst_mult_3_556  $ (!Xd_0__inst_mult_3_272  $ (Xd_0__inst_mult_2_548 )) ) + ( Xd_0__inst_mult_3_382  ) + ( Xd_0__inst_mult_3_381  ))
// Xd_0__inst_mult_3_386  = SHARE((!Xd_0__inst_mult_3_556  & (Xd_0__inst_mult_3_272  & Xd_0__inst_mult_2_548 )) # (Xd_0__inst_mult_3_556  & ((Xd_0__inst_mult_2_548 ) # (Xd_0__inst_mult_3_272 ))))

	.dataa(!Xd_0__inst_mult_3_556 ),
	.datab(!Xd_0__inst_mult_3_272 ),
	.datac(!Xd_0__inst_mult_2_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_381 ),
	.sharein(Xd_0__inst_mult_3_382 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_384 ),
	.cout(Xd_0__inst_mult_3_385 ),
	.shareout(Xd_0__inst_mult_3_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_0_112 (
// Equation(s):
// Xd_0__inst_mult_0_360  = SUM(( !Xd_0__inst_mult_0_536  $ (!Xd_0__inst_mult_0_540  $ (Xd_0__inst_mult_0_544 )) ) + ( Xd_0__inst_mult_0_358  ) + ( Xd_0__inst_mult_0_357  ))
// Xd_0__inst_mult_0_361  = CARRY(( !Xd_0__inst_mult_0_536  $ (!Xd_0__inst_mult_0_540  $ (Xd_0__inst_mult_0_544 )) ) + ( Xd_0__inst_mult_0_358  ) + ( Xd_0__inst_mult_0_357  ))
// Xd_0__inst_mult_0_362  = SHARE((!Xd_0__inst_mult_0_536  & (Xd_0__inst_mult_0_540  & Xd_0__inst_mult_0_544 )) # (Xd_0__inst_mult_0_536  & ((Xd_0__inst_mult_0_544 ) # (Xd_0__inst_mult_0_540 ))))

	.dataa(!Xd_0__inst_mult_0_536 ),
	.datab(!Xd_0__inst_mult_0_540 ),
	.datac(!Xd_0__inst_mult_0_544 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_357 ),
	.sharein(Xd_0__inst_mult_0_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_360 ),
	.cout(Xd_0__inst_mult_0_361 ),
	.shareout(Xd_0__inst_mult_0_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_111 (
// Equation(s):
// Xd_0__inst_mult_1_356  = SUM(( GND ) + ( Xd_0__inst_mult_1_350  ) + ( Xd_0__inst_mult_1_349  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_349 ),
	.sharein(Xd_0__inst_mult_1_350 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_356 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000171700006969),
	.shared_arith("on")
) Xd_0__inst_mult_1_112 (
// Equation(s):
// Xd_0__inst_mult_1_360  = SUM(( !Xd_0__inst_mult_1_540  $ (!Xd_0__inst_mult_1_544  $ (Xd_0__inst_mult_1_548 )) ) + ( Xd_0__inst_mult_1_354  ) + ( Xd_0__inst_mult_1_353  ))
// Xd_0__inst_mult_1_361  = CARRY(( !Xd_0__inst_mult_1_540  $ (!Xd_0__inst_mult_1_544  $ (Xd_0__inst_mult_1_548 )) ) + ( Xd_0__inst_mult_1_354  ) + ( Xd_0__inst_mult_1_353  ))
// Xd_0__inst_mult_1_362  = SHARE((!Xd_0__inst_mult_1_540  & (Xd_0__inst_mult_1_544  & Xd_0__inst_mult_1_548 )) # (Xd_0__inst_mult_1_540  & ((Xd_0__inst_mult_1_548 ) # (Xd_0__inst_mult_1_544 ))))

	.dataa(!Xd_0__inst_mult_1_540 ),
	.datab(!Xd_0__inst_mult_1_544 ),
	.datac(!Xd_0__inst_mult_1_548 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_353 ),
	.sharein(Xd_0__inst_mult_1_354 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_360 ),
	.cout(Xd_0__inst_mult_1_361 ),
	.shareout(Xd_0__inst_mult_1_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_160 (
// Equation(s):
// Xd_0__inst_mult_6_540  = SUM(( (din_a[80] & din_b[79]) ) + ( Xd_0__inst_mult_6_530  ) + ( Xd_0__inst_mult_6_529  ))
// Xd_0__inst_mult_6_541  = CARRY(( (din_a[80] & din_b[79]) ) + ( Xd_0__inst_mult_6_530  ) + ( Xd_0__inst_mult_6_529  ))
// Xd_0__inst_mult_6_542  = SHARE((din_b[79] & din_a[81]))

	.dataa(!din_a[80]),
	.datab(!din_b[79]),
	.datac(!din_a[81]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_529 ),
	.sharein(Xd_0__inst_mult_6_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_540 ),
	.cout(Xd_0__inst_mult_6_541 ),
	.shareout(Xd_0__inst_mult_6_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_161 (
// Equation(s):
// Xd_0__inst_mult_6_544  = SUM(( (!din_a[79] & (((din_a[78] & din_b[81])))) # (din_a[79] & (!din_b[80] $ (((!din_a[78]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_6_534  ) + ( Xd_0__inst_mult_6_533  ))
// Xd_0__inst_mult_6_545  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[81])))) # (din_a[79] & (!din_b[80] $ (((!din_a[78]) # (!din_b[81]))))) ) + ( Xd_0__inst_mult_6_534  ) + ( Xd_0__inst_mult_6_533  ))
// Xd_0__inst_mult_6_546  = SHARE((din_a[79] & (din_b[80] & (din_a[78] & din_b[81]))))

	.dataa(!din_a[79]),
	.datab(!din_b[80]),
	.datac(!din_a[78]),
	.datad(!din_b[81]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_533 ),
	.sharein(Xd_0__inst_mult_6_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_544 ),
	.cout(Xd_0__inst_mult_6_545 ),
	.shareout(Xd_0__inst_mult_6_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_162 (
// Equation(s):
// Xd_0__inst_mult_6_548  = SUM(( GND ) + ( Xd_0__inst_mult_6_538  ) + ( Xd_0__inst_mult_6_537  ))
// Xd_0__inst_mult_6_549  = CARRY(( GND ) + ( Xd_0__inst_mult_6_538  ) + ( Xd_0__inst_mult_6_537  ))
// Xd_0__inst_mult_6_550  = SHARE(VCC)

	.dataa(!din_a[75]),
	.datab(!din_b[73]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_537 ),
	.sharein(Xd_0__inst_mult_6_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_548 ),
	.cout(Xd_0__inst_mult_6_549 ),
	.shareout(Xd_0__inst_mult_6_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_160 (
// Equation(s):
// Xd_0__inst_mult_7_540  = SUM(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_7_530  ) + ( Xd_0__inst_mult_7_529  ))
// Xd_0__inst_mult_7_541  = CARRY(( (din_a[92] & din_b[91]) ) + ( Xd_0__inst_mult_7_530  ) + ( Xd_0__inst_mult_7_529  ))
// Xd_0__inst_mult_7_542  = SHARE((din_b[91] & din_a[93]))

	.dataa(!din_a[92]),
	.datab(!din_b[91]),
	.datac(!din_a[93]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_529 ),
	.sharein(Xd_0__inst_mult_7_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_540 ),
	.cout(Xd_0__inst_mult_7_541 ),
	.shareout(Xd_0__inst_mult_7_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_161 (
// Equation(s):
// Xd_0__inst_mult_7_544  = SUM(( (!din_a[91] & (((din_a[90] & din_b[93])))) # (din_a[91] & (!din_b[92] $ (((!din_a[90]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_7_534  ) + ( Xd_0__inst_mult_7_533  ))
// Xd_0__inst_mult_7_545  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[93])))) # (din_a[91] & (!din_b[92] $ (((!din_a[90]) # (!din_b[93]))))) ) + ( Xd_0__inst_mult_7_534  ) + ( Xd_0__inst_mult_7_533  ))
// Xd_0__inst_mult_7_546  = SHARE((din_a[91] & (din_b[92] & (din_a[90] & din_b[93]))))

	.dataa(!din_a[91]),
	.datab(!din_b[92]),
	.datac(!din_a[90]),
	.datad(!din_b[93]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_533 ),
	.sharein(Xd_0__inst_mult_7_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_544 ),
	.cout(Xd_0__inst_mult_7_545 ),
	.shareout(Xd_0__inst_mult_7_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_115 (
// Equation(s):
// Xd_0__inst_mult_4_360  = SUM(( GND ) + ( Xd_0__inst_mult_7_538  ) + ( Xd_0__inst_mult_7_537  ))
// Xd_0__inst_mult_4_361  = CARRY(( GND ) + ( Xd_0__inst_mult_7_538  ) + ( Xd_0__inst_mult_7_537  ))
// Xd_0__inst_mult_4_362  = SHARE(VCC)

	.dataa(!din_a[50]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_537 ),
	.sharein(Xd_0__inst_mult_7_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_360 ),
	.cout(Xd_0__inst_mult_4_361 ),
	.shareout(Xd_0__inst_mult_4_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_4_116 (
// Equation(s):
// Xd_0__inst_mult_4_364  = SUM(( !Xd_0__inst_mult_4_552  $ (!Xd_0__inst_mult_4_556 ) ) + ( Xd_0__inst_mult_4_358  ) + ( Xd_0__inst_mult_4_357  ))
// Xd_0__inst_mult_4_365  = CARRY(( !Xd_0__inst_mult_4_552  $ (!Xd_0__inst_mult_4_556 ) ) + ( Xd_0__inst_mult_4_358  ) + ( Xd_0__inst_mult_4_357  ))
// Xd_0__inst_mult_4_366  = SHARE((Xd_0__inst_mult_4_552  & Xd_0__inst_mult_4_556 ))

	.dataa(!Xd_0__inst_mult_4_552 ),
	.datab(!Xd_0__inst_mult_4_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_357 ),
	.sharein(Xd_0__inst_mult_4_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_364 ),
	.cout(Xd_0__inst_mult_4_365 ),
	.shareout(Xd_0__inst_mult_4_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_39 (
// Equation(s):
// Xd_0__inst_mult_4_39_sumout  = SUM(( (din_a[58] & din_b[54]) ) + ( Xd_0__inst_mult_7_69  ) + ( Xd_0__inst_mult_7_68  ))
// Xd_0__inst_mult_4_40  = CARRY(( (din_a[58] & din_b[54]) ) + ( Xd_0__inst_mult_7_69  ) + ( Xd_0__inst_mult_7_68  ))
// Xd_0__inst_mult_4_41  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_68 ),
	.sharein(Xd_0__inst_mult_7_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_39_sumout ),
	.cout(Xd_0__inst_mult_4_40 ),
	.shareout(Xd_0__inst_mult_4_41 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_5_115 (
// Equation(s):
// Xd_0__inst_mult_5_360  = SUM(( !Xd_0__inst_mult_5_552  $ (!Xd_0__inst_mult_5_556 ) ) + ( Xd_0__inst_mult_5_358  ) + ( Xd_0__inst_mult_5_357  ))
// Xd_0__inst_mult_5_361  = CARRY(( !Xd_0__inst_mult_5_552  $ (!Xd_0__inst_mult_5_556 ) ) + ( Xd_0__inst_mult_5_358  ) + ( Xd_0__inst_mult_5_357  ))
// Xd_0__inst_mult_5_362  = SHARE((Xd_0__inst_mult_5_552  & Xd_0__inst_mult_5_556 ))

	.dataa(!Xd_0__inst_mult_5_552 ),
	.datab(!Xd_0__inst_mult_5_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_357 ),
	.sharein(Xd_0__inst_mult_5_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_360 ),
	.cout(Xd_0__inst_mult_5_361 ),
	.shareout(Xd_0__inst_mult_5_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_51 (
// Equation(s):
// Xd_0__inst_mult_5_51_sumout  = SUM(( (din_a[70] & din_b[66]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_52  = CARRY(( (din_a[70] & din_b[66]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_53  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_51_sumout ),
	.cout(Xd_0__inst_mult_5_52 ),
	.shareout(Xd_0__inst_mult_5_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_2_115 (
// Equation(s):
// Xd_0__inst_mult_2_360  = SUM(( !Xd_0__inst_mult_2_552  $ (!Xd_0__inst_mult_2_556 ) ) + ( Xd_0__inst_mult_2_358  ) + ( Xd_0__inst_mult_2_357  ))
// Xd_0__inst_mult_2_361  = CARRY(( !Xd_0__inst_mult_2_552  $ (!Xd_0__inst_mult_2_556 ) ) + ( Xd_0__inst_mult_2_358  ) + ( Xd_0__inst_mult_2_357  ))
// Xd_0__inst_mult_2_362  = SHARE((Xd_0__inst_mult_2_552  & Xd_0__inst_mult_2_556 ))

	.dataa(!Xd_0__inst_mult_2_552 ),
	.datab(!Xd_0__inst_mult_2_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_357 ),
	.sharein(Xd_0__inst_mult_2_358 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_360 ),
	.cout(Xd_0__inst_mult_2_361 ),
	.shareout(Xd_0__inst_mult_2_362 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_51 (
// Equation(s):
// Xd_0__inst_mult_2_51_sumout  = SUM(( (din_a[34] & din_b[30]) ) + ( Xd_0__inst_mult_5_53  ) + ( Xd_0__inst_mult_5_52  ))
// Xd_0__inst_mult_2_52  = CARRY(( (din_a[34] & din_b[30]) ) + ( Xd_0__inst_mult_5_53  ) + ( Xd_0__inst_mult_5_52  ))
// Xd_0__inst_mult_2_53  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_52 ),
	.sharein(Xd_0__inst_mult_5_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_51_sumout ),
	.cout(Xd_0__inst_mult_2_52 ),
	.shareout(Xd_0__inst_mult_2_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_3_119 (
// Equation(s):
// Xd_0__inst_mult_3_388  = SUM(( !Xd_0__inst_mult_3_560  $ (!Xd_0__inst_mult_3_188 ) ) + ( Xd_0__inst_mult_3_386  ) + ( Xd_0__inst_mult_3_385  ))
// Xd_0__inst_mult_3_389  = CARRY(( !Xd_0__inst_mult_3_560  $ (!Xd_0__inst_mult_3_188 ) ) + ( Xd_0__inst_mult_3_386  ) + ( Xd_0__inst_mult_3_385  ))
// Xd_0__inst_mult_3_390  = SHARE((Xd_0__inst_mult_3_560  & Xd_0__inst_mult_3_188 ))

	.dataa(!Xd_0__inst_mult_3_560 ),
	.datab(!Xd_0__inst_mult_3_188 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_385 ),
	.sharein(Xd_0__inst_mult_3_386 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_388 ),
	.cout(Xd_0__inst_mult_3_389 ),
	.shareout(Xd_0__inst_mult_3_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_0_113 (
// Equation(s):
// Xd_0__inst_mult_0_364  = SUM(( !Xd_0__inst_mult_0_548  $ (!Xd_0__inst_mult_0_552 ) ) + ( Xd_0__inst_mult_0_362  ) + ( Xd_0__inst_mult_0_361  ))
// Xd_0__inst_mult_0_365  = CARRY(( !Xd_0__inst_mult_0_548  $ (!Xd_0__inst_mult_0_552 ) ) + ( Xd_0__inst_mult_0_362  ) + ( Xd_0__inst_mult_0_361  ))
// Xd_0__inst_mult_0_366  = SHARE((Xd_0__inst_mult_0_548  & Xd_0__inst_mult_0_552 ))

	.dataa(!Xd_0__inst_mult_0_548 ),
	.datab(!Xd_0__inst_mult_0_552 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_361 ),
	.sharein(Xd_0__inst_mult_0_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_364 ),
	.cout(Xd_0__inst_mult_0_365 ),
	.shareout(Xd_0__inst_mult_0_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_51 (
// Equation(s):
// Xd_0__inst_mult_0_51_sumout  = SUM(( (din_a[10] & din_b[6]) ) + ( Xd_0__inst_mult_5_61  ) + ( Xd_0__inst_mult_5_60  ))
// Xd_0__inst_mult_0_52  = CARRY(( (din_a[10] & din_b[6]) ) + ( Xd_0__inst_mult_5_61  ) + ( Xd_0__inst_mult_5_60  ))
// Xd_0__inst_mult_0_53  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_60 ),
	.sharein(Xd_0__inst_mult_5_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_51_sumout ),
	.cout(Xd_0__inst_mult_0_52 ),
	.shareout(Xd_0__inst_mult_0_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100006666),
	.shared_arith("on")
) Xd_0__inst_mult_1_113 (
// Equation(s):
// Xd_0__inst_mult_1_364  = SUM(( !Xd_0__inst_mult_1_552  $ (!Xd_0__inst_mult_1_556 ) ) + ( Xd_0__inst_mult_1_362  ) + ( Xd_0__inst_mult_1_361  ))
// Xd_0__inst_mult_1_365  = CARRY(( !Xd_0__inst_mult_1_552  $ (!Xd_0__inst_mult_1_556 ) ) + ( Xd_0__inst_mult_1_362  ) + ( Xd_0__inst_mult_1_361  ))
// Xd_0__inst_mult_1_366  = SHARE((Xd_0__inst_mult_1_552  & Xd_0__inst_mult_1_556 ))

	.dataa(!Xd_0__inst_mult_1_552 ),
	.datab(!Xd_0__inst_mult_1_556 ),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_361 ),
	.sharein(Xd_0__inst_mult_1_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_364 ),
	.cout(Xd_0__inst_mult_1_365 ),
	.shareout(Xd_0__inst_mult_1_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_51 (
// Equation(s):
// Xd_0__inst_mult_1_51_sumout  = SUM(( (din_a[22] & din_b[18]) ) + ( Xd_0__inst_mult_0_53  ) + ( Xd_0__inst_mult_0_52  ))
// Xd_0__inst_mult_1_52  = CARRY(( (din_a[22] & din_b[18]) ) + ( Xd_0__inst_mult_0_53  ) + ( Xd_0__inst_mult_0_52  ))
// Xd_0__inst_mult_1_53  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_52 ),
	.sharein(Xd_0__inst_mult_0_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_51_sumout ),
	.cout(Xd_0__inst_mult_1_52 ),
	.shareout(Xd_0__inst_mult_1_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_163 (
// Equation(s):
// Xd_0__inst_mult_6_552  = SUM(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_6_542  ) + ( Xd_0__inst_mult_6_541  ))
// Xd_0__inst_mult_6_553  = CARRY(( (din_a[80] & din_b[80]) ) + ( Xd_0__inst_mult_6_542  ) + ( Xd_0__inst_mult_6_541  ))
// Xd_0__inst_mult_6_554  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[80]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_541 ),
	.sharein(Xd_0__inst_mult_6_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_552 ),
	.cout(Xd_0__inst_mult_6_553 ),
	.shareout(Xd_0__inst_mult_6_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_164 (
// Equation(s):
// Xd_0__inst_mult_6_556  = SUM(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_546  ) + ( Xd_0__inst_mult_6_545  ))
// Xd_0__inst_mult_6_557  = CARRY(( (!din_a[79] & (((din_a[78] & din_b[82])))) # (din_a[79] & (!din_b[81] $ (((!din_a[78]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_546  ) + ( Xd_0__inst_mult_6_545  ))
// Xd_0__inst_mult_6_558  = SHARE((din_a[79] & (din_b[81] & (din_a[78] & din_b[82]))))

	.dataa(!din_a[79]),
	.datab(!din_b[81]),
	.datac(!din_a[78]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_545 ),
	.sharein(Xd_0__inst_mult_6_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_556 ),
	.cout(Xd_0__inst_mult_6_557 ),
	.shareout(Xd_0__inst_mult_6_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_162 (
// Equation(s):
// Xd_0__inst_mult_7_548  = SUM(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_7_542  ) + ( Xd_0__inst_mult_7_541  ))
// Xd_0__inst_mult_7_549  = CARRY(( (din_a[92] & din_b[92]) ) + ( Xd_0__inst_mult_7_542  ) + ( Xd_0__inst_mult_7_541  ))
// Xd_0__inst_mult_7_550  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[92]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_541 ),
	.sharein(Xd_0__inst_mult_7_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_548 ),
	.cout(Xd_0__inst_mult_7_549 ),
	.shareout(Xd_0__inst_mult_7_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_163 (
// Equation(s):
// Xd_0__inst_mult_7_552  = SUM(( (!din_a[91] & (((din_a[90] & din_b[94])))) # (din_a[91] & (!din_b[93] $ (((!din_a[90]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_546  ) + ( Xd_0__inst_mult_7_545  ))
// Xd_0__inst_mult_7_553  = CARRY(( (!din_a[91] & (((din_a[90] & din_b[94])))) # (din_a[91] & (!din_b[93] $ (((!din_a[90]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_546  ) + ( Xd_0__inst_mult_7_545  ))
// Xd_0__inst_mult_7_554  = SHARE((din_a[91] & (din_b[93] & (din_a[90] & din_b[94]))))

	.dataa(!din_a[91]),
	.datab(!din_b[93]),
	.datac(!din_a[90]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_545 ),
	.sharein(Xd_0__inst_mult_7_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_552 ),
	.cout(Xd_0__inst_mult_7_553 ),
	.shareout(Xd_0__inst_mult_7_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_4_117 (
// Equation(s):
// Xd_0__inst_mult_4_368  = SUM(( !Xd_0__inst_mult_4_560  $ (!Xd_0__inst_mult_4_564  $ (((din_a[57] & din_b[56])))) ) + ( Xd_0__inst_mult_4_366  ) + ( Xd_0__inst_mult_4_365  ))
// Xd_0__inst_mult_4_369  = CARRY(( !Xd_0__inst_mult_4_560  $ (!Xd_0__inst_mult_4_564  $ (((din_a[57] & din_b[56])))) ) + ( Xd_0__inst_mult_4_366  ) + ( Xd_0__inst_mult_4_365  ))
// Xd_0__inst_mult_4_370  = SHARE((!Xd_0__inst_mult_4_560  & (Xd_0__inst_mult_4_564  & (din_a[57] & din_b[56]))) # (Xd_0__inst_mult_4_560  & (((din_a[57] & din_b[56])) # (Xd_0__inst_mult_4_564 ))))

	.dataa(!Xd_0__inst_mult_4_560 ),
	.datab(!Xd_0__inst_mult_4_564 ),
	.datac(!din_a[57]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_365 ),
	.sharein(Xd_0__inst_mult_4_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_368 ),
	.cout(Xd_0__inst_mult_4_369 ),
	.shareout(Xd_0__inst_mult_4_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_43 (
// Equation(s):
// Xd_0__inst_mult_4_43_sumout  = SUM(( (din_a[58] & din_b[55]) ) + ( Xd_0__inst_mult_1_53  ) + ( Xd_0__inst_mult_1_52  ))
// Xd_0__inst_mult_4_44  = CARRY(( (din_a[58] & din_b[55]) ) + ( Xd_0__inst_mult_1_53  ) + ( Xd_0__inst_mult_1_52  ))
// Xd_0__inst_mult_4_45  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[55]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_52 ),
	.sharein(Xd_0__inst_mult_1_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_43_sumout ),
	.cout(Xd_0__inst_mult_4_44 ),
	.shareout(Xd_0__inst_mult_4_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_5_116 (
// Equation(s):
// Xd_0__inst_mult_5_364  = SUM(( !Xd_0__inst_mult_5_560  $ (!Xd_0__inst_mult_5_564  $ (((din_a[69] & din_b[68])))) ) + ( Xd_0__inst_mult_5_362  ) + ( Xd_0__inst_mult_5_361  ))
// Xd_0__inst_mult_5_365  = CARRY(( !Xd_0__inst_mult_5_560  $ (!Xd_0__inst_mult_5_564  $ (((din_a[69] & din_b[68])))) ) + ( Xd_0__inst_mult_5_362  ) + ( Xd_0__inst_mult_5_361  ))
// Xd_0__inst_mult_5_366  = SHARE((!Xd_0__inst_mult_5_560  & (Xd_0__inst_mult_5_564  & (din_a[69] & din_b[68]))) # (Xd_0__inst_mult_5_560  & (((din_a[69] & din_b[68])) # (Xd_0__inst_mult_5_564 ))))

	.dataa(!Xd_0__inst_mult_5_560 ),
	.datab(!Xd_0__inst_mult_5_564 ),
	.datac(!din_a[69]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_361 ),
	.sharein(Xd_0__inst_mult_5_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_364 ),
	.cout(Xd_0__inst_mult_5_365 ),
	.shareout(Xd_0__inst_mult_5_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_55 (
// Equation(s):
// Xd_0__inst_mult_5_55_sumout  = SUM(( (din_a[70] & din_b[67]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_56  = CARRY(( (din_a[70] & din_b[67]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_57  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_55_sumout ),
	.cout(Xd_0__inst_mult_5_56 ),
	.shareout(Xd_0__inst_mult_5_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_2_116 (
// Equation(s):
// Xd_0__inst_mult_2_364  = SUM(( !Xd_0__inst_mult_2_560  $ (!Xd_0__inst_mult_2_564  $ (((din_a[33] & din_b[32])))) ) + ( Xd_0__inst_mult_2_362  ) + ( Xd_0__inst_mult_2_361  ))
// Xd_0__inst_mult_2_365  = CARRY(( !Xd_0__inst_mult_2_560  $ (!Xd_0__inst_mult_2_564  $ (((din_a[33] & din_b[32])))) ) + ( Xd_0__inst_mult_2_362  ) + ( Xd_0__inst_mult_2_361  ))
// Xd_0__inst_mult_2_366  = SHARE((!Xd_0__inst_mult_2_560  & (Xd_0__inst_mult_2_564  & (din_a[33] & din_b[32]))) # (Xd_0__inst_mult_2_560  & (((din_a[33] & din_b[32])) # (Xd_0__inst_mult_2_564 ))))

	.dataa(!Xd_0__inst_mult_2_560 ),
	.datab(!Xd_0__inst_mult_2_564 ),
	.datac(!din_a[33]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_361 ),
	.sharein(Xd_0__inst_mult_2_362 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_364 ),
	.cout(Xd_0__inst_mult_2_365 ),
	.shareout(Xd_0__inst_mult_2_366 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_55 (
// Equation(s):
// Xd_0__inst_mult_2_55_sumout  = SUM(( (din_a[34] & din_b[31]) ) + ( Xd_0__inst_mult_5_57  ) + ( Xd_0__inst_mult_5_56  ))
// Xd_0__inst_mult_2_56  = CARRY(( (din_a[34] & din_b[31]) ) + ( Xd_0__inst_mult_5_57  ) + ( Xd_0__inst_mult_5_56  ))
// Xd_0__inst_mult_2_57  = SHARE(GND)

	.dataa(!din_a[34]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_56 ),
	.sharein(Xd_0__inst_mult_5_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_55_sumout ),
	.cout(Xd_0__inst_mult_2_56 ),
	.shareout(Xd_0__inst_mult_2_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_3_120 (
// Equation(s):
// Xd_0__inst_mult_3_392  = SUM(( !Xd_0__inst_mult_3_564  $ (!Xd_0__inst_mult_3_180  $ (((din_a[45] & din_b[44])))) ) + ( Xd_0__inst_mult_3_390  ) + ( Xd_0__inst_mult_3_389  ))
// Xd_0__inst_mult_3_393  = CARRY(( !Xd_0__inst_mult_3_564  $ (!Xd_0__inst_mult_3_180  $ (((din_a[45] & din_b[44])))) ) + ( Xd_0__inst_mult_3_390  ) + ( Xd_0__inst_mult_3_389  ))
// Xd_0__inst_mult_3_394  = SHARE((!Xd_0__inst_mult_3_564  & (Xd_0__inst_mult_3_180  & (din_a[45] & din_b[44]))) # (Xd_0__inst_mult_3_564  & (((din_a[45] & din_b[44])) # (Xd_0__inst_mult_3_180 ))))

	.dataa(!Xd_0__inst_mult_3_564 ),
	.datab(!Xd_0__inst_mult_3_180 ),
	.datac(!din_a[45]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_389 ),
	.sharein(Xd_0__inst_mult_3_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_392 ),
	.cout(Xd_0__inst_mult_3_393 ),
	.shareout(Xd_0__inst_mult_3_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_43 (
// Equation(s):
// Xd_0__inst_mult_3_43_sumout  = SUM(( (din_a[46] & din_b[43]) ) + ( Xd_0__inst_mult_2_57  ) + ( Xd_0__inst_mult_2_56  ))
// Xd_0__inst_mult_3_44  = CARRY(( (din_a[46] & din_b[43]) ) + ( Xd_0__inst_mult_2_57  ) + ( Xd_0__inst_mult_2_56  ))
// Xd_0__inst_mult_3_45  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_56 ),
	.sharein(Xd_0__inst_mult_2_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_43_sumout ),
	.cout(Xd_0__inst_mult_3_44 ),
	.shareout(Xd_0__inst_mult_3_45 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_0_114 (
// Equation(s):
// Xd_0__inst_mult_0_368  = SUM(( !Xd_0__inst_mult_0_556  $ (!Xd_0__inst_mult_0_560  $ (((din_a[9] & din_b[8])))) ) + ( Xd_0__inst_mult_0_366  ) + ( Xd_0__inst_mult_0_365  ))
// Xd_0__inst_mult_0_369  = CARRY(( !Xd_0__inst_mult_0_556  $ (!Xd_0__inst_mult_0_560  $ (((din_a[9] & din_b[8])))) ) + ( Xd_0__inst_mult_0_366  ) + ( Xd_0__inst_mult_0_365  ))
// Xd_0__inst_mult_0_370  = SHARE((!Xd_0__inst_mult_0_556  & (Xd_0__inst_mult_0_560  & (din_a[9] & din_b[8]))) # (Xd_0__inst_mult_0_556  & (((din_a[9] & din_b[8])) # (Xd_0__inst_mult_0_560 ))))

	.dataa(!Xd_0__inst_mult_0_556 ),
	.datab(!Xd_0__inst_mult_0_560 ),
	.datac(!din_a[9]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_365 ),
	.sharein(Xd_0__inst_mult_0_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_368 ),
	.cout(Xd_0__inst_mult_0_369 ),
	.shareout(Xd_0__inst_mult_0_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_55 (
// Equation(s):
// Xd_0__inst_mult_0_55_sumout  = SUM(( (din_a[10] & din_b[7]) ) + ( Xd_0__inst_mult_3_45  ) + ( Xd_0__inst_mult_3_44  ))
// Xd_0__inst_mult_0_56  = CARRY(( (din_a[10] & din_b[7]) ) + ( Xd_0__inst_mult_3_45  ) + ( Xd_0__inst_mult_3_44  ))
// Xd_0__inst_mult_0_57  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_44 ),
	.sharein(Xd_0__inst_mult_3_45 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_55_sumout ),
	.cout(Xd_0__inst_mult_0_56 ),
	.shareout(Xd_0__inst_mult_0_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111700006669),
	.shared_arith("on")
) Xd_0__inst_mult_1_114 (
// Equation(s):
// Xd_0__inst_mult_1_368  = SUM(( !Xd_0__inst_mult_1_560  $ (!Xd_0__inst_mult_1_564  $ (((din_a[21] & din_b[20])))) ) + ( Xd_0__inst_mult_1_366  ) + ( Xd_0__inst_mult_1_365  ))
// Xd_0__inst_mult_1_369  = CARRY(( !Xd_0__inst_mult_1_560  $ (!Xd_0__inst_mult_1_564  $ (((din_a[21] & din_b[20])))) ) + ( Xd_0__inst_mult_1_366  ) + ( Xd_0__inst_mult_1_365  ))
// Xd_0__inst_mult_1_370  = SHARE((!Xd_0__inst_mult_1_560  & (Xd_0__inst_mult_1_564  & (din_a[21] & din_b[20]))) # (Xd_0__inst_mult_1_560  & (((din_a[21] & din_b[20])) # (Xd_0__inst_mult_1_564 ))))

	.dataa(!Xd_0__inst_mult_1_560 ),
	.datab(!Xd_0__inst_mult_1_564 ),
	.datac(!din_a[21]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_365 ),
	.sharein(Xd_0__inst_mult_1_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_368 ),
	.cout(Xd_0__inst_mult_1_369 ),
	.shareout(Xd_0__inst_mult_1_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_55 (
// Equation(s):
// Xd_0__inst_mult_1_55_sumout  = SUM(( (din_a[22] & din_b[19]) ) + ( Xd_0__inst_mult_0_57  ) + ( Xd_0__inst_mult_0_56  ))
// Xd_0__inst_mult_1_56  = CARRY(( (din_a[22] & din_b[19]) ) + ( Xd_0__inst_mult_0_57  ) + ( Xd_0__inst_mult_0_56  ))
// Xd_0__inst_mult_1_57  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_56 ),
	.sharein(Xd_0__inst_mult_0_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_55_sumout ),
	.cout(Xd_0__inst_mult_1_56 ),
	.shareout(Xd_0__inst_mult_1_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_165 (
// Equation(s):
// Xd_0__inst_mult_6_560  = SUM(( GND ) + ( Xd_0__inst_mult_6_554  ) + ( Xd_0__inst_mult_6_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_553 ),
	.sharein(Xd_0__inst_mult_6_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_6_166 (
// Equation(s):
// Xd_0__inst_mult_6_564  = SUM(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_558  ) + ( Xd_0__inst_mult_6_557  ))
// Xd_0__inst_mult_6_565  = CARRY(( (!din_a[80] & (((din_a[79] & din_b[82])))) # (din_a[80] & (!din_b[81] $ (((!din_a[79]) # (!din_b[82]))))) ) + ( Xd_0__inst_mult_6_558  ) + ( Xd_0__inst_mult_6_557  ))
// Xd_0__inst_mult_6_566  = SHARE((din_a[80] & (din_b[81] & (din_a[79] & din_b[82]))))

	.dataa(!din_a[80]),
	.datab(!din_b[81]),
	.datac(!din_a[79]),
	.datad(!din_b[82]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_557 ),
	.sharein(Xd_0__inst_mult_6_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_564 ),
	.cout(Xd_0__inst_mult_6_565 ),
	.shareout(Xd_0__inst_mult_6_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_164 (
// Equation(s):
// Xd_0__inst_mult_7_556  = SUM(( GND ) + ( Xd_0__inst_mult_7_550  ) + ( Xd_0__inst_mult_7_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_549 ),
	.sharein(Xd_0__inst_mult_7_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_7_165 (
// Equation(s):
// Xd_0__inst_mult_7_560  = SUM(( (!din_a[92] & (((din_a[91] & din_b[94])))) # (din_a[92] & (!din_b[93] $ (((!din_a[91]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_554  ) + ( Xd_0__inst_mult_7_553  ))
// Xd_0__inst_mult_7_561  = CARRY(( (!din_a[92] & (((din_a[91] & din_b[94])))) # (din_a[92] & (!din_b[93] $ (((!din_a[91]) # (!din_b[94]))))) ) + ( Xd_0__inst_mult_7_554  ) + ( Xd_0__inst_mult_7_553  ))
// Xd_0__inst_mult_7_562  = SHARE((din_a[92] & (din_b[93] & (din_a[91] & din_b[94]))))

	.dataa(!din_a[92]),
	.datab(!din_b[93]),
	.datac(!din_a[91]),
	.datad(!din_b[94]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_553 ),
	.sharein(Xd_0__inst_mult_7_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_560 ),
	.cout(Xd_0__inst_mult_7_561 ),
	.shareout(Xd_0__inst_mult_7_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_118 (
// Equation(s):
// Xd_0__inst_mult_4_372  = SUM(( !Xd_0__inst_mult_4_568  $ (((!din_a[57]) # (!din_b[57]))) ) + ( Xd_0__inst_mult_4_370  ) + ( Xd_0__inst_mult_4_369  ))
// Xd_0__inst_mult_4_373  = CARRY(( !Xd_0__inst_mult_4_568  $ (((!din_a[57]) # (!din_b[57]))) ) + ( Xd_0__inst_mult_4_370  ) + ( Xd_0__inst_mult_4_369  ))
// Xd_0__inst_mult_4_374  = SHARE((din_a[57] & (din_b[57] & Xd_0__inst_mult_4_568 )))

	.dataa(!din_a[57]),
	.datab(!din_b[57]),
	.datac(!Xd_0__inst_mult_4_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_369 ),
	.sharein(Xd_0__inst_mult_4_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_372 ),
	.cout(Xd_0__inst_mult_4_373 ),
	.shareout(Xd_0__inst_mult_4_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_47 (
// Equation(s):
// Xd_0__inst_mult_4_47_sumout  = SUM(( (din_a[58] & din_b[56]) ) + ( Xd_0__inst_mult_1_57  ) + ( Xd_0__inst_mult_1_56  ))
// Xd_0__inst_mult_4_48  = CARRY(( (din_a[58] & din_b[56]) ) + ( Xd_0__inst_mult_1_57  ) + ( Xd_0__inst_mult_1_56  ))
// Xd_0__inst_mult_4_49  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_56 ),
	.sharein(Xd_0__inst_mult_1_57 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_47_sumout ),
	.cout(Xd_0__inst_mult_4_48 ),
	.shareout(Xd_0__inst_mult_4_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_117 (
// Equation(s):
// Xd_0__inst_mult_5_368  = SUM(( !Xd_0__inst_mult_5_568  $ (((!din_a[69]) # (!din_b[69]))) ) + ( Xd_0__inst_mult_5_366  ) + ( Xd_0__inst_mult_5_365  ))
// Xd_0__inst_mult_5_369  = CARRY(( !Xd_0__inst_mult_5_568  $ (((!din_a[69]) # (!din_b[69]))) ) + ( Xd_0__inst_mult_5_366  ) + ( Xd_0__inst_mult_5_365  ))
// Xd_0__inst_mult_5_370  = SHARE((din_a[69] & (din_b[69] & Xd_0__inst_mult_5_568 )))

	.dataa(!din_a[69]),
	.datab(!din_b[69]),
	.datac(!Xd_0__inst_mult_5_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_365 ),
	.sharein(Xd_0__inst_mult_5_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_368 ),
	.cout(Xd_0__inst_mult_5_369 ),
	.shareout(Xd_0__inst_mult_5_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_59 (
// Equation(s):
// Xd_0__inst_mult_5_59_sumout  = SUM(( (din_a[70] & din_b[68]) ) + ( Xd_0__inst_mult_2_53  ) + ( Xd_0__inst_mult_2_52  ))
// Xd_0__inst_mult_5_60  = CARRY(( (din_a[70] & din_b[68]) ) + ( Xd_0__inst_mult_2_53  ) + ( Xd_0__inst_mult_2_52  ))
// Xd_0__inst_mult_5_61  = SHARE(GND)

	.dataa(!din_a[70]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_52 ),
	.sharein(Xd_0__inst_mult_2_53 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_59_sumout ),
	.cout(Xd_0__inst_mult_5_60 ),
	.shareout(Xd_0__inst_mult_5_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_117 (
// Equation(s):
// Xd_0__inst_mult_2_368  = SUM(( !Xd_0__inst_mult_2_568  $ (((!din_a[33]) # (!din_b[33]))) ) + ( Xd_0__inst_mult_2_366  ) + ( Xd_0__inst_mult_2_365  ))
// Xd_0__inst_mult_2_369  = CARRY(( !Xd_0__inst_mult_2_568  $ (((!din_a[33]) # (!din_b[33]))) ) + ( Xd_0__inst_mult_2_366  ) + ( Xd_0__inst_mult_2_365  ))
// Xd_0__inst_mult_2_370  = SHARE((din_a[33] & (din_b[33] & Xd_0__inst_mult_2_568 )))

	.dataa(!din_a[33]),
	.datab(!din_b[33]),
	.datac(!Xd_0__inst_mult_2_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_365 ),
	.sharein(Xd_0__inst_mult_2_366 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_368 ),
	.cout(Xd_0__inst_mult_2_369 ),
	.shareout(Xd_0__inst_mult_2_370 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_121 (
// Equation(s):
// Xd_0__inst_mult_3_396  = SUM(( !Xd_0__inst_mult_3_173  $ (((!din_a[45]) # (!din_b[45]))) ) + ( Xd_0__inst_mult_3_394  ) + ( Xd_0__inst_mult_3_393  ))
// Xd_0__inst_mult_3_397  = CARRY(( !Xd_0__inst_mult_3_173  $ (((!din_a[45]) # (!din_b[45]))) ) + ( Xd_0__inst_mult_3_394  ) + ( Xd_0__inst_mult_3_393  ))
// Xd_0__inst_mult_3_398  = SHARE((din_a[45] & (din_b[45] & Xd_0__inst_mult_3_173 )))

	.dataa(!din_a[45]),
	.datab(!din_b[45]),
	.datac(!Xd_0__inst_mult_3_173 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_393 ),
	.sharein(Xd_0__inst_mult_3_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_396 ),
	.cout(Xd_0__inst_mult_3_397 ),
	.shareout(Xd_0__inst_mult_3_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_47 (
// Equation(s):
// Xd_0__inst_mult_3_47_sumout  = SUM(( (din_a[46] & din_b[44]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_48  = CARRY(( (din_a[46] & din_b[44]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_49  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_47_sumout ),
	.cout(Xd_0__inst_mult_3_48 ),
	.shareout(Xd_0__inst_mult_3_49 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_115 (
// Equation(s):
// Xd_0__inst_mult_0_372  = SUM(( !Xd_0__inst_mult_0_564  $ (((!din_a[9]) # (!din_b[9]))) ) + ( Xd_0__inst_mult_0_370  ) + ( Xd_0__inst_mult_0_369  ))
// Xd_0__inst_mult_0_373  = CARRY(( !Xd_0__inst_mult_0_564  $ (((!din_a[9]) # (!din_b[9]))) ) + ( Xd_0__inst_mult_0_370  ) + ( Xd_0__inst_mult_0_369  ))
// Xd_0__inst_mult_0_374  = SHARE((din_a[9] & (din_b[9] & Xd_0__inst_mult_0_564 )))

	.dataa(!din_a[9]),
	.datab(!din_b[9]),
	.datac(!Xd_0__inst_mult_0_564 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_369 ),
	.sharein(Xd_0__inst_mult_0_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_372 ),
	.cout(Xd_0__inst_mult_0_373 ),
	.shareout(Xd_0__inst_mult_0_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_115 (
// Equation(s):
// Xd_0__inst_mult_1_372  = SUM(( !Xd_0__inst_mult_1_568  $ (((!din_a[21]) # (!din_b[21]))) ) + ( Xd_0__inst_mult_1_370  ) + ( Xd_0__inst_mult_1_369  ))
// Xd_0__inst_mult_1_373  = CARRY(( !Xd_0__inst_mult_1_568  $ (((!din_a[21]) # (!din_b[21]))) ) + ( Xd_0__inst_mult_1_370  ) + ( Xd_0__inst_mult_1_369  ))
// Xd_0__inst_mult_1_374  = SHARE((din_a[21] & (din_b[21] & Xd_0__inst_mult_1_568 )))

	.dataa(!din_a[21]),
	.datab(!din_b[21]),
	.datac(!Xd_0__inst_mult_1_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_369 ),
	.sharein(Xd_0__inst_mult_1_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_372 ),
	.cout(Xd_0__inst_mult_1_373 ),
	.shareout(Xd_0__inst_mult_1_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_167 (
// Equation(s):
// Xd_0__inst_mult_6_568  = SUM(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_6_566  ) + ( Xd_0__inst_mult_6_565  ))
// Xd_0__inst_mult_6_569  = CARRY(( (din_a[80] & din_b[82]) ) + ( Xd_0__inst_mult_6_566  ) + ( Xd_0__inst_mult_6_565  ))
// Xd_0__inst_mult_6_570  = SHARE(GND)

	.dataa(!din_a[80]),
	.datab(!din_b[82]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_565 ),
	.sharein(Xd_0__inst_mult_6_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_568 ),
	.cout(Xd_0__inst_mult_6_569 ),
	.shareout(Xd_0__inst_mult_6_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_166 (
// Equation(s):
// Xd_0__inst_mult_7_564  = SUM(( (din_a[92] & din_b[94]) ) + ( Xd_0__inst_mult_7_562  ) + ( Xd_0__inst_mult_7_561  ))
// Xd_0__inst_mult_7_565  = CARRY(( (din_a[92] & din_b[94]) ) + ( Xd_0__inst_mult_7_562  ) + ( Xd_0__inst_mult_7_561  ))
// Xd_0__inst_mult_7_566  = SHARE(GND)

	.dataa(!din_a[92]),
	.datab(!din_b[94]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_561 ),
	.sharein(Xd_0__inst_mult_7_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_564 ),
	.cout(Xd_0__inst_mult_7_565 ),
	.shareout(Xd_0__inst_mult_7_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_4_119 (
// Equation(s):
// Xd_0__inst_mult_4_376  = SUM(( !Xd_0__inst_mult_4_572  $ (((!din_a[57]) # (!din_b[58]))) ) + ( Xd_0__inst_mult_4_374  ) + ( Xd_0__inst_mult_4_373  ))
// Xd_0__inst_mult_4_377  = CARRY(( !Xd_0__inst_mult_4_572  $ (((!din_a[57]) # (!din_b[58]))) ) + ( Xd_0__inst_mult_4_374  ) + ( Xd_0__inst_mult_4_373  ))
// Xd_0__inst_mult_4_378  = SHARE((din_a[57] & (din_b[58] & Xd_0__inst_mult_4_572 )))

	.dataa(!din_a[57]),
	.datab(!din_b[58]),
	.datac(!Xd_0__inst_mult_4_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_373 ),
	.sharein(Xd_0__inst_mult_4_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_376 ),
	.cout(Xd_0__inst_mult_4_377 ),
	.shareout(Xd_0__inst_mult_4_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_51 (
// Equation(s):
// Xd_0__inst_mult_4_51_sumout  = SUM(( (din_a[58] & din_b[57]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_52  = CARRY(( (din_a[58] & din_b[57]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_53  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[57]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_51_sumout ),
	.cout(Xd_0__inst_mult_4_52 ),
	.shareout(Xd_0__inst_mult_4_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_5_118 (
// Equation(s):
// Xd_0__inst_mult_5_372  = SUM(( !Xd_0__inst_mult_5_572  $ (((!din_a[69]) # (!din_b[70]))) ) + ( Xd_0__inst_mult_5_370  ) + ( Xd_0__inst_mult_5_369  ))
// Xd_0__inst_mult_5_373  = CARRY(( !Xd_0__inst_mult_5_572  $ (((!din_a[69]) # (!din_b[70]))) ) + ( Xd_0__inst_mult_5_370  ) + ( Xd_0__inst_mult_5_369  ))
// Xd_0__inst_mult_5_374  = SHARE((din_a[69] & (din_b[70] & Xd_0__inst_mult_5_572 )))

	.dataa(!din_a[69]),
	.datab(!din_b[70]),
	.datac(!Xd_0__inst_mult_5_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_369 ),
	.sharein(Xd_0__inst_mult_5_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_372 ),
	.cout(Xd_0__inst_mult_5_373 ),
	.shareout(Xd_0__inst_mult_5_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_2_118 (
// Equation(s):
// Xd_0__inst_mult_2_372  = SUM(( !Xd_0__inst_mult_2_572  $ (((!din_a[33]) # (!din_b[34]))) ) + ( Xd_0__inst_mult_2_370  ) + ( Xd_0__inst_mult_2_369  ))
// Xd_0__inst_mult_2_373  = CARRY(( !Xd_0__inst_mult_2_572  $ (((!din_a[33]) # (!din_b[34]))) ) + ( Xd_0__inst_mult_2_370  ) + ( Xd_0__inst_mult_2_369  ))
// Xd_0__inst_mult_2_374  = SHARE((din_a[33] & (din_b[34] & Xd_0__inst_mult_2_572 )))

	.dataa(!din_a[33]),
	.datab(!din_b[34]),
	.datac(!Xd_0__inst_mult_2_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_369 ),
	.sharein(Xd_0__inst_mult_2_370 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_372 ),
	.cout(Xd_0__inst_mult_2_373 ),
	.shareout(Xd_0__inst_mult_2_374 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_3_122 (
// Equation(s):
// Xd_0__inst_mult_3_400  = SUM(( !Xd_0__inst_mult_3_169  $ (((!din_a[45]) # (!din_b[46]))) ) + ( Xd_0__inst_mult_3_398  ) + ( Xd_0__inst_mult_3_397  ))
// Xd_0__inst_mult_3_401  = CARRY(( !Xd_0__inst_mult_3_169  $ (((!din_a[45]) # (!din_b[46]))) ) + ( Xd_0__inst_mult_3_398  ) + ( Xd_0__inst_mult_3_397  ))
// Xd_0__inst_mult_3_402  = SHARE((din_a[45] & (din_b[46] & Xd_0__inst_mult_3_169 )))

	.dataa(!din_a[45]),
	.datab(!din_b[46]),
	.datac(!Xd_0__inst_mult_3_169 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_397 ),
	.sharein(Xd_0__inst_mult_3_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_400 ),
	.cout(Xd_0__inst_mult_3_401 ),
	.shareout(Xd_0__inst_mult_3_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_51 (
// Equation(s):
// Xd_0__inst_mult_3_51_sumout  = SUM(( (din_a[46] & din_b[45]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_52  = CARRY(( (din_a[46] & din_b[45]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_53  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[45]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_51_sumout ),
	.cout(Xd_0__inst_mult_3_52 ),
	.shareout(Xd_0__inst_mult_3_53 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_0_116 (
// Equation(s):
// Xd_0__inst_mult_0_376  = SUM(( !Xd_0__inst_mult_0_568  $ (((!din_a[9]) # (!din_b[10]))) ) + ( Xd_0__inst_mult_0_374  ) + ( Xd_0__inst_mult_0_373  ))
// Xd_0__inst_mult_0_377  = CARRY(( !Xd_0__inst_mult_0_568  $ (((!din_a[9]) # (!din_b[10]))) ) + ( Xd_0__inst_mult_0_374  ) + ( Xd_0__inst_mult_0_373  ))
// Xd_0__inst_mult_0_378  = SHARE((din_a[9] & (din_b[10] & Xd_0__inst_mult_0_568 )))

	.dataa(!din_a[9]),
	.datab(!din_b[10]),
	.datac(!Xd_0__inst_mult_0_568 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_373 ),
	.sharein(Xd_0__inst_mult_0_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_376 ),
	.cout(Xd_0__inst_mult_0_377 ),
	.shareout(Xd_0__inst_mult_0_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000010100001E1E),
	.shared_arith("on")
) Xd_0__inst_mult_1_116 (
// Equation(s):
// Xd_0__inst_mult_1_376  = SUM(( !Xd_0__inst_mult_1_572  $ (((!din_a[21]) # (!din_b[22]))) ) + ( Xd_0__inst_mult_1_374  ) + ( Xd_0__inst_mult_1_373  ))
// Xd_0__inst_mult_1_377  = CARRY(( !Xd_0__inst_mult_1_572  $ (((!din_a[21]) # (!din_b[22]))) ) + ( Xd_0__inst_mult_1_374  ) + ( Xd_0__inst_mult_1_373  ))
// Xd_0__inst_mult_1_378  = SHARE((din_a[21] & (din_b[22] & Xd_0__inst_mult_1_572 )))

	.dataa(!din_a[21]),
	.datab(!din_b[22]),
	.datac(!Xd_0__inst_mult_1_572 ),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_373 ),
	.sharein(Xd_0__inst_mult_1_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_376 ),
	.cout(Xd_0__inst_mult_1_377 ),
	.shareout(Xd_0__inst_mult_1_378 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_168 (
// Equation(s):
// Xd_0__inst_mult_6_572  = SUM(( GND ) + ( Xd_0__inst_mult_6_570  ) + ( Xd_0__inst_mult_6_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_569 ),
	.sharein(Xd_0__inst_mult_6_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_6_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_167 (
// Equation(s):
// Xd_0__inst_mult_7_568  = SUM(( GND ) + ( Xd_0__inst_mult_7_566  ) + ( Xd_0__inst_mult_7_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_565 ),
	.sharein(Xd_0__inst_mult_7_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_120 (
// Equation(s):
// Xd_0__inst_mult_4_380  = SUM(( GND ) + ( Xd_0__inst_mult_4_378  ) + ( Xd_0__inst_mult_4_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_377 ),
	.sharein(Xd_0__inst_mult_4_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_55 (
// Equation(s):
// Xd_0__inst_mult_4_55_sumout  = SUM(( (din_a[58] & din_b[58]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_56  = CARRY(( (din_a[58] & din_b[58]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_57  = SHARE(GND)

	.dataa(!din_a[58]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_55_sumout ),
	.cout(Xd_0__inst_mult_4_56 ),
	.shareout(Xd_0__inst_mult_4_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_119 (
// Equation(s):
// Xd_0__inst_mult_5_376  = SUM(( GND ) + ( Xd_0__inst_mult_5_374  ) + ( Xd_0__inst_mult_5_373  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_373 ),
	.sharein(Xd_0__inst_mult_5_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_376 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_119 (
// Equation(s):
// Xd_0__inst_mult_2_376  = SUM(( GND ) + ( Xd_0__inst_mult_2_374  ) + ( Xd_0__inst_mult_2_373  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_373 ),
	.sharein(Xd_0__inst_mult_2_374 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_376 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_123 (
// Equation(s):
// Xd_0__inst_mult_3_404  = SUM(( GND ) + ( Xd_0__inst_mult_3_402  ) + ( Xd_0__inst_mult_3_401  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_401 ),
	.sharein(Xd_0__inst_mult_3_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_404 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_55 (
// Equation(s):
// Xd_0__inst_mult_3_55_sumout  = SUM(( (din_a[46] & din_b[46]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_56  = CARRY(( (din_a[46] & din_b[46]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_57  = SHARE(GND)

	.dataa(!din_a[46]),
	.datab(!din_b[46]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_3_55_sumout ),
	.cout(Xd_0__inst_mult_3_56 ),
	.shareout(Xd_0__inst_mult_3_57 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_117 (
// Equation(s):
// Xd_0__inst_mult_0_380  = SUM(( GND ) + ( Xd_0__inst_mult_0_378  ) + ( Xd_0__inst_mult_0_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_377 ),
	.sharein(Xd_0__inst_mult_0_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_117 (
// Equation(s):
// Xd_0__inst_mult_1_380  = SUM(( GND ) + ( Xd_0__inst_mult_1_378  ) + ( Xd_0__inst_mult_1_377  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_377 ),
	.sharein(Xd_0__inst_mult_1_378 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_380 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_124 (
// Equation(s):
// Xd_0__inst_mult_3_408  = SUM(( (!din_a[45] & (((din_a[44] & din_b[40])))) # (din_a[45] & (!din_b[39] $ (((!din_a[44]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_514  ) + ( Xd_0__inst_mult_3_513  ))
// Xd_0__inst_mult_3_409  = CARRY(( (!din_a[45] & (((din_a[44] & din_b[40])))) # (din_a[45] & (!din_b[39] $ (((!din_a[44]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_514  ) + ( Xd_0__inst_mult_3_513  ))
// Xd_0__inst_mult_3_410  = SHARE((din_a[45] & (din_b[39] & (din_a[44] & din_b[40]))))

	.dataa(!din_a[45]),
	.datab(!din_b[39]),
	.datac(!din_a[44]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_513 ),
	.sharein(Xd_0__inst_mult_3_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_408 ),
	.cout(Xd_0__inst_mult_3_409 ),
	.shareout(Xd_0__inst_mult_3_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_125 (
// Equation(s):
// Xd_0__inst_mult_3_412  = SUM(( GND ) + ( Xd_0__inst_mult_3_510  ) + ( Xd_0__inst_mult_3_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_509 ),
	.sharein(Xd_0__inst_mult_3_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_412 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_118 (
// Equation(s):
// Xd_0__inst_mult_0_384  = SUM(( (!din_a[9] & (((din_a[8] & din_b[4])))) # (din_a[9] & (!din_b[3] $ (((!din_a[8]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_486  ) + ( Xd_0__inst_mult_0_485  ))
// Xd_0__inst_mult_0_385  = CARRY(( (!din_a[9] & (((din_a[8] & din_b[4])))) # (din_a[9] & (!din_b[3] $ (((!din_a[8]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_486  ) + ( Xd_0__inst_mult_0_485  ))
// Xd_0__inst_mult_0_386  = SHARE((din_a[9] & (din_b[3] & (din_a[8] & din_b[4]))))

	.dataa(!din_a[9]),
	.datab(!din_b[3]),
	.datac(!din_a[8]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_485 ),
	.sharein(Xd_0__inst_mult_0_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_384 ),
	.cout(Xd_0__inst_mult_0_385 ),
	.shareout(Xd_0__inst_mult_0_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_119 (
// Equation(s):
// Xd_0__inst_mult_0_388  = SUM(( GND ) + ( Xd_0__inst_mult_0_482  ) + ( Xd_0__inst_mult_0_481  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_481 ),
	.sharein(Xd_0__inst_mult_0_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_388 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_126 (
// Equation(s):
// Xd_0__inst_mult_3_416  = SUM(( (din_a[40] & din_b[45]) ) + ( Xd_0__inst_mult_3_534  ) + ( Xd_0__inst_mult_3_533  ))
// Xd_0__inst_mult_3_417  = CARRY(( (din_a[40] & din_b[45]) ) + ( Xd_0__inst_mult_3_534  ) + ( Xd_0__inst_mult_3_533  ))
// Xd_0__inst_mult_3_418  = SHARE((din_a[40] & din_b[46]))

	.dataa(!din_a[40]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_533 ),
	.sharein(Xd_0__inst_mult_3_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_416 ),
	.cout(Xd_0__inst_mult_3_417 ),
	.shareout(Xd_0__inst_mult_3_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_121 (
// Equation(s):
// Xd_0__inst_mult_4_384  = SUM(( (!din_a[50] & (((din_a[51] & din_b[48])))) # (din_a[50] & (!din_b[49] $ (((!din_a[51]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_250  ) + ( Xd_0__inst_mult_4_249  ))
// Xd_0__inst_mult_4_385  = CARRY(( (!din_a[50] & (((din_a[51] & din_b[48])))) # (din_a[50] & (!din_b[49] $ (((!din_a[51]) # (!din_b[48]))))) ) + ( Xd_0__inst_mult_4_250  ) + ( Xd_0__inst_mult_4_249  ))
// Xd_0__inst_mult_4_386  = SHARE((din_a[50] & (din_b[49] & (din_a[51] & din_b[48]))))

	.dataa(!din_a[50]),
	.datab(!din_b[49]),
	.datac(!din_a[51]),
	.datad(!din_b[48]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_249 ),
	.sharein(Xd_0__inst_mult_4_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_384 ),
	.cout(Xd_0__inst_mult_4_385 ),
	.shareout(Xd_0__inst_mult_4_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_122 (
// Equation(s):
// Xd_0__inst_mult_4_388  = SUM(( (din_a[45] & din_b[36]) ) + ( Xd_0__inst_mult_2_69  ) + ( Xd_0__inst_mult_2_68  ))
// Xd_0__inst_mult_4_389  = CARRY(( (din_a[45] & din_b[36]) ) + ( Xd_0__inst_mult_2_69  ) + ( Xd_0__inst_mult_2_68  ))
// Xd_0__inst_mult_4_390  = SHARE(Xd_0__inst_mult_4_384 )

	.dataa(!din_a[45]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_4_384 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_68 ),
	.sharein(Xd_0__inst_mult_2_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_388 ),
	.cout(Xd_0__inst_mult_4_389 ),
	.shareout(Xd_0__inst_mult_4_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_120 (
// Equation(s):
// Xd_0__inst_mult_5_380  = SUM(( (!din_a[62] & (((din_a[63] & din_b[60])))) # (din_a[62] & (!din_b[61] $ (((!din_a[63]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_250  ) + ( Xd_0__inst_mult_5_249  ))
// Xd_0__inst_mult_5_381  = CARRY(( (!din_a[62] & (((din_a[63] & din_b[60])))) # (din_a[62] & (!din_b[61] $ (((!din_a[63]) # (!din_b[60]))))) ) + ( Xd_0__inst_mult_5_250  ) + ( Xd_0__inst_mult_5_249  ))
// Xd_0__inst_mult_5_382  = SHARE((din_a[62] & (din_b[61] & (din_a[63] & din_b[60]))))

	.dataa(!din_a[62]),
	.datab(!din_b[61]),
	.datac(!din_a[63]),
	.datad(!din_b[60]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_249 ),
	.sharein(Xd_0__inst_mult_5_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_380 ),
	.cout(Xd_0__inst_mult_5_381 ),
	.shareout(Xd_0__inst_mult_5_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_121 (
// Equation(s):
// Xd_0__inst_mult_5_384  = SUM(( (din_a[8] & din_b[0]) ) + ( Xd_0__inst_mult_3_65  ) + ( Xd_0__inst_mult_3_64  ))
// Xd_0__inst_mult_5_385  = CARRY(( (din_a[8] & din_b[0]) ) + ( Xd_0__inst_mult_3_65  ) + ( Xd_0__inst_mult_3_64  ))
// Xd_0__inst_mult_5_386  = SHARE(Xd_0__inst_mult_5_380 )

	.dataa(!din_a[8]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_5_380 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_64 ),
	.sharein(Xd_0__inst_mult_3_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_384 ),
	.cout(Xd_0__inst_mult_5_385 ),
	.shareout(Xd_0__inst_mult_5_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_120 (
// Equation(s):
// Xd_0__inst_mult_2_380  = SUM(( (!din_a[26] & (((din_a[27] & din_b[24])))) # (din_a[26] & (!din_b[25] $ (((!din_a[27]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_250  ) + ( Xd_0__inst_mult_2_249  ))
// Xd_0__inst_mult_2_381  = CARRY(( (!din_a[26] & (((din_a[27] & din_b[24])))) # (din_a[26] & (!din_b[25] $ (((!din_a[27]) # (!din_b[24]))))) ) + ( Xd_0__inst_mult_2_250  ) + ( Xd_0__inst_mult_2_249  ))
// Xd_0__inst_mult_2_382  = SHARE((din_a[26] & (din_b[25] & (din_a[27] & din_b[24]))))

	.dataa(!din_a[26]),
	.datab(!din_b[25]),
	.datac(!din_a[27]),
	.datad(!din_b[24]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_249 ),
	.sharein(Xd_0__inst_mult_2_250 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_380 ),
	.cout(Xd_0__inst_mult_2_381 ),
	.shareout(Xd_0__inst_mult_2_382 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000FF00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_121 (
// Equation(s):
// Xd_0__inst_mult_2_384  = SUM(( (din_a[19] & din_b[12]) ) + ( Xd_0__inst_mult_0_65  ) + ( Xd_0__inst_mult_0_64  ))
// Xd_0__inst_mult_2_385  = CARRY(( (din_a[19] & din_b[12]) ) + ( Xd_0__inst_mult_0_65  ) + ( Xd_0__inst_mult_0_64  ))
// Xd_0__inst_mult_2_386  = SHARE(Xd_0__inst_mult_2_380 )

	.dataa(!din_a[19]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(!Xd_0__inst_mult_2_380 ),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_64 ),
	.sharein(Xd_0__inst_mult_0_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_384 ),
	.cout(Xd_0__inst_mult_2_385 ),
	.shareout(Xd_0__inst_mult_2_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_127 (
// Equation(s):
// Xd_0__inst_mult_3_420  = SUM(( (!din_a[38] & (((din_a[39] & din_b[36])))) # (din_a[38] & (!din_b[37] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_282  ) + ( Xd_0__inst_mult_3_281  ))
// Xd_0__inst_mult_3_421  = CARRY(( (!din_a[38] & (((din_a[39] & din_b[36])))) # (din_a[38] & (!din_b[37] $ (((!din_a[39]) # (!din_b[36]))))) ) + ( Xd_0__inst_mult_3_282  ) + ( Xd_0__inst_mult_3_281  ))
// Xd_0__inst_mult_3_422  = SHARE((din_a[38] & (din_b[37] & (din_a[39] & din_b[36]))))

	.dataa(!din_a[38]),
	.datab(!din_b[37]),
	.datac(!din_a[39]),
	.datad(!din_b[36]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_281 ),
	.sharein(Xd_0__inst_mult_3_282 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_420 ),
	.cout(Xd_0__inst_mult_3_421 ),
	.shareout(Xd_0__inst_mult_3_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_128 (
// Equation(s):
// Xd_0__inst_mult_3_425  = CARRY(( GND ) + ( Xd_0__inst_mult_2_61  ) + ( Xd_0__inst_mult_2_60  ))
// Xd_0__inst_mult_3_426  = SHARE(Xd_0__inst_mult_3_420 )

	.dataa(!Xd_0__inst_mult_3_420 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_60 ),
	.sharein(Xd_0__inst_mult_2_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_425 ),
	.shareout(Xd_0__inst_mult_3_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_120 (
// Equation(s):
// Xd_0__inst_mult_0_392  = SUM(( (!din_a[2] & (((din_a[3] & din_b[0])))) # (din_a[2] & (!din_b[1] $ (((!din_a[3]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_262  ) + ( Xd_0__inst_mult_0_261  ))
// Xd_0__inst_mult_0_393  = CARRY(( (!din_a[2] & (((din_a[3] & din_b[0])))) # (din_a[2] & (!din_b[1] $ (((!din_a[3]) # (!din_b[0]))))) ) + ( Xd_0__inst_mult_0_262  ) + ( Xd_0__inst_mult_0_261  ))
// Xd_0__inst_mult_0_394  = SHARE((din_a[2] & (din_b[1] & (din_a[3] & din_b[0]))))

	.dataa(!din_a[2]),
	.datab(!din_b[1]),
	.datac(!din_a[3]),
	.datad(!din_b[0]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_261 ),
	.sharein(Xd_0__inst_mult_0_262 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_392 ),
	.cout(Xd_0__inst_mult_0_393 ),
	.shareout(Xd_0__inst_mult_0_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000555500000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_121 (
// Equation(s):
// Xd_0__inst_mult_0_397  = CARRY(( GND ) + ( Xd_0__inst_mult_4_61  ) + ( Xd_0__inst_mult_4_60  ))
// Xd_0__inst_mult_0_398  = SHARE(Xd_0__inst_mult_0_392 )

	.dataa(!Xd_0__inst_mult_0_392 ),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_60 ),
	.sharein(Xd_0__inst_mult_4_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_397 ),
	.shareout(Xd_0__inst_mult_0_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_63 (
// Equation(s):
// Xd_0__inst_mult_5_63_sumout  = SUM(( (din_a[67] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_64  = CARRY(( (din_a[67] & din_b[60]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_65  = SHARE(GND)

	.dataa(!din_a[67]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_5_63_sumout ),
	.cout(Xd_0__inst_mult_5_64 ),
	.shareout(Xd_0__inst_mult_5_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_123 (
// Equation(s):
// Xd_0__inst_mult_4_393  = CARRY(( (din_a[51] & din_b[49]) ) + ( Xd_0__inst_mult_4_578  ) + ( Xd_0__inst_mult_4_577  ))
// Xd_0__inst_mult_4_394  = SHARE((din_a[50] & din_b[50]))

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(!din_a[50]),
	.datad(!din_b[50]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_577 ),
	.sharein(Xd_0__inst_mult_4_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_393 ),
	.shareout(Xd_0__inst_mult_4_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_122 (
// Equation(s):
// Xd_0__inst_mult_5_389  = CARRY(( (din_a[63] & din_b[61]) ) + ( Xd_0__inst_mult_5_578  ) + ( Xd_0__inst_mult_5_577  ))
// Xd_0__inst_mult_5_390  = SHARE((din_a[62] & din_b[62]))

	.dataa(!din_a[63]),
	.datab(!din_b[61]),
	.datac(!din_a[62]),
	.datad(!din_b[62]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_577 ),
	.sharein(Xd_0__inst_mult_5_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_389 ),
	.shareout(Xd_0__inst_mult_5_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_122 (
// Equation(s):
// Xd_0__inst_mult_2_389  = CARRY(( (din_a[27] & din_b[25]) ) + ( Xd_0__inst_mult_2_578  ) + ( Xd_0__inst_mult_2_577  ))
// Xd_0__inst_mult_2_390  = SHARE((din_a[26] & din_b[26]))

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(!din_a[26]),
	.datad(!din_b[26]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_577 ),
	.sharein(Xd_0__inst_mult_2_578 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_389 ),
	.shareout(Xd_0__inst_mult_2_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_129 (
// Equation(s):
// Xd_0__inst_mult_3_429  = CARRY(( (din_a[39] & din_b[37]) ) + ( Xd_0__inst_mult_3_570  ) + ( Xd_0__inst_mult_3_569  ))
// Xd_0__inst_mult_3_430  = SHARE((din_a[38] & din_b[38]))

	.dataa(!din_a[39]),
	.datab(!din_b[37]),
	.datac(!din_a[38]),
	.datad(!din_b[38]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_569 ),
	.sharein(Xd_0__inst_mult_3_570 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_429 ),
	.shareout(Xd_0__inst_mult_3_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_122 (
// Equation(s):
// Xd_0__inst_mult_0_401  = CARRY(( (din_a[3] & din_b[1]) ) + ( Xd_0__inst_mult_0_574  ) + ( Xd_0__inst_mult_0_573  ))
// Xd_0__inst_mult_0_402  = SHARE((din_a[2] & din_b[2]))

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(!din_a[2]),
	.datad(!din_b[2]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_573 ),
	.sharein(Xd_0__inst_mult_0_574 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_401 ),
	.shareout(Xd_0__inst_mult_0_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_118 (
// Equation(s):
// Xd_0__inst_mult_1_385  = CARRY(( (din_a[15] & din_b[13]) ) + ( Xd_0__inst_mult_1_550  ) + ( Xd_0__inst_mult_1_549  ))
// Xd_0__inst_mult_1_386  = SHARE((din_a[14] & din_b[14]))

	.dataa(!din_a[15]),
	.datab(!din_b[13]),
	.datac(!din_a[14]),
	.datad(!din_b[14]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_549 ),
	.sharein(Xd_0__inst_mult_1_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_385 ),
	.shareout(Xd_0__inst_mult_1_386 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_168 (
// Equation(s):
// Xd_0__inst_mult_7_572  = SUM(( GND ) + ( Xd_0__inst_mult_4_542  ) + ( Xd_0__inst_mult_4_541  ))
// Xd_0__inst_mult_7_573  = CARRY(( GND ) + ( Xd_0__inst_mult_4_542  ) + ( Xd_0__inst_mult_4_541  ))
// Xd_0__inst_mult_7_574  = SHARE(VCC)

	.dataa(!din_a[87]),
	.datab(!din_b[85]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_541 ),
	.sharein(Xd_0__inst_mult_4_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_7_572 ),
	.cout(Xd_0__inst_mult_7_573 ),
	.shareout(Xd_0__inst_mult_7_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_124 (
// Equation(s):
// Xd_0__inst_mult_4_396  = SUM(( (din_a[53] & din_b[48]) ) + ( Xd_0__inst_mult_4_266  ) + ( Xd_0__inst_mult_4_265  ))
// Xd_0__inst_mult_4_397  = CARRY(( (din_a[53] & din_b[48]) ) + ( Xd_0__inst_mult_4_266  ) + ( Xd_0__inst_mult_4_265  ))
// Xd_0__inst_mult_4_398  = SHARE((din_b[48] & din_a[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[48]),
	.datac(!din_a[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_265 ),
	.sharein(Xd_0__inst_mult_4_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_396 ),
	.cout(Xd_0__inst_mult_4_397 ),
	.shareout(Xd_0__inst_mult_4_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_125 (
// Equation(s):
// Xd_0__inst_mult_4_400  = SUM(( (din_a[51] & din_b[50]) ) + ( Xd_0__inst_mult_4_270  ) + ( Xd_0__inst_mult_4_269  ))
// Xd_0__inst_mult_4_401  = CARRY(( (din_a[51] & din_b[50]) ) + ( Xd_0__inst_mult_4_270  ) + ( Xd_0__inst_mult_4_269  ))
// Xd_0__inst_mult_4_402  = SHARE((din_b[50] & din_a[52]))

	.dataa(!din_a[51]),
	.datab(!din_b[50]),
	.datac(!din_a[52]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_269 ),
	.sharein(Xd_0__inst_mult_4_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_400 ),
	.cout(Xd_0__inst_mult_4_401 ),
	.shareout(Xd_0__inst_mult_4_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_59 (
// Equation(s):
// Xd_0__inst_mult_0_59_sumout  = SUM(( (din_a[10] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_60  = CARRY(( (din_a[10] & din_b[0]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_61  = SHARE(GND)

	.dataa(!din_a[10]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_0_59_sumout ),
	.cout(Xd_0__inst_mult_0_60 ),
	.shareout(Xd_0__inst_mult_0_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_123 (
// Equation(s):
// Xd_0__inst_mult_5_392  = SUM(( (din_a[65] & din_b[60]) ) + ( Xd_0__inst_mult_5_266  ) + ( Xd_0__inst_mult_5_265  ))
// Xd_0__inst_mult_5_393  = CARRY(( (din_a[65] & din_b[60]) ) + ( Xd_0__inst_mult_5_266  ) + ( Xd_0__inst_mult_5_265  ))
// Xd_0__inst_mult_5_394  = SHARE((din_b[60] & din_a[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[60]),
	.datac(!din_a[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_265 ),
	.sharein(Xd_0__inst_mult_5_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_392 ),
	.cout(Xd_0__inst_mult_5_393 ),
	.shareout(Xd_0__inst_mult_5_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_124 (
// Equation(s):
// Xd_0__inst_mult_5_396  = SUM(( (din_a[63] & din_b[62]) ) + ( Xd_0__inst_mult_5_270  ) + ( Xd_0__inst_mult_5_269  ))
// Xd_0__inst_mult_5_397  = CARRY(( (din_a[63] & din_b[62]) ) + ( Xd_0__inst_mult_5_270  ) + ( Xd_0__inst_mult_5_269  ))
// Xd_0__inst_mult_5_398  = SHARE((din_b[62] & din_a[64]))

	.dataa(!din_a[63]),
	.datab(!din_b[62]),
	.datac(!din_a[64]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_269 ),
	.sharein(Xd_0__inst_mult_5_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_396 ),
	.cout(Xd_0__inst_mult_5_397 ),
	.shareout(Xd_0__inst_mult_5_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_123 (
// Equation(s):
// Xd_0__inst_mult_2_392  = SUM(( (din_a[29] & din_b[24]) ) + ( Xd_0__inst_mult_2_266  ) + ( Xd_0__inst_mult_2_265  ))
// Xd_0__inst_mult_2_393  = CARRY(( (din_a[29] & din_b[24]) ) + ( Xd_0__inst_mult_2_266  ) + ( Xd_0__inst_mult_2_265  ))
// Xd_0__inst_mult_2_394  = SHARE((din_b[24] & din_a[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[24]),
	.datac(!din_a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_265 ),
	.sharein(Xd_0__inst_mult_2_266 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_392 ),
	.cout(Xd_0__inst_mult_2_393 ),
	.shareout(Xd_0__inst_mult_2_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_124 (
// Equation(s):
// Xd_0__inst_mult_2_396  = SUM(( (din_a[27] & din_b[26]) ) + ( Xd_0__inst_mult_2_270  ) + ( Xd_0__inst_mult_2_269  ))
// Xd_0__inst_mult_2_397  = CARRY(( (din_a[27] & din_b[26]) ) + ( Xd_0__inst_mult_2_270  ) + ( Xd_0__inst_mult_2_269  ))
// Xd_0__inst_mult_2_398  = SHARE((din_b[26] & din_a[28]))

	.dataa(!din_a[27]),
	.datab(!din_b[26]),
	.datac(!din_a[28]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_269 ),
	.sharein(Xd_0__inst_mult_2_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_396 ),
	.cout(Xd_0__inst_mult_2_397 ),
	.shareout(Xd_0__inst_mult_2_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_130 (
// Equation(s):
// Xd_0__inst_mult_3_432  = SUM(( (din_a[41] & din_b[36]) ) + ( Xd_0__inst_mult_3_310  ) + ( Xd_0__inst_mult_3_309  ))
// Xd_0__inst_mult_3_433  = CARRY(( (din_a[41] & din_b[36]) ) + ( Xd_0__inst_mult_3_310  ) + ( Xd_0__inst_mult_3_309  ))
// Xd_0__inst_mult_3_434  = SHARE((din_b[36] & din_a[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[36]),
	.datac(!din_a[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_309 ),
	.sharein(Xd_0__inst_mult_3_310 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_432 ),
	.cout(Xd_0__inst_mult_3_433 ),
	.shareout(Xd_0__inst_mult_3_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_131 (
// Equation(s):
// Xd_0__inst_mult_3_436  = SUM(( (din_a[39] & din_b[38]) ) + ( Xd_0__inst_mult_3_314  ) + ( Xd_0__inst_mult_3_313  ))
// Xd_0__inst_mult_3_437  = CARRY(( (din_a[39] & din_b[38]) ) + ( Xd_0__inst_mult_3_314  ) + ( Xd_0__inst_mult_3_313  ))
// Xd_0__inst_mult_3_438  = SHARE((din_b[38] & din_a[40]))

	.dataa(!din_a[39]),
	.datab(!din_b[38]),
	.datac(!din_a[40]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_313 ),
	.sharein(Xd_0__inst_mult_3_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_436 ),
	.cout(Xd_0__inst_mult_3_437 ),
	.shareout(Xd_0__inst_mult_3_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_59 (
// Equation(s):
// Xd_0__inst_mult_1_59_sumout  = SUM(( (din_a[22] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_60  = CARRY(( (din_a[22] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_61  = SHARE(GND)

	.dataa(!din_a[22]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_59_sumout ),
	.cout(Xd_0__inst_mult_1_60 ),
	.shareout(Xd_0__inst_mult_1_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_123 (
// Equation(s):
// Xd_0__inst_mult_0_404  = SUM(( (din_a[5] & din_b[0]) ) + ( Xd_0__inst_mult_0_286  ) + ( Xd_0__inst_mult_0_285  ))
// Xd_0__inst_mult_0_405  = CARRY(( (din_a[5] & din_b[0]) ) + ( Xd_0__inst_mult_0_286  ) + ( Xd_0__inst_mult_0_285  ))
// Xd_0__inst_mult_0_406  = SHARE((din_b[0] & din_a[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[0]),
	.datac(!din_a[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_285 ),
	.sharein(Xd_0__inst_mult_0_286 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_404 ),
	.cout(Xd_0__inst_mult_0_405 ),
	.shareout(Xd_0__inst_mult_0_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_124 (
// Equation(s):
// Xd_0__inst_mult_0_408  = SUM(( (din_a[3] & din_b[2]) ) + ( Xd_0__inst_mult_0_290  ) + ( Xd_0__inst_mult_0_289  ))
// Xd_0__inst_mult_0_409  = CARRY(( (din_a[3] & din_b[2]) ) + ( Xd_0__inst_mult_0_290  ) + ( Xd_0__inst_mult_0_289  ))
// Xd_0__inst_mult_0_410  = SHARE((din_b[2] & din_a[4]))

	.dataa(!din_a[3]),
	.datab(!din_b[2]),
	.datac(!din_a[4]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_289 ),
	.sharein(Xd_0__inst_mult_0_290 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_408 ),
	.cout(Xd_0__inst_mult_0_409 ),
	.shareout(Xd_0__inst_mult_0_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_119 (
// Equation(s):
// Xd_0__inst_mult_1_388  = SUM(( (din_a[17] & din_b[12]) ) + ( Xd_0__inst_mult_1_270  ) + ( Xd_0__inst_mult_1_269  ))
// Xd_0__inst_mult_1_389  = CARRY(( (din_a[17] & din_b[12]) ) + ( Xd_0__inst_mult_1_270  ) + ( Xd_0__inst_mult_1_269  ))
// Xd_0__inst_mult_1_390  = SHARE((din_b[12] & din_a[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[12]),
	.datac(!din_a[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_269 ),
	.sharein(Xd_0__inst_mult_1_270 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_388 ),
	.cout(Xd_0__inst_mult_1_389 ),
	.shareout(Xd_0__inst_mult_1_390 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_120 (
// Equation(s):
// Xd_0__inst_mult_1_392  = SUM(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_1_274  ) + ( Xd_0__inst_mult_1_273  ))
// Xd_0__inst_mult_1_393  = CARRY(( (din_a[15] & din_b[14]) ) + ( Xd_0__inst_mult_1_274  ) + ( Xd_0__inst_mult_1_273  ))
// Xd_0__inst_mult_1_394  = SHARE((din_b[14] & din_a[16]))

	.dataa(!din_a[15]),
	.datab(!din_b[14]),
	.datac(!din_a[16]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_273 ),
	.sharein(Xd_0__inst_mult_1_274 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_392 ),
	.cout(Xd_0__inst_mult_1_393 ),
	.shareout(Xd_0__inst_mult_1_394 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_126 (
// Equation(s):
// Xd_0__inst_mult_4_404  = SUM(( (din_a[53] & din_b[49]) ) + ( Xd_0__inst_mult_4_398  ) + ( Xd_0__inst_mult_4_397  ))
// Xd_0__inst_mult_4_405  = CARRY(( (din_a[53] & din_b[49]) ) + ( Xd_0__inst_mult_4_398  ) + ( Xd_0__inst_mult_4_397  ))
// Xd_0__inst_mult_4_406  = SHARE((din_b[49] & din_a[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[49]),
	.datac(!din_a[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_397 ),
	.sharein(Xd_0__inst_mult_4_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_404 ),
	.cout(Xd_0__inst_mult_4_405 ),
	.shareout(Xd_0__inst_mult_4_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_127 (
// Equation(s):
// Xd_0__inst_mult_4_408  = SUM(( (!din_a[51] & (((din_a[50] & din_b[52])))) # (din_a[51] & (!din_b[51] $ (((!din_a[50]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_402  ) + ( Xd_0__inst_mult_4_401  ))
// Xd_0__inst_mult_4_409  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[52])))) # (din_a[51] & (!din_b[51] $ (((!din_a[50]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_402  ) + ( Xd_0__inst_mult_4_401  ))
// Xd_0__inst_mult_4_410  = SHARE((din_a[51] & (din_b[51] & (din_a[50] & din_b[52]))))

	.dataa(!din_a[51]),
	.datab(!din_b[51]),
	.datac(!din_a[50]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_401 ),
	.sharein(Xd_0__inst_mult_4_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_408 ),
	.cout(Xd_0__inst_mult_4_409 ),
	.shareout(Xd_0__inst_mult_4_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_125 (
// Equation(s):
// Xd_0__inst_mult_5_400  = SUM(( (din_a[65] & din_b[61]) ) + ( Xd_0__inst_mult_5_394  ) + ( Xd_0__inst_mult_5_393  ))
// Xd_0__inst_mult_5_401  = CARRY(( (din_a[65] & din_b[61]) ) + ( Xd_0__inst_mult_5_394  ) + ( Xd_0__inst_mult_5_393  ))
// Xd_0__inst_mult_5_402  = SHARE((din_b[61] & din_a[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[61]),
	.datac(!din_a[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_393 ),
	.sharein(Xd_0__inst_mult_5_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_400 ),
	.cout(Xd_0__inst_mult_5_401 ),
	.shareout(Xd_0__inst_mult_5_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_126 (
// Equation(s):
// Xd_0__inst_mult_5_404  = SUM(( (!din_a[63] & (((din_a[62] & din_b[64])))) # (din_a[63] & (!din_b[63] $ (((!din_a[62]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_398  ) + ( Xd_0__inst_mult_5_397  ))
// Xd_0__inst_mult_5_405  = CARRY(( (!din_a[63] & (((din_a[62] & din_b[64])))) # (din_a[63] & (!din_b[63] $ (((!din_a[62]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_398  ) + ( Xd_0__inst_mult_5_397  ))
// Xd_0__inst_mult_5_406  = SHARE((din_a[63] & (din_b[63] & (din_a[62] & din_b[64]))))

	.dataa(!din_a[63]),
	.datab(!din_b[63]),
	.datac(!din_a[62]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_397 ),
	.sharein(Xd_0__inst_mult_5_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_404 ),
	.cout(Xd_0__inst_mult_5_405 ),
	.shareout(Xd_0__inst_mult_5_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_125 (
// Equation(s):
// Xd_0__inst_mult_2_400  = SUM(( (din_a[29] & din_b[25]) ) + ( Xd_0__inst_mult_2_394  ) + ( Xd_0__inst_mult_2_393  ))
// Xd_0__inst_mult_2_401  = CARRY(( (din_a[29] & din_b[25]) ) + ( Xd_0__inst_mult_2_394  ) + ( Xd_0__inst_mult_2_393  ))
// Xd_0__inst_mult_2_402  = SHARE((din_b[25] & din_a[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[25]),
	.datac(!din_a[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_393 ),
	.sharein(Xd_0__inst_mult_2_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_400 ),
	.cout(Xd_0__inst_mult_2_401 ),
	.shareout(Xd_0__inst_mult_2_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_126 (
// Equation(s):
// Xd_0__inst_mult_2_404  = SUM(( (!din_a[27] & (((din_a[26] & din_b[28])))) # (din_a[27] & (!din_b[27] $ (((!din_a[26]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_398  ) + ( Xd_0__inst_mult_2_397  ))
// Xd_0__inst_mult_2_405  = CARRY(( (!din_a[27] & (((din_a[26] & din_b[28])))) # (din_a[27] & (!din_b[27] $ (((!din_a[26]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_398  ) + ( Xd_0__inst_mult_2_397  ))
// Xd_0__inst_mult_2_406  = SHARE((din_a[27] & (din_b[27] & (din_a[26] & din_b[28]))))

	.dataa(!din_a[27]),
	.datab(!din_b[27]),
	.datac(!din_a[26]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_397 ),
	.sharein(Xd_0__inst_mult_2_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_404 ),
	.cout(Xd_0__inst_mult_2_405 ),
	.shareout(Xd_0__inst_mult_2_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_132 (
// Equation(s):
// Xd_0__inst_mult_3_440  = SUM(( (din_a[41] & din_b[37]) ) + ( Xd_0__inst_mult_3_434  ) + ( Xd_0__inst_mult_3_433  ))
// Xd_0__inst_mult_3_441  = CARRY(( (din_a[41] & din_b[37]) ) + ( Xd_0__inst_mult_3_434  ) + ( Xd_0__inst_mult_3_433  ))
// Xd_0__inst_mult_3_442  = SHARE((din_b[37] & din_a[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[37]),
	.datac(!din_a[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_433 ),
	.sharein(Xd_0__inst_mult_3_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_440 ),
	.cout(Xd_0__inst_mult_3_441 ),
	.shareout(Xd_0__inst_mult_3_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_133 (
// Equation(s):
// Xd_0__inst_mult_3_444  = SUM(( (!din_a[39] & (((din_a[38] & din_b[40])))) # (din_a[39] & (!din_b[39] $ (((!din_a[38]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_438  ) + ( Xd_0__inst_mult_3_437  ))
// Xd_0__inst_mult_3_445  = CARRY(( (!din_a[39] & (((din_a[38] & din_b[40])))) # (din_a[39] & (!din_b[39] $ (((!din_a[38]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_438  ) + ( Xd_0__inst_mult_3_437  ))
// Xd_0__inst_mult_3_446  = SHARE((din_a[39] & (din_b[39] & (din_a[38] & din_b[40]))))

	.dataa(!din_a[39]),
	.datab(!din_b[39]),
	.datac(!din_a[38]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_437 ),
	.sharein(Xd_0__inst_mult_3_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_444 ),
	.cout(Xd_0__inst_mult_3_445 ),
	.shareout(Xd_0__inst_mult_3_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_125 (
// Equation(s):
// Xd_0__inst_mult_0_412  = SUM(( (din_a[5] & din_b[1]) ) + ( Xd_0__inst_mult_0_406  ) + ( Xd_0__inst_mult_0_405  ))
// Xd_0__inst_mult_0_413  = CARRY(( (din_a[5] & din_b[1]) ) + ( Xd_0__inst_mult_0_406  ) + ( Xd_0__inst_mult_0_405  ))
// Xd_0__inst_mult_0_414  = SHARE((din_b[1] & din_a[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[1]),
	.datac(!din_a[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_405 ),
	.sharein(Xd_0__inst_mult_0_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_412 ),
	.cout(Xd_0__inst_mult_0_413 ),
	.shareout(Xd_0__inst_mult_0_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_126 (
// Equation(s):
// Xd_0__inst_mult_0_416  = SUM(( (!din_a[3] & (((din_a[2] & din_b[4])))) # (din_a[3] & (!din_b[3] $ (((!din_a[2]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_410  ) + ( Xd_0__inst_mult_0_409  ))
// Xd_0__inst_mult_0_417  = CARRY(( (!din_a[3] & (((din_a[2] & din_b[4])))) # (din_a[3] & (!din_b[3] $ (((!din_a[2]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_410  ) + ( Xd_0__inst_mult_0_409  ))
// Xd_0__inst_mult_0_418  = SHARE((din_a[3] & (din_b[3] & (din_a[2] & din_b[4]))))

	.dataa(!din_a[3]),
	.datab(!din_b[3]),
	.datac(!din_a[2]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_409 ),
	.sharein(Xd_0__inst_mult_0_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_416 ),
	.cout(Xd_0__inst_mult_0_417 ),
	.shareout(Xd_0__inst_mult_0_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_121 (
// Equation(s):
// Xd_0__inst_mult_1_396  = SUM(( (din_a[17] & din_b[13]) ) + ( Xd_0__inst_mult_1_390  ) + ( Xd_0__inst_mult_1_389  ))
// Xd_0__inst_mult_1_397  = CARRY(( (din_a[17] & din_b[13]) ) + ( Xd_0__inst_mult_1_390  ) + ( Xd_0__inst_mult_1_389  ))
// Xd_0__inst_mult_1_398  = SHARE((din_b[13] & din_a[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[13]),
	.datac(!din_a[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_389 ),
	.sharein(Xd_0__inst_mult_1_390 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_396 ),
	.cout(Xd_0__inst_mult_1_397 ),
	.shareout(Xd_0__inst_mult_1_398 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_122 (
// Equation(s):
// Xd_0__inst_mult_1_400  = SUM(( (!din_a[15] & (((din_a[14] & din_b[16])))) # (din_a[15] & (!din_b[15] $ (((!din_a[14]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_394  ) + ( Xd_0__inst_mult_1_393  ))
// Xd_0__inst_mult_1_401  = CARRY(( (!din_a[15] & (((din_a[14] & din_b[16])))) # (din_a[15] & (!din_b[15] $ (((!din_a[14]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_394  ) + ( Xd_0__inst_mult_1_393  ))
// Xd_0__inst_mult_1_402  = SHARE((din_a[15] & (din_b[15] & (din_a[14] & din_b[16]))))

	.dataa(!din_a[15]),
	.datab(!din_b[15]),
	.datac(!din_a[14]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_393 ),
	.sharein(Xd_0__inst_mult_1_394 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_400 ),
	.cout(Xd_0__inst_mult_1_401 ),
	.shareout(Xd_0__inst_mult_1_402 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_128 (
// Equation(s):
// Xd_0__inst_mult_4_412  = SUM(( (din_a[53] & din_b[50]) ) + ( Xd_0__inst_mult_4_406  ) + ( Xd_0__inst_mult_4_405  ))
// Xd_0__inst_mult_4_413  = CARRY(( (din_a[53] & din_b[50]) ) + ( Xd_0__inst_mult_4_406  ) + ( Xd_0__inst_mult_4_405  ))
// Xd_0__inst_mult_4_414  = SHARE((din_a[55] & din_b[49]))

	.dataa(!din_a[53]),
	.datab(!din_b[50]),
	.datac(!din_a[55]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_405 ),
	.sharein(Xd_0__inst_mult_4_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_412 ),
	.cout(Xd_0__inst_mult_4_413 ),
	.shareout(Xd_0__inst_mult_4_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_129 (
// Equation(s):
// Xd_0__inst_mult_4_416  = SUM(( (!din_a[52] & (((din_a[51] & din_b[52])))) # (din_a[52] & (!din_b[51] $ (((!din_a[51]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_410  ) + ( Xd_0__inst_mult_4_409  ))
// Xd_0__inst_mult_4_417  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[52])))) # (din_a[52] & (!din_b[51] $ (((!din_a[51]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_410  ) + ( Xd_0__inst_mult_4_409  ))
// Xd_0__inst_mult_4_418  = SHARE((din_a[52] & (din_b[51] & (din_a[51] & din_b[52]))))

	.dataa(!din_a[52]),
	.datab(!din_b[51]),
	.datac(!din_a[51]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_409 ),
	.sharein(Xd_0__inst_mult_4_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_416 ),
	.cout(Xd_0__inst_mult_4_417 ),
	.shareout(Xd_0__inst_mult_4_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_59 (
// Equation(s):
// Xd_0__inst_mult_4_59_sumout  = SUM(( (din_a[55] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_60  = CARRY(( (din_a[55] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_61  = SHARE(GND)

	.dataa(!din_a[55]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_59_sumout ),
	.cout(Xd_0__inst_mult_4_60 ),
	.shareout(Xd_0__inst_mult_4_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_127 (
// Equation(s):
// Xd_0__inst_mult_5_408  = SUM(( (din_a[65] & din_b[62]) ) + ( Xd_0__inst_mult_5_402  ) + ( Xd_0__inst_mult_5_401  ))
// Xd_0__inst_mult_5_409  = CARRY(( (din_a[65] & din_b[62]) ) + ( Xd_0__inst_mult_5_402  ) + ( Xd_0__inst_mult_5_401  ))
// Xd_0__inst_mult_5_410  = SHARE((din_a[67] & din_b[61]))

	.dataa(!din_a[65]),
	.datab(!din_b[62]),
	.datac(!din_a[67]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_401 ),
	.sharein(Xd_0__inst_mult_5_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_408 ),
	.cout(Xd_0__inst_mult_5_409 ),
	.shareout(Xd_0__inst_mult_5_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_128 (
// Equation(s):
// Xd_0__inst_mult_5_412  = SUM(( (!din_a[64] & (((din_a[63] & din_b[64])))) # (din_a[64] & (!din_b[63] $ (((!din_a[63]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_406  ) + ( Xd_0__inst_mult_5_405  ))
// Xd_0__inst_mult_5_413  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[64])))) # (din_a[64] & (!din_b[63] $ (((!din_a[63]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_406  ) + ( Xd_0__inst_mult_5_405  ))
// Xd_0__inst_mult_5_414  = SHARE((din_a[64] & (din_b[63] & (din_a[63] & din_b[64]))))

	.dataa(!din_a[64]),
	.datab(!din_b[63]),
	.datac(!din_a[63]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_405 ),
	.sharein(Xd_0__inst_mult_5_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_412 ),
	.cout(Xd_0__inst_mult_5_413 ),
	.shareout(Xd_0__inst_mult_5_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_127 (
// Equation(s):
// Xd_0__inst_mult_2_408  = SUM(( (din_a[29] & din_b[26]) ) + ( Xd_0__inst_mult_2_402  ) + ( Xd_0__inst_mult_2_401  ))
// Xd_0__inst_mult_2_409  = CARRY(( (din_a[29] & din_b[26]) ) + ( Xd_0__inst_mult_2_402  ) + ( Xd_0__inst_mult_2_401  ))
// Xd_0__inst_mult_2_410  = SHARE((din_a[31] & din_b[25]))

	.dataa(!din_a[29]),
	.datab(!din_b[26]),
	.datac(!din_a[31]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_401 ),
	.sharein(Xd_0__inst_mult_2_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_408 ),
	.cout(Xd_0__inst_mult_2_409 ),
	.shareout(Xd_0__inst_mult_2_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_128 (
// Equation(s):
// Xd_0__inst_mult_2_412  = SUM(( (!din_a[28] & (((din_a[27] & din_b[28])))) # (din_a[28] & (!din_b[27] $ (((!din_a[27]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_406  ) + ( Xd_0__inst_mult_2_405  ))
// Xd_0__inst_mult_2_413  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[28])))) # (din_a[28] & (!din_b[27] $ (((!din_a[27]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_406  ) + ( Xd_0__inst_mult_2_405  ))
// Xd_0__inst_mult_2_414  = SHARE((din_a[28] & (din_b[27] & (din_a[27] & din_b[28]))))

	.dataa(!din_a[28]),
	.datab(!din_b[27]),
	.datac(!din_a[27]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_405 ),
	.sharein(Xd_0__inst_mult_2_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_412 ),
	.cout(Xd_0__inst_mult_2_413 ),
	.shareout(Xd_0__inst_mult_2_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_59 (
// Equation(s):
// Xd_0__inst_mult_2_59_sumout  = SUM(( (din_a[31] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_60  = CARRY(( (din_a[31] & din_b[24]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_61  = SHARE(GND)

	.dataa(!din_a[31]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_2_59_sumout ),
	.cout(Xd_0__inst_mult_2_60 ),
	.shareout(Xd_0__inst_mult_2_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_134 (
// Equation(s):
// Xd_0__inst_mult_3_448  = SUM(( (din_a[41] & din_b[38]) ) + ( Xd_0__inst_mult_3_442  ) + ( Xd_0__inst_mult_3_441  ))
// Xd_0__inst_mult_3_449  = CARRY(( (din_a[41] & din_b[38]) ) + ( Xd_0__inst_mult_3_442  ) + ( Xd_0__inst_mult_3_441  ))
// Xd_0__inst_mult_3_450  = SHARE((din_a[43] & din_b[37]))

	.dataa(!din_a[41]),
	.datab(!din_b[38]),
	.datac(!din_a[43]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_441 ),
	.sharein(Xd_0__inst_mult_3_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_448 ),
	.cout(Xd_0__inst_mult_3_449 ),
	.shareout(Xd_0__inst_mult_3_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_135 (
// Equation(s):
// Xd_0__inst_mult_3_452  = SUM(( (!din_a[40] & (((din_a[39] & din_b[40])))) # (din_a[40] & (!din_b[39] $ (((!din_a[39]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_446  ) + ( Xd_0__inst_mult_3_445  ))
// Xd_0__inst_mult_3_453  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[40])))) # (din_a[40] & (!din_b[39] $ (((!din_a[39]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_446  ) + ( Xd_0__inst_mult_3_445  ))
// Xd_0__inst_mult_3_454  = SHARE((din_a[40] & (din_b[39] & (din_a[39] & din_b[40]))))

	.dataa(!din_a[40]),
	.datab(!din_b[39]),
	.datac(!din_a[39]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_445 ),
	.sharein(Xd_0__inst_mult_3_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_452 ),
	.cout(Xd_0__inst_mult_3_453 ),
	.shareout(Xd_0__inst_mult_3_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_59 (
// Equation(s):
// Xd_0__inst_mult_3_59_sumout  = SUM(( (din_a[43] & din_b[36]) ) + ( Xd_0__inst_mult_4_69  ) + ( Xd_0__inst_mult_4_68  ))
// Xd_0__inst_mult_3_60  = CARRY(( (din_a[43] & din_b[36]) ) + ( Xd_0__inst_mult_4_69  ) + ( Xd_0__inst_mult_4_68  ))
// Xd_0__inst_mult_3_61  = SHARE(GND)

	.dataa(!din_a[43]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_68 ),
	.sharein(Xd_0__inst_mult_4_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_59_sumout ),
	.cout(Xd_0__inst_mult_3_60 ),
	.shareout(Xd_0__inst_mult_3_61 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_127 (
// Equation(s):
// Xd_0__inst_mult_0_420  = SUM(( (din_a[5] & din_b[2]) ) + ( Xd_0__inst_mult_0_414  ) + ( Xd_0__inst_mult_0_413  ))
// Xd_0__inst_mult_0_421  = CARRY(( (din_a[5] & din_b[2]) ) + ( Xd_0__inst_mult_0_414  ) + ( Xd_0__inst_mult_0_413  ))
// Xd_0__inst_mult_0_422  = SHARE((din_a[7] & din_b[1]))

	.dataa(!din_a[5]),
	.datab(!din_b[2]),
	.datac(!din_a[7]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_413 ),
	.sharein(Xd_0__inst_mult_0_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_420 ),
	.cout(Xd_0__inst_mult_0_421 ),
	.shareout(Xd_0__inst_mult_0_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_128 (
// Equation(s):
// Xd_0__inst_mult_0_424  = SUM(( (!din_a[4] & (((din_a[3] & din_b[4])))) # (din_a[4] & (!din_b[3] $ (((!din_a[3]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_418  ) + ( Xd_0__inst_mult_0_417  ))
// Xd_0__inst_mult_0_425  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[4])))) # (din_a[4] & (!din_b[3] $ (((!din_a[3]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_418  ) + ( Xd_0__inst_mult_0_417  ))
// Xd_0__inst_mult_0_426  = SHARE((din_a[4] & (din_b[3] & (din_a[3] & din_b[4]))))

	.dataa(!din_a[4]),
	.datab(!din_b[3]),
	.datac(!din_a[3]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_417 ),
	.sharein(Xd_0__inst_mult_0_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_424 ),
	.cout(Xd_0__inst_mult_0_425 ),
	.shareout(Xd_0__inst_mult_0_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_63 (
// Equation(s):
// Xd_0__inst_mult_0_63_sumout  = SUM(( (din_a[7] & din_b[0]) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_0_64  = CARRY(( (din_a[7] & din_b[0]) ) + ( Xd_0__inst_mult_7_37  ) + ( Xd_0__inst_mult_7_36  ))
// Xd_0__inst_mult_0_65  = SHARE(GND)

	.dataa(!din_a[7]),
	.datab(!din_b[0]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_36 ),
	.sharein(Xd_0__inst_mult_7_37 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_63_sumout ),
	.cout(Xd_0__inst_mult_0_64 ),
	.shareout(Xd_0__inst_mult_0_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_123 (
// Equation(s):
// Xd_0__inst_mult_1_404  = SUM(( (din_a[17] & din_b[14]) ) + ( Xd_0__inst_mult_1_398  ) + ( Xd_0__inst_mult_1_397  ))
// Xd_0__inst_mult_1_405  = CARRY(( (din_a[17] & din_b[14]) ) + ( Xd_0__inst_mult_1_398  ) + ( Xd_0__inst_mult_1_397  ))
// Xd_0__inst_mult_1_406  = SHARE((din_a[19] & din_b[13]))

	.dataa(!din_a[17]),
	.datab(!din_b[14]),
	.datac(!din_a[19]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_397 ),
	.sharein(Xd_0__inst_mult_1_398 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_404 ),
	.cout(Xd_0__inst_mult_1_405 ),
	.shareout(Xd_0__inst_mult_1_406 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_124 (
// Equation(s):
// Xd_0__inst_mult_1_408  = SUM(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_402  ) + ( Xd_0__inst_mult_1_401  ))
// Xd_0__inst_mult_1_409  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[16])))) # (din_a[16] & (!din_b[15] $ (((!din_a[15]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_402  ) + ( Xd_0__inst_mult_1_401  ))
// Xd_0__inst_mult_1_410  = SHARE((din_a[16] & (din_b[15] & (din_a[15] & din_b[16]))))

	.dataa(!din_a[16]),
	.datab(!din_b[15]),
	.datac(!din_a[15]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_401 ),
	.sharein(Xd_0__inst_mult_1_402 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_408 ),
	.cout(Xd_0__inst_mult_1_409 ),
	.shareout(Xd_0__inst_mult_1_410 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_130 (
// Equation(s):
// Xd_0__inst_mult_4_420  = SUM(( (din_a[54] & din_b[50]) ) + ( Xd_0__inst_mult_4_414  ) + ( Xd_0__inst_mult_4_413  ))
// Xd_0__inst_mult_4_421  = CARRY(( (din_a[54] & din_b[50]) ) + ( Xd_0__inst_mult_4_414  ) + ( Xd_0__inst_mult_4_413  ))
// Xd_0__inst_mult_4_422  = SHARE((din_a[56] & din_b[49]))

	.dataa(!din_a[54]),
	.datab(!din_b[50]),
	.datac(!din_a[56]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_413 ),
	.sharein(Xd_0__inst_mult_4_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_420 ),
	.cout(Xd_0__inst_mult_4_421 ),
	.shareout(Xd_0__inst_mult_4_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_131 (
// Equation(s):
// Xd_0__inst_mult_4_424  = SUM(( (!din_a[53] & (((din_a[52] & din_b[52])))) # (din_a[53] & (!din_b[51] $ (((!din_a[52]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_418  ) + ( Xd_0__inst_mult_4_417  ))
// Xd_0__inst_mult_4_425  = CARRY(( (!din_a[53] & (((din_a[52] & din_b[52])))) # (din_a[53] & (!din_b[51] $ (((!din_a[52]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_418  ) + ( Xd_0__inst_mult_4_417  ))
// Xd_0__inst_mult_4_426  = SHARE((din_a[53] & (din_b[51] & (din_a[52] & din_b[52]))))

	.dataa(!din_a[53]),
	.datab(!din_b[51]),
	.datac(!din_a[52]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_417 ),
	.sharein(Xd_0__inst_mult_4_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_424 ),
	.cout(Xd_0__inst_mult_4_425 ),
	.shareout(Xd_0__inst_mult_4_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_63 (
// Equation(s):
// Xd_0__inst_mult_4_63_sumout  = SUM(( (din_a[56] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_64  = CARRY(( (din_a[56] & din_b[48]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_65  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_4_63_sumout ),
	.cout(Xd_0__inst_mult_4_64 ),
	.shareout(Xd_0__inst_mult_4_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_132 (
// Equation(s):
// Xd_0__inst_mult_4_428  = SUM(( (!din_a[50] & (((din_a[51] & din_b[53])))) # (din_a[50] & (!din_b[54] $ (((!din_a[51]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_294  ) + ( Xd_0__inst_mult_4_293  ))
// Xd_0__inst_mult_4_429  = CARRY(( (!din_a[50] & (((din_a[51] & din_b[53])))) # (din_a[50] & (!din_b[54] $ (((!din_a[51]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_294  ) + ( Xd_0__inst_mult_4_293  ))
// Xd_0__inst_mult_4_430  = SHARE((din_a[50] & (din_b[54] & (din_a[51] & din_b[53]))))

	.dataa(!din_a[50]),
	.datab(!din_b[54]),
	.datac(!din_a[51]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_293 ),
	.sharein(Xd_0__inst_mult_4_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_428 ),
	.cout(Xd_0__inst_mult_4_429 ),
	.shareout(Xd_0__inst_mult_4_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_133 (
// Equation(s):
// Xd_0__inst_mult_4_433  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_434  = SHARE((din_a[48] & din_b[56]))

	.dataa(!din_a[48]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_433 ),
	.shareout(Xd_0__inst_mult_4_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_129 (
// Equation(s):
// Xd_0__inst_mult_5_416  = SUM(( (din_a[66] & din_b[62]) ) + ( Xd_0__inst_mult_5_410  ) + ( Xd_0__inst_mult_5_409  ))
// Xd_0__inst_mult_5_417  = CARRY(( (din_a[66] & din_b[62]) ) + ( Xd_0__inst_mult_5_410  ) + ( Xd_0__inst_mult_5_409  ))
// Xd_0__inst_mult_5_418  = SHARE((din_a[68] & din_b[61]))

	.dataa(!din_a[66]),
	.datab(!din_b[62]),
	.datac(!din_a[68]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_409 ),
	.sharein(Xd_0__inst_mult_5_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_416 ),
	.cout(Xd_0__inst_mult_5_417 ),
	.shareout(Xd_0__inst_mult_5_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_130 (
// Equation(s):
// Xd_0__inst_mult_5_420  = SUM(( (!din_a[65] & (((din_a[64] & din_b[64])))) # (din_a[65] & (!din_b[63] $ (((!din_a[64]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_414  ) + ( Xd_0__inst_mult_5_413  ))
// Xd_0__inst_mult_5_421  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[64])))) # (din_a[65] & (!din_b[63] $ (((!din_a[64]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_414  ) + ( Xd_0__inst_mult_5_413  ))
// Xd_0__inst_mult_5_422  = SHARE((din_a[65] & (din_b[63] & (din_a[64] & din_b[64]))))

	.dataa(!din_a[65]),
	.datab(!din_b[63]),
	.datac(!din_a[64]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_413 ),
	.sharein(Xd_0__inst_mult_5_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_420 ),
	.cout(Xd_0__inst_mult_5_421 ),
	.shareout(Xd_0__inst_mult_5_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_67 (
// Equation(s):
// Xd_0__inst_mult_5_67_sumout  = SUM(( (din_a[68] & din_b[60]) ) + ( Xd_0__inst_mult_4_65  ) + ( Xd_0__inst_mult_4_64  ))
// Xd_0__inst_mult_5_68  = CARRY(( (din_a[68] & din_b[60]) ) + ( Xd_0__inst_mult_4_65  ) + ( Xd_0__inst_mult_4_64  ))
// Xd_0__inst_mult_5_69  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[60]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_64 ),
	.sharein(Xd_0__inst_mult_4_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_67_sumout ),
	.cout(Xd_0__inst_mult_5_68 ),
	.shareout(Xd_0__inst_mult_5_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_131 (
// Equation(s):
// Xd_0__inst_mult_5_424  = SUM(( (!din_a[62] & (((din_a[63] & din_b[65])))) # (din_a[62] & (!din_b[66] $ (((!din_a[63]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_294  ) + ( Xd_0__inst_mult_5_293  ))
// Xd_0__inst_mult_5_425  = CARRY(( (!din_a[62] & (((din_a[63] & din_b[65])))) # (din_a[62] & (!din_b[66] $ (((!din_a[63]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_294  ) + ( Xd_0__inst_mult_5_293  ))
// Xd_0__inst_mult_5_426  = SHARE((din_a[62] & (din_b[66] & (din_a[63] & din_b[65]))))

	.dataa(!din_a[62]),
	.datab(!din_b[66]),
	.datac(!din_a[63]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_293 ),
	.sharein(Xd_0__inst_mult_5_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_424 ),
	.cout(Xd_0__inst_mult_5_425 ),
	.shareout(Xd_0__inst_mult_5_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_132 (
// Equation(s):
// Xd_0__inst_mult_5_429  = CARRY(( GND ) + ( Xd_0__inst_mult_6_61  ) + ( Xd_0__inst_mult_6_60  ))
// Xd_0__inst_mult_5_430  = SHARE((din_a[60] & din_b[68]))

	.dataa(!din_a[60]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_60 ),
	.sharein(Xd_0__inst_mult_6_61 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_429 ),
	.shareout(Xd_0__inst_mult_5_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_129 (
// Equation(s):
// Xd_0__inst_mult_2_416  = SUM(( (din_a[30] & din_b[26]) ) + ( Xd_0__inst_mult_2_410  ) + ( Xd_0__inst_mult_2_409  ))
// Xd_0__inst_mult_2_417  = CARRY(( (din_a[30] & din_b[26]) ) + ( Xd_0__inst_mult_2_410  ) + ( Xd_0__inst_mult_2_409  ))
// Xd_0__inst_mult_2_418  = SHARE((din_a[32] & din_b[25]))

	.dataa(!din_a[30]),
	.datab(!din_b[26]),
	.datac(!din_a[32]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_409 ),
	.sharein(Xd_0__inst_mult_2_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_416 ),
	.cout(Xd_0__inst_mult_2_417 ),
	.shareout(Xd_0__inst_mult_2_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_130 (
// Equation(s):
// Xd_0__inst_mult_2_420  = SUM(( (!din_a[29] & (((din_a[28] & din_b[28])))) # (din_a[29] & (!din_b[27] $ (((!din_a[28]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_414  ) + ( Xd_0__inst_mult_2_413  ))
// Xd_0__inst_mult_2_421  = CARRY(( (!din_a[29] & (((din_a[28] & din_b[28])))) # (din_a[29] & (!din_b[27] $ (((!din_a[28]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_414  ) + ( Xd_0__inst_mult_2_413  ))
// Xd_0__inst_mult_2_422  = SHARE((din_a[29] & (din_b[27] & (din_a[28] & din_b[28]))))

	.dataa(!din_a[29]),
	.datab(!din_b[27]),
	.datac(!din_a[28]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_413 ),
	.sharein(Xd_0__inst_mult_2_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_420 ),
	.cout(Xd_0__inst_mult_2_421 ),
	.shareout(Xd_0__inst_mult_2_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_63 (
// Equation(s):
// Xd_0__inst_mult_2_63_sumout  = SUM(( (din_a[32] & din_b[24]) ) + ( Xd_0__inst_mult_5_69  ) + ( Xd_0__inst_mult_5_68  ))
// Xd_0__inst_mult_2_64  = CARRY(( (din_a[32] & din_b[24]) ) + ( Xd_0__inst_mult_5_69  ) + ( Xd_0__inst_mult_5_68  ))
// Xd_0__inst_mult_2_65  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_68 ),
	.sharein(Xd_0__inst_mult_5_69 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_63_sumout ),
	.cout(Xd_0__inst_mult_2_64 ),
	.shareout(Xd_0__inst_mult_2_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_131 (
// Equation(s):
// Xd_0__inst_mult_2_424  = SUM(( (!din_a[26] & (((din_a[27] & din_b[29])))) # (din_a[26] & (!din_b[30] $ (((!din_a[27]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_294  ) + ( Xd_0__inst_mult_2_293  ))
// Xd_0__inst_mult_2_425  = CARRY(( (!din_a[26] & (((din_a[27] & din_b[29])))) # (din_a[26] & (!din_b[30] $ (((!din_a[27]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_294  ) + ( Xd_0__inst_mult_2_293  ))
// Xd_0__inst_mult_2_426  = SHARE((din_a[26] & (din_b[30] & (din_a[27] & din_b[29]))))

	.dataa(!din_a[26]),
	.datab(!din_b[30]),
	.datac(!din_a[27]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_293 ),
	.sharein(Xd_0__inst_mult_2_294 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_424 ),
	.cout(Xd_0__inst_mult_2_425 ),
	.shareout(Xd_0__inst_mult_2_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_132 (
// Equation(s):
// Xd_0__inst_mult_2_429  = CARRY(( GND ) + ( Xd_0__inst_mult_4_45  ) + ( Xd_0__inst_mult_4_44  ))
// Xd_0__inst_mult_2_430  = SHARE((din_a[24] & din_b[32]))

	.dataa(!din_a[24]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_44 ),
	.sharein(Xd_0__inst_mult_4_45 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_429 ),
	.shareout(Xd_0__inst_mult_2_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_136 (
// Equation(s):
// Xd_0__inst_mult_3_456  = SUM(( (din_a[42] & din_b[38]) ) + ( Xd_0__inst_mult_3_450  ) + ( Xd_0__inst_mult_3_449  ))
// Xd_0__inst_mult_3_457  = CARRY(( (din_a[42] & din_b[38]) ) + ( Xd_0__inst_mult_3_450  ) + ( Xd_0__inst_mult_3_449  ))
// Xd_0__inst_mult_3_458  = SHARE((din_a[44] & din_b[37]))

	.dataa(!din_a[42]),
	.datab(!din_b[38]),
	.datac(!din_a[44]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_449 ),
	.sharein(Xd_0__inst_mult_3_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_456 ),
	.cout(Xd_0__inst_mult_3_457 ),
	.shareout(Xd_0__inst_mult_3_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_137 (
// Equation(s):
// Xd_0__inst_mult_3_460  = SUM(( (!din_a[41] & (((din_a[40] & din_b[40])))) # (din_a[41] & (!din_b[39] $ (((!din_a[40]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_454  ) + ( Xd_0__inst_mult_3_453  ))
// Xd_0__inst_mult_3_461  = CARRY(( (!din_a[41] & (((din_a[40] & din_b[40])))) # (din_a[41] & (!din_b[39] $ (((!din_a[40]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_454  ) + ( Xd_0__inst_mult_3_453  ))
// Xd_0__inst_mult_3_462  = SHARE((din_a[41] & (din_b[39] & (din_a[40] & din_b[40]))))

	.dataa(!din_a[41]),
	.datab(!din_b[39]),
	.datac(!din_a[40]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_453 ),
	.sharein(Xd_0__inst_mult_3_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_460 ),
	.cout(Xd_0__inst_mult_3_461 ),
	.shareout(Xd_0__inst_mult_3_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_63 (
// Equation(s):
// Xd_0__inst_mult_3_63_sumout  = SUM(( (din_a[44] & din_b[36]) ) + ( Xd_0__inst_mult_2_65  ) + ( Xd_0__inst_mult_2_64  ))
// Xd_0__inst_mult_3_64  = CARRY(( (din_a[44] & din_b[36]) ) + ( Xd_0__inst_mult_2_65  ) + ( Xd_0__inst_mult_2_64  ))
// Xd_0__inst_mult_3_65  = SHARE(GND)

	.dataa(!din_a[44]),
	.datab(!din_b[36]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_64 ),
	.sharein(Xd_0__inst_mult_2_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_63_sumout ),
	.cout(Xd_0__inst_mult_3_64 ),
	.shareout(Xd_0__inst_mult_3_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_138 (
// Equation(s):
// Xd_0__inst_mult_3_464  = SUM(( (!din_a[38] & (((din_a[39] & din_b[41])))) # (din_a[38] & (!din_b[42] $ (((!din_a[39]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_338  ) + ( Xd_0__inst_mult_3_337  ))
// Xd_0__inst_mult_3_465  = CARRY(( (!din_a[38] & (((din_a[39] & din_b[41])))) # (din_a[38] & (!din_b[42] $ (((!din_a[39]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_338  ) + ( Xd_0__inst_mult_3_337  ))
// Xd_0__inst_mult_3_466  = SHARE((din_a[38] & (din_b[42] & (din_a[39] & din_b[41]))))

	.dataa(!din_a[38]),
	.datab(!din_b[42]),
	.datac(!din_a[39]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_337 ),
	.sharein(Xd_0__inst_mult_3_338 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_464 ),
	.cout(Xd_0__inst_mult_3_465 ),
	.shareout(Xd_0__inst_mult_3_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_139 (
// Equation(s):
// Xd_0__inst_mult_3_469  = CARRY(( GND ) + ( Xd_0__inst_mult_4_49  ) + ( Xd_0__inst_mult_4_48  ))
// Xd_0__inst_mult_3_470  = SHARE((din_a[36] & din_b[44]))

	.dataa(!din_a[36]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_48 ),
	.sharein(Xd_0__inst_mult_4_49 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_469 ),
	.shareout(Xd_0__inst_mult_3_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_129 (
// Equation(s):
// Xd_0__inst_mult_0_428  = SUM(( (din_a[6] & din_b[2]) ) + ( Xd_0__inst_mult_0_422  ) + ( Xd_0__inst_mult_0_421  ))
// Xd_0__inst_mult_0_429  = CARRY(( (din_a[6] & din_b[2]) ) + ( Xd_0__inst_mult_0_422  ) + ( Xd_0__inst_mult_0_421  ))
// Xd_0__inst_mult_0_430  = SHARE((din_a[8] & din_b[1]))

	.dataa(!din_a[6]),
	.datab(!din_b[2]),
	.datac(!din_a[8]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_421 ),
	.sharein(Xd_0__inst_mult_0_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_428 ),
	.cout(Xd_0__inst_mult_0_429 ),
	.shareout(Xd_0__inst_mult_0_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_130 (
// Equation(s):
// Xd_0__inst_mult_0_432  = SUM(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_426  ) + ( Xd_0__inst_mult_0_425  ))
// Xd_0__inst_mult_0_433  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[4])))) # (din_a[5] & (!din_b[3] $ (((!din_a[4]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_426  ) + ( Xd_0__inst_mult_0_425  ))
// Xd_0__inst_mult_0_434  = SHARE((din_a[5] & (din_b[3] & (din_a[4] & din_b[4]))))

	.dataa(!din_a[5]),
	.datab(!din_b[3]),
	.datac(!din_a[4]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_425 ),
	.sharein(Xd_0__inst_mult_0_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_432 ),
	.cout(Xd_0__inst_mult_0_433 ),
	.shareout(Xd_0__inst_mult_0_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_131 (
// Equation(s):
// Xd_0__inst_mult_0_436  = SUM(( (!din_a[2] & (((din_a[3] & din_b[5])))) # (din_a[2] & (!din_b[6] $ (((!din_a[3]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_314  ) + ( Xd_0__inst_mult_0_313  ))
// Xd_0__inst_mult_0_437  = CARRY(( (!din_a[2] & (((din_a[3] & din_b[5])))) # (din_a[2] & (!din_b[6] $ (((!din_a[3]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_314  ) + ( Xd_0__inst_mult_0_313  ))
// Xd_0__inst_mult_0_438  = SHARE((din_a[2] & (din_b[6] & (din_a[3] & din_b[5]))))

	.dataa(!din_a[2]),
	.datab(!din_b[6]),
	.datac(!din_a[3]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_313 ),
	.sharein(Xd_0__inst_mult_0_314 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_436 ),
	.cout(Xd_0__inst_mult_0_437 ),
	.shareout(Xd_0__inst_mult_0_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_132 (
// Equation(s):
// Xd_0__inst_mult_0_441  = CARRY(( GND ) + ( Xd_0__inst_i29_15  ) + ( Xd_0__inst_i29_14  ))
// Xd_0__inst_mult_0_442  = SHARE((din_a[0] & din_b[8]))

	.dataa(!din_a[0]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_i29_14 ),
	.sharein(Xd_0__inst_i29_15 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_441 ),
	.shareout(Xd_0__inst_mult_0_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_125 (
// Equation(s):
// Xd_0__inst_mult_1_412  = SUM(( (din_a[18] & din_b[14]) ) + ( Xd_0__inst_mult_1_406  ) + ( Xd_0__inst_mult_1_405  ))
// Xd_0__inst_mult_1_413  = CARRY(( (din_a[18] & din_b[14]) ) + ( Xd_0__inst_mult_1_406  ) + ( Xd_0__inst_mult_1_405  ))
// Xd_0__inst_mult_1_414  = SHARE((din_a[20] & din_b[13]))

	.dataa(!din_a[18]),
	.datab(!din_b[14]),
	.datac(!din_a[20]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_405 ),
	.sharein(Xd_0__inst_mult_1_406 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_412 ),
	.cout(Xd_0__inst_mult_1_413 ),
	.shareout(Xd_0__inst_mult_1_414 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_126 (
// Equation(s):
// Xd_0__inst_mult_1_416  = SUM(( (!din_a[17] & (((din_a[16] & din_b[16])))) # (din_a[17] & (!din_b[15] $ (((!din_a[16]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_410  ) + ( Xd_0__inst_mult_1_409  ))
// Xd_0__inst_mult_1_417  = CARRY(( (!din_a[17] & (((din_a[16] & din_b[16])))) # (din_a[17] & (!din_b[15] $ (((!din_a[16]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_410  ) + ( Xd_0__inst_mult_1_409  ))
// Xd_0__inst_mult_1_418  = SHARE((din_a[17] & (din_b[15] & (din_a[16] & din_b[16]))))

	.dataa(!din_a[17]),
	.datab(!din_b[15]),
	.datac(!din_a[16]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_409 ),
	.sharein(Xd_0__inst_mult_1_410 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_416 ),
	.cout(Xd_0__inst_mult_1_417 ),
	.shareout(Xd_0__inst_mult_1_418 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_63 (
// Equation(s):
// Xd_0__inst_mult_1_63_sumout  = SUM(( (din_a[20] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_64  = CARRY(( (din_a[20] & din_b[12]) ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_65  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[12]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(Xd_0__inst_mult_1_63_sumout ),
	.cout(Xd_0__inst_mult_1_64 ),
	.shareout(Xd_0__inst_mult_1_65 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_127 (
// Equation(s):
// Xd_0__inst_mult_1_420  = SUM(( (!din_a[14] & (((din_a[15] & din_b[17])))) # (din_a[14] & (!din_b[18] $ (((!din_a[15]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_298  ) + ( Xd_0__inst_mult_1_297  ))
// Xd_0__inst_mult_1_421  = CARRY(( (!din_a[14] & (((din_a[15] & din_b[17])))) # (din_a[14] & (!din_b[18] $ (((!din_a[15]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_298  ) + ( Xd_0__inst_mult_1_297  ))
// Xd_0__inst_mult_1_422  = SHARE((din_a[14] & (din_b[18] & (din_a[15] & din_b[17]))))

	.dataa(!din_a[14]),
	.datab(!din_b[18]),
	.datac(!din_a[15]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_297 ),
	.sharein(Xd_0__inst_mult_1_298 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_420 ),
	.cout(Xd_0__inst_mult_1_421 ),
	.shareout(Xd_0__inst_mult_1_422 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_128 (
// Equation(s):
// Xd_0__inst_mult_1_425  = CARRY(( GND ) + ( Xd_0__inst_mult_6_41  ) + ( Xd_0__inst_mult_6_40  ))
// Xd_0__inst_mult_1_426  = SHARE((din_a[12] & din_b[20]))

	.dataa(!din_a[12]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_40 ),
	.sharein(Xd_0__inst_mult_6_41 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_425 ),
	.shareout(Xd_0__inst_mult_1_426 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_134 (
// Equation(s):
// Xd_0__inst_mult_4_436  = SUM(( (din_a[55] & din_b[50]) ) + ( Xd_0__inst_mult_4_422  ) + ( Xd_0__inst_mult_4_421  ))
// Xd_0__inst_mult_4_437  = CARRY(( (din_a[55] & din_b[50]) ) + ( Xd_0__inst_mult_4_422  ) + ( Xd_0__inst_mult_4_421  ))
// Xd_0__inst_mult_4_438  = SHARE((din_a[57] & din_b[49]))

	.dataa(!din_a[55]),
	.datab(!din_b[50]),
	.datac(!din_a[57]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_421 ),
	.sharein(Xd_0__inst_mult_4_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_436 ),
	.cout(Xd_0__inst_mult_4_437 ),
	.shareout(Xd_0__inst_mult_4_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_135 (
// Equation(s):
// Xd_0__inst_mult_4_440  = SUM(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_426  ) + ( Xd_0__inst_mult_4_425  ))
// Xd_0__inst_mult_4_441  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[52])))) # (din_a[54] & (!din_b[51] $ (((!din_a[53]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_426  ) + ( Xd_0__inst_mult_4_425  ))
// Xd_0__inst_mult_4_442  = SHARE((din_a[54] & (din_b[51] & (din_a[53] & din_b[52]))))

	.dataa(!din_a[54]),
	.datab(!din_b[51]),
	.datac(!din_a[53]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_425 ),
	.sharein(Xd_0__inst_mult_4_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_440 ),
	.cout(Xd_0__inst_mult_4_441 ),
	.shareout(Xd_0__inst_mult_4_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_67 (
// Equation(s):
// Xd_0__inst_mult_4_67_sumout  = SUM(( (din_a[57] & din_b[48]) ) + ( Xd_0__inst_mult_1_65  ) + ( Xd_0__inst_mult_1_64  ))
// Xd_0__inst_mult_4_68  = CARRY(( (din_a[57] & din_b[48]) ) + ( Xd_0__inst_mult_1_65  ) + ( Xd_0__inst_mult_1_64  ))
// Xd_0__inst_mult_4_69  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[48]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_64 ),
	.sharein(Xd_0__inst_mult_1_65 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_67_sumout ),
	.cout(Xd_0__inst_mult_4_68 ),
	.shareout(Xd_0__inst_mult_4_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_136 (
// Equation(s):
// Xd_0__inst_mult_4_444  = SUM(( (!din_a[51] & (((din_a[52] & din_b[53])))) # (din_a[51] & (!din_b[54] $ (((!din_a[52]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_430  ) + ( Xd_0__inst_mult_4_429  ))
// Xd_0__inst_mult_4_445  = CARRY(( (!din_a[51] & (((din_a[52] & din_b[53])))) # (din_a[51] & (!din_b[54] $ (((!din_a[52]) # (!din_b[53]))))) ) + ( Xd_0__inst_mult_4_430  ) + ( Xd_0__inst_mult_4_429  ))
// Xd_0__inst_mult_4_446  = SHARE((din_a[51] & (din_b[54] & (din_a[52] & din_b[53]))))

	.dataa(!din_a[51]),
	.datab(!din_b[54]),
	.datac(!din_a[52]),
	.datad(!din_b[53]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_429 ),
	.sharein(Xd_0__inst_mult_4_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_444 ),
	.cout(Xd_0__inst_mult_4_445 ),
	.shareout(Xd_0__inst_mult_4_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_137 (
// Equation(s):
// Xd_0__inst_mult_4_448  = SUM(( (din_a[48] & din_b[57]) ) + ( Xd_0__inst_mult_4_582  ) + ( Xd_0__inst_mult_4_581  ))
// Xd_0__inst_mult_4_449  = CARRY(( (din_a[48] & din_b[57]) ) + ( Xd_0__inst_mult_4_582  ) + ( Xd_0__inst_mult_4_581  ))
// Xd_0__inst_mult_4_450  = SHARE((din_a[48] & din_b[58]))

	.dataa(!din_a[48]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_581 ),
	.sharein(Xd_0__inst_mult_4_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_448 ),
	.cout(Xd_0__inst_mult_4_449 ),
	.shareout(Xd_0__inst_mult_4_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_133 (
// Equation(s):
// Xd_0__inst_mult_5_432  = SUM(( (din_a[67] & din_b[62]) ) + ( Xd_0__inst_mult_5_418  ) + ( Xd_0__inst_mult_5_417  ))
// Xd_0__inst_mult_5_433  = CARRY(( (din_a[67] & din_b[62]) ) + ( Xd_0__inst_mult_5_418  ) + ( Xd_0__inst_mult_5_417  ))
// Xd_0__inst_mult_5_434  = SHARE((din_a[69] & din_b[61]))

	.dataa(!din_a[67]),
	.datab(!din_b[62]),
	.datac(!din_a[69]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_417 ),
	.sharein(Xd_0__inst_mult_5_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_432 ),
	.cout(Xd_0__inst_mult_5_433 ),
	.shareout(Xd_0__inst_mult_5_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_134 (
// Equation(s):
// Xd_0__inst_mult_5_436  = SUM(( (!din_a[66] & (((din_a[65] & din_b[64])))) # (din_a[66] & (!din_b[63] $ (((!din_a[65]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_422  ) + ( Xd_0__inst_mult_5_421  ))
// Xd_0__inst_mult_5_437  = CARRY(( (!din_a[66] & (((din_a[65] & din_b[64])))) # (din_a[66] & (!din_b[63] $ (((!din_a[65]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_422  ) + ( Xd_0__inst_mult_5_421  ))
// Xd_0__inst_mult_5_438  = SHARE((din_a[66] & (din_b[63] & (din_a[65] & din_b[64]))))

	.dataa(!din_a[66]),
	.datab(!din_b[63]),
	.datac(!din_a[65]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_421 ),
	.sharein(Xd_0__inst_mult_5_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_436 ),
	.cout(Xd_0__inst_mult_5_437 ),
	.shareout(Xd_0__inst_mult_5_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_135 (
// Equation(s):
// Xd_0__inst_mult_5_440  = SUM(( (!din_a[63] & (((din_a[64] & din_b[65])))) # (din_a[63] & (!din_b[66] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_426  ) + ( Xd_0__inst_mult_5_425  ))
// Xd_0__inst_mult_5_441  = CARRY(( (!din_a[63] & (((din_a[64] & din_b[65])))) # (din_a[63] & (!din_b[66] $ (((!din_a[64]) # (!din_b[65]))))) ) + ( Xd_0__inst_mult_5_426  ) + ( Xd_0__inst_mult_5_425  ))
// Xd_0__inst_mult_5_442  = SHARE((din_a[63] & (din_b[66] & (din_a[64] & din_b[65]))))

	.dataa(!din_a[63]),
	.datab(!din_b[66]),
	.datac(!din_a[64]),
	.datad(!din_b[65]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_425 ),
	.sharein(Xd_0__inst_mult_5_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_440 ),
	.cout(Xd_0__inst_mult_5_441 ),
	.shareout(Xd_0__inst_mult_5_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_136 (
// Equation(s):
// Xd_0__inst_mult_5_444  = SUM(( (din_a[60] & din_b[69]) ) + ( Xd_0__inst_mult_5_582  ) + ( Xd_0__inst_mult_5_581  ))
// Xd_0__inst_mult_5_445  = CARRY(( (din_a[60] & din_b[69]) ) + ( Xd_0__inst_mult_5_582  ) + ( Xd_0__inst_mult_5_581  ))
// Xd_0__inst_mult_5_446  = SHARE((din_a[60] & din_b[70]))

	.dataa(!din_a[60]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_581 ),
	.sharein(Xd_0__inst_mult_5_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_444 ),
	.cout(Xd_0__inst_mult_5_445 ),
	.shareout(Xd_0__inst_mult_5_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_133 (
// Equation(s):
// Xd_0__inst_mult_2_432  = SUM(( (din_a[31] & din_b[26]) ) + ( Xd_0__inst_mult_2_418  ) + ( Xd_0__inst_mult_2_417  ))
// Xd_0__inst_mult_2_433  = CARRY(( (din_a[31] & din_b[26]) ) + ( Xd_0__inst_mult_2_418  ) + ( Xd_0__inst_mult_2_417  ))
// Xd_0__inst_mult_2_434  = SHARE((din_a[33] & din_b[25]))

	.dataa(!din_a[31]),
	.datab(!din_b[26]),
	.datac(!din_a[33]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_417 ),
	.sharein(Xd_0__inst_mult_2_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_432 ),
	.cout(Xd_0__inst_mult_2_433 ),
	.shareout(Xd_0__inst_mult_2_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_134 (
// Equation(s):
// Xd_0__inst_mult_2_436  = SUM(( (!din_a[30] & (((din_a[29] & din_b[28])))) # (din_a[30] & (!din_b[27] $ (((!din_a[29]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_422  ) + ( Xd_0__inst_mult_2_421  ))
// Xd_0__inst_mult_2_437  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[28])))) # (din_a[30] & (!din_b[27] $ (((!din_a[29]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_422  ) + ( Xd_0__inst_mult_2_421  ))
// Xd_0__inst_mult_2_438  = SHARE((din_a[30] & (din_b[27] & (din_a[29] & din_b[28]))))

	.dataa(!din_a[30]),
	.datab(!din_b[27]),
	.datac(!din_a[29]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_421 ),
	.sharein(Xd_0__inst_mult_2_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_436 ),
	.cout(Xd_0__inst_mult_2_437 ),
	.shareout(Xd_0__inst_mult_2_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_67 (
// Equation(s):
// Xd_0__inst_mult_2_67_sumout  = SUM(( (din_a[33] & din_b[24]) ) + ( Xd_0__inst_mult_3_61  ) + ( Xd_0__inst_mult_3_60  ))
// Xd_0__inst_mult_2_68  = CARRY(( (din_a[33] & din_b[24]) ) + ( Xd_0__inst_mult_3_61  ) + ( Xd_0__inst_mult_3_60  ))
// Xd_0__inst_mult_2_69  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[24]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_60 ),
	.sharein(Xd_0__inst_mult_3_61 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_67_sumout ),
	.cout(Xd_0__inst_mult_2_68 ),
	.shareout(Xd_0__inst_mult_2_69 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_135 (
// Equation(s):
// Xd_0__inst_mult_2_440  = SUM(( (!din_a[27] & (((din_a[28] & din_b[29])))) # (din_a[27] & (!din_b[30] $ (((!din_a[28]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_426  ) + ( Xd_0__inst_mult_2_425  ))
// Xd_0__inst_mult_2_441  = CARRY(( (!din_a[27] & (((din_a[28] & din_b[29])))) # (din_a[27] & (!din_b[30] $ (((!din_a[28]) # (!din_b[29]))))) ) + ( Xd_0__inst_mult_2_426  ) + ( Xd_0__inst_mult_2_425  ))
// Xd_0__inst_mult_2_442  = SHARE((din_a[27] & (din_b[30] & (din_a[28] & din_b[29]))))

	.dataa(!din_a[27]),
	.datab(!din_b[30]),
	.datac(!din_a[28]),
	.datad(!din_b[29]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_425 ),
	.sharein(Xd_0__inst_mult_2_426 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_440 ),
	.cout(Xd_0__inst_mult_2_441 ),
	.shareout(Xd_0__inst_mult_2_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_136 (
// Equation(s):
// Xd_0__inst_mult_2_444  = SUM(( (din_a[24] & din_b[33]) ) + ( Xd_0__inst_mult_2_582  ) + ( Xd_0__inst_mult_2_581  ))
// Xd_0__inst_mult_2_445  = CARRY(( (din_a[24] & din_b[33]) ) + ( Xd_0__inst_mult_2_582  ) + ( Xd_0__inst_mult_2_581  ))
// Xd_0__inst_mult_2_446  = SHARE((din_a[24] & din_b[34]))

	.dataa(!din_a[24]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_581 ),
	.sharein(Xd_0__inst_mult_2_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_444 ),
	.cout(Xd_0__inst_mult_2_445 ),
	.shareout(Xd_0__inst_mult_2_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_140 (
// Equation(s):
// Xd_0__inst_mult_3_472  = SUM(( (din_a[43] & din_b[38]) ) + ( Xd_0__inst_mult_3_458  ) + ( Xd_0__inst_mult_3_457  ))
// Xd_0__inst_mult_3_473  = CARRY(( (din_a[43] & din_b[38]) ) + ( Xd_0__inst_mult_3_458  ) + ( Xd_0__inst_mult_3_457  ))
// Xd_0__inst_mult_3_474  = SHARE((din_a[45] & din_b[37]))

	.dataa(!din_a[43]),
	.datab(!din_b[38]),
	.datac(!din_a[45]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_457 ),
	.sharein(Xd_0__inst_mult_3_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_472 ),
	.cout(Xd_0__inst_mult_3_473 ),
	.shareout(Xd_0__inst_mult_3_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_141 (
// Equation(s):
// Xd_0__inst_mult_3_476  = SUM(( (!din_a[42] & (((din_a[41] & din_b[40])))) # (din_a[42] & (!din_b[39] $ (((!din_a[41]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_462  ) + ( Xd_0__inst_mult_3_461  ))
// Xd_0__inst_mult_3_477  = CARRY(( (!din_a[42] & (((din_a[41] & din_b[40])))) # (din_a[42] & (!din_b[39] $ (((!din_a[41]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_462  ) + ( Xd_0__inst_mult_3_461  ))
// Xd_0__inst_mult_3_478  = SHARE((din_a[42] & (din_b[39] & (din_a[41] & din_b[40]))))

	.dataa(!din_a[42]),
	.datab(!din_b[39]),
	.datac(!din_a[41]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_461 ),
	.sharein(Xd_0__inst_mult_3_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_476 ),
	.cout(Xd_0__inst_mult_3_477 ),
	.shareout(Xd_0__inst_mult_3_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_142 (
// Equation(s):
// Xd_0__inst_mult_3_480  = SUM(( (!din_a[39] & (((din_a[40] & din_b[41])))) # (din_a[39] & (!din_b[42] $ (((!din_a[40]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_466  ) + ( Xd_0__inst_mult_3_465  ))
// Xd_0__inst_mult_3_481  = CARRY(( (!din_a[39] & (((din_a[40] & din_b[41])))) # (din_a[39] & (!din_b[42] $ (((!din_a[40]) # (!din_b[41]))))) ) + ( Xd_0__inst_mult_3_466  ) + ( Xd_0__inst_mult_3_465  ))
// Xd_0__inst_mult_3_482  = SHARE((din_a[39] & (din_b[42] & (din_a[40] & din_b[41]))))

	.dataa(!din_a[39]),
	.datab(!din_b[42]),
	.datac(!din_a[40]),
	.datad(!din_b[41]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_465 ),
	.sharein(Xd_0__inst_mult_3_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_480 ),
	.cout(Xd_0__inst_mult_3_481 ),
	.shareout(Xd_0__inst_mult_3_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_143 (
// Equation(s):
// Xd_0__inst_mult_3_484  = SUM(( (din_a[36] & din_b[45]) ) + ( Xd_0__inst_mult_3_574  ) + ( Xd_0__inst_mult_3_573  ))
// Xd_0__inst_mult_3_485  = CARRY(( (din_a[36] & din_b[45]) ) + ( Xd_0__inst_mult_3_574  ) + ( Xd_0__inst_mult_3_573  ))
// Xd_0__inst_mult_3_486  = SHARE((din_a[36] & din_b[46]))

	.dataa(!din_a[36]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_573 ),
	.sharein(Xd_0__inst_mult_3_574 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_484 ),
	.cout(Xd_0__inst_mult_3_485 ),
	.shareout(Xd_0__inst_mult_3_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_133 (
// Equation(s):
// Xd_0__inst_mult_0_444  = SUM(( (din_a[7] & din_b[2]) ) + ( Xd_0__inst_mult_0_430  ) + ( Xd_0__inst_mult_0_429  ))
// Xd_0__inst_mult_0_445  = CARRY(( (din_a[7] & din_b[2]) ) + ( Xd_0__inst_mult_0_430  ) + ( Xd_0__inst_mult_0_429  ))
// Xd_0__inst_mult_0_446  = SHARE((din_a[9] & din_b[1]))

	.dataa(!din_a[7]),
	.datab(!din_b[2]),
	.datac(!din_a[9]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_429 ),
	.sharein(Xd_0__inst_mult_0_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_444 ),
	.cout(Xd_0__inst_mult_0_445 ),
	.shareout(Xd_0__inst_mult_0_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_134 (
// Equation(s):
// Xd_0__inst_mult_0_448  = SUM(( (!din_a[6] & (((din_a[5] & din_b[4])))) # (din_a[6] & (!din_b[3] $ (((!din_a[5]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_434  ) + ( Xd_0__inst_mult_0_433  ))
// Xd_0__inst_mult_0_449  = CARRY(( (!din_a[6] & (((din_a[5] & din_b[4])))) # (din_a[6] & (!din_b[3] $ (((!din_a[5]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_434  ) + ( Xd_0__inst_mult_0_433  ))
// Xd_0__inst_mult_0_450  = SHARE((din_a[6] & (din_b[3] & (din_a[5] & din_b[4]))))

	.dataa(!din_a[6]),
	.datab(!din_b[3]),
	.datac(!din_a[5]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_433 ),
	.sharein(Xd_0__inst_mult_0_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_448 ),
	.cout(Xd_0__inst_mult_0_449 ),
	.shareout(Xd_0__inst_mult_0_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_135 (
// Equation(s):
// Xd_0__inst_mult_0_452  = SUM(( (!din_a[3] & (((din_a[4] & din_b[5])))) # (din_a[3] & (!din_b[6] $ (((!din_a[4]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_438  ) + ( Xd_0__inst_mult_0_437  ))
// Xd_0__inst_mult_0_453  = CARRY(( (!din_a[3] & (((din_a[4] & din_b[5])))) # (din_a[3] & (!din_b[6] $ (((!din_a[4]) # (!din_b[5]))))) ) + ( Xd_0__inst_mult_0_438  ) + ( Xd_0__inst_mult_0_437  ))
// Xd_0__inst_mult_0_454  = SHARE((din_a[3] & (din_b[6] & (din_a[4] & din_b[5]))))

	.dataa(!din_a[3]),
	.datab(!din_b[6]),
	.datac(!din_a[4]),
	.datad(!din_b[5]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_437 ),
	.sharein(Xd_0__inst_mult_0_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_452 ),
	.cout(Xd_0__inst_mult_0_453 ),
	.shareout(Xd_0__inst_mult_0_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_136 (
// Equation(s):
// Xd_0__inst_mult_0_456  = SUM(( (din_a[0] & din_b[9]) ) + ( Xd_0__inst_mult_0_578  ) + ( Xd_0__inst_mult_0_577  ))
// Xd_0__inst_mult_0_457  = CARRY(( (din_a[0] & din_b[9]) ) + ( Xd_0__inst_mult_0_578  ) + ( Xd_0__inst_mult_0_577  ))
// Xd_0__inst_mult_0_458  = SHARE((din_a[0] & din_b[10]))

	.dataa(!din_a[0]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_577 ),
	.sharein(Xd_0__inst_mult_0_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_456 ),
	.cout(Xd_0__inst_mult_0_457 ),
	.shareout(Xd_0__inst_mult_0_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_129 (
// Equation(s):
// Xd_0__inst_mult_1_428  = SUM(( (din_a[19] & din_b[14]) ) + ( Xd_0__inst_mult_1_414  ) + ( Xd_0__inst_mult_1_413  ))
// Xd_0__inst_mult_1_429  = CARRY(( (din_a[19] & din_b[14]) ) + ( Xd_0__inst_mult_1_414  ) + ( Xd_0__inst_mult_1_413  ))
// Xd_0__inst_mult_1_430  = SHARE((din_a[21] & din_b[13]))

	.dataa(!din_a[19]),
	.datab(!din_b[14]),
	.datac(!din_a[21]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_413 ),
	.sharein(Xd_0__inst_mult_1_414 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_428 ),
	.cout(Xd_0__inst_mult_1_429 ),
	.shareout(Xd_0__inst_mult_1_430 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_130 (
// Equation(s):
// Xd_0__inst_mult_1_432  = SUM(( (!din_a[18] & (((din_a[17] & din_b[16])))) # (din_a[18] & (!din_b[15] $ (((!din_a[17]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_418  ) + ( Xd_0__inst_mult_1_417  ))
// Xd_0__inst_mult_1_433  = CARRY(( (!din_a[18] & (((din_a[17] & din_b[16])))) # (din_a[18] & (!din_b[15] $ (((!din_a[17]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_418  ) + ( Xd_0__inst_mult_1_417  ))
// Xd_0__inst_mult_1_434  = SHARE((din_a[18] & (din_b[15] & (din_a[17] & din_b[16]))))

	.dataa(!din_a[18]),
	.datab(!din_b[15]),
	.datac(!din_a[17]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_417 ),
	.sharein(Xd_0__inst_mult_1_418 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_432 ),
	.cout(Xd_0__inst_mult_1_433 ),
	.shareout(Xd_0__inst_mult_1_434 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_131 (
// Equation(s):
// Xd_0__inst_mult_1_436  = SUM(( (!din_a[15] & (((din_a[16] & din_b[17])))) # (din_a[15] & (!din_b[18] $ (((!din_a[16]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_422  ) + ( Xd_0__inst_mult_1_421  ))
// Xd_0__inst_mult_1_437  = CARRY(( (!din_a[15] & (((din_a[16] & din_b[17])))) # (din_a[15] & (!din_b[18] $ (((!din_a[16]) # (!din_b[17]))))) ) + ( Xd_0__inst_mult_1_422  ) + ( Xd_0__inst_mult_1_421  ))
// Xd_0__inst_mult_1_438  = SHARE((din_a[15] & (din_b[18] & (din_a[16] & din_b[17]))))

	.dataa(!din_a[15]),
	.datab(!din_b[18]),
	.datac(!din_a[16]),
	.datad(!din_b[17]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_421 ),
	.sharein(Xd_0__inst_mult_1_422 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_436 ),
	.cout(Xd_0__inst_mult_1_437 ),
	.shareout(Xd_0__inst_mult_1_438 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_132 (
// Equation(s):
// Xd_0__inst_mult_1_440  = SUM(( (din_a[12] & din_b[21]) ) + ( Xd_0__inst_mult_1_578  ) + ( Xd_0__inst_mult_1_577  ))
// Xd_0__inst_mult_1_441  = CARRY(( (din_a[12] & din_b[21]) ) + ( Xd_0__inst_mult_1_578  ) + ( Xd_0__inst_mult_1_577  ))
// Xd_0__inst_mult_1_442  = SHARE((din_a[12] & din_b[22]))

	.dataa(!din_a[12]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_577 ),
	.sharein(Xd_0__inst_mult_1_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_440 ),
	.cout(Xd_0__inst_mult_1_441 ),
	.shareout(Xd_0__inst_mult_1_442 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_6_169 (
// Equation(s):
// Xd_0__inst_mult_6_577  = CARRY(( (din_a[74] & din_b[79]) ) + ( Xd_0__inst_mult_6_586  ) + ( Xd_0__inst_mult_6_585  ))
// Xd_0__inst_mult_6_578  = SHARE((din_a[73] & din_b[80]))

	.dataa(!din_a[74]),
	.datab(!din_b[79]),
	.datac(!din_a[73]),
	.datad(!din_b[80]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_6_585 ),
	.sharein(Xd_0__inst_mult_6_586 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_577 ),
	.shareout(Xd_0__inst_mult_6_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_7_169 (
// Equation(s):
// Xd_0__inst_mult_7_577  = CARRY(( (din_a[86] & din_b[91]) ) + ( Xd_0__inst_mult_7_586  ) + ( Xd_0__inst_mult_7_585  ))
// Xd_0__inst_mult_7_578  = SHARE((din_a[85] & din_b[92]))

	.dataa(!din_a[86]),
	.datab(!din_b[91]),
	.datac(!din_a[85]),
	.datad(!din_b[92]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_7_585 ),
	.sharein(Xd_0__inst_mult_7_586 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_577 ),
	.shareout(Xd_0__inst_mult_7_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_138 (
// Equation(s):
// Xd_0__inst_mult_4_452  = SUM(( (din_a[56] & din_b[50]) ) + ( Xd_0__inst_mult_4_438  ) + ( Xd_0__inst_mult_4_437  ))
// Xd_0__inst_mult_4_453  = CARRY(( (din_a[56] & din_b[50]) ) + ( Xd_0__inst_mult_4_438  ) + ( Xd_0__inst_mult_4_437  ))
// Xd_0__inst_mult_4_454  = SHARE((din_a[58] & din_b[49]))

	.dataa(!din_a[56]),
	.datab(!din_b[50]),
	.datac(!din_a[58]),
	.datad(!din_b[49]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_437 ),
	.sharein(Xd_0__inst_mult_4_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_452 ),
	.cout(Xd_0__inst_mult_4_453 ),
	.shareout(Xd_0__inst_mult_4_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_139 (
// Equation(s):
// Xd_0__inst_mult_4_456  = SUM(( (!din_a[55] & (((din_a[54] & din_b[52])))) # (din_a[55] & (!din_b[51] $ (((!din_a[54]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_442  ) + ( Xd_0__inst_mult_4_441  ))
// Xd_0__inst_mult_4_457  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[52])))) # (din_a[55] & (!din_b[51] $ (((!din_a[54]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_442  ) + ( Xd_0__inst_mult_4_441  ))
// Xd_0__inst_mult_4_458  = SHARE((din_a[55] & (din_b[51] & (din_a[54] & din_b[52]))))

	.dataa(!din_a[55]),
	.datab(!din_b[51]),
	.datac(!din_a[54]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_441 ),
	.sharein(Xd_0__inst_mult_4_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_456 ),
	.cout(Xd_0__inst_mult_4_457 ),
	.shareout(Xd_0__inst_mult_4_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_140 (
// Equation(s):
// Xd_0__inst_mult_4_460  = SUM(( (din_a[53] & din_b[53]) ) + ( Xd_0__inst_mult_4_446  ) + ( Xd_0__inst_mult_4_445  ))
// Xd_0__inst_mult_4_461  = CARRY(( (din_a[53] & din_b[53]) ) + ( Xd_0__inst_mult_4_446  ) + ( Xd_0__inst_mult_4_445  ))
// Xd_0__inst_mult_4_462  = SHARE((din_a[53] & din_b[54]))

	.dataa(!din_a[53]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_445 ),
	.sharein(Xd_0__inst_mult_4_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_460 ),
	.cout(Xd_0__inst_mult_4_461 ),
	.shareout(Xd_0__inst_mult_4_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_141 (
// Equation(s):
// Xd_0__inst_mult_4_464  = SUM(( (din_a[49] & din_b[57]) ) + ( Xd_0__inst_mult_4_450  ) + ( Xd_0__inst_mult_4_449  ))
// Xd_0__inst_mult_4_465  = CARRY(( (din_a[49] & din_b[57]) ) + ( Xd_0__inst_mult_4_450  ) + ( Xd_0__inst_mult_4_449  ))
// Xd_0__inst_mult_4_466  = SHARE((din_a[49] & din_b[58]))

	.dataa(!din_a[49]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_449 ),
	.sharein(Xd_0__inst_mult_4_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_464 ),
	.cout(Xd_0__inst_mult_4_465 ),
	.shareout(Xd_0__inst_mult_4_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_142 (
// Equation(s):
// Xd_0__inst_mult_4_468  = SUM(( (!din_a[51] & (((din_a[50] & din_b[56])))) # (din_a[51] & (!din_b[55] $ (((!din_a[50]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_586  ) + ( Xd_0__inst_mult_4_585  ))
// Xd_0__inst_mult_4_469  = CARRY(( (!din_a[51] & (((din_a[50] & din_b[56])))) # (din_a[51] & (!din_b[55] $ (((!din_a[50]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_586  ) + ( Xd_0__inst_mult_4_585  ))
// Xd_0__inst_mult_4_470  = SHARE((din_a[51] & (din_b[55] & (din_a[50] & din_b[56]))))

	.dataa(!din_a[51]),
	.datab(!din_b[55]),
	.datac(!din_a[50]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_585 ),
	.sharein(Xd_0__inst_mult_4_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_468 ),
	.cout(Xd_0__inst_mult_4_469 ),
	.shareout(Xd_0__inst_mult_4_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_137 (
// Equation(s):
// Xd_0__inst_mult_5_448  = SUM(( (din_a[68] & din_b[62]) ) + ( Xd_0__inst_mult_5_434  ) + ( Xd_0__inst_mult_5_433  ))
// Xd_0__inst_mult_5_449  = CARRY(( (din_a[68] & din_b[62]) ) + ( Xd_0__inst_mult_5_434  ) + ( Xd_0__inst_mult_5_433  ))
// Xd_0__inst_mult_5_450  = SHARE((din_a[70] & din_b[61]))

	.dataa(!din_a[68]),
	.datab(!din_b[62]),
	.datac(!din_a[70]),
	.datad(!din_b[61]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_433 ),
	.sharein(Xd_0__inst_mult_5_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_448 ),
	.cout(Xd_0__inst_mult_5_449 ),
	.shareout(Xd_0__inst_mult_5_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_138 (
// Equation(s):
// Xd_0__inst_mult_5_452  = SUM(( (!din_a[67] & (((din_a[66] & din_b[64])))) # (din_a[67] & (!din_b[63] $ (((!din_a[66]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_438  ) + ( Xd_0__inst_mult_5_437  ))
// Xd_0__inst_mult_5_453  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[64])))) # (din_a[67] & (!din_b[63] $ (((!din_a[66]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_438  ) + ( Xd_0__inst_mult_5_437  ))
// Xd_0__inst_mult_5_454  = SHARE((din_a[67] & (din_b[63] & (din_a[66] & din_b[64]))))

	.dataa(!din_a[67]),
	.datab(!din_b[63]),
	.datac(!din_a[66]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_437 ),
	.sharein(Xd_0__inst_mult_5_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_452 ),
	.cout(Xd_0__inst_mult_5_453 ),
	.shareout(Xd_0__inst_mult_5_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_139 (
// Equation(s):
// Xd_0__inst_mult_5_456  = SUM(( (din_a[65] & din_b[65]) ) + ( Xd_0__inst_mult_5_442  ) + ( Xd_0__inst_mult_5_441  ))
// Xd_0__inst_mult_5_457  = CARRY(( (din_a[65] & din_b[65]) ) + ( Xd_0__inst_mult_5_442  ) + ( Xd_0__inst_mult_5_441  ))
// Xd_0__inst_mult_5_458  = SHARE((din_a[65] & din_b[66]))

	.dataa(!din_a[65]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_441 ),
	.sharein(Xd_0__inst_mult_5_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_456 ),
	.cout(Xd_0__inst_mult_5_457 ),
	.shareout(Xd_0__inst_mult_5_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_140 (
// Equation(s):
// Xd_0__inst_mult_5_460  = SUM(( (din_a[61] & din_b[69]) ) + ( Xd_0__inst_mult_5_446  ) + ( Xd_0__inst_mult_5_445  ))
// Xd_0__inst_mult_5_461  = CARRY(( (din_a[61] & din_b[69]) ) + ( Xd_0__inst_mult_5_446  ) + ( Xd_0__inst_mult_5_445  ))
// Xd_0__inst_mult_5_462  = SHARE((din_a[61] & din_b[70]))

	.dataa(!din_a[61]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_445 ),
	.sharein(Xd_0__inst_mult_5_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_460 ),
	.cout(Xd_0__inst_mult_5_461 ),
	.shareout(Xd_0__inst_mult_5_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_141 (
// Equation(s):
// Xd_0__inst_mult_5_464  = SUM(( (!din_a[63] & (((din_a[62] & din_b[68])))) # (din_a[63] & (!din_b[67] $ (((!din_a[62]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_586  ) + ( Xd_0__inst_mult_5_585  ))
// Xd_0__inst_mult_5_465  = CARRY(( (!din_a[63] & (((din_a[62] & din_b[68])))) # (din_a[63] & (!din_b[67] $ (((!din_a[62]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_586  ) + ( Xd_0__inst_mult_5_585  ))
// Xd_0__inst_mult_5_466  = SHARE((din_a[63] & (din_b[67] & (din_a[62] & din_b[68]))))

	.dataa(!din_a[63]),
	.datab(!din_b[67]),
	.datac(!din_a[62]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_585 ),
	.sharein(Xd_0__inst_mult_5_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_464 ),
	.cout(Xd_0__inst_mult_5_465 ),
	.shareout(Xd_0__inst_mult_5_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_137 (
// Equation(s):
// Xd_0__inst_mult_2_448  = SUM(( (din_a[32] & din_b[26]) ) + ( Xd_0__inst_mult_2_434  ) + ( Xd_0__inst_mult_2_433  ))
// Xd_0__inst_mult_2_449  = CARRY(( (din_a[32] & din_b[26]) ) + ( Xd_0__inst_mult_2_434  ) + ( Xd_0__inst_mult_2_433  ))
// Xd_0__inst_mult_2_450  = SHARE((din_a[34] & din_b[25]))

	.dataa(!din_a[32]),
	.datab(!din_b[26]),
	.datac(!din_a[34]),
	.datad(!din_b[25]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_433 ),
	.sharein(Xd_0__inst_mult_2_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_448 ),
	.cout(Xd_0__inst_mult_2_449 ),
	.shareout(Xd_0__inst_mult_2_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_138 (
// Equation(s):
// Xd_0__inst_mult_2_452  = SUM(( (!din_a[31] & (((din_a[30] & din_b[28])))) # (din_a[31] & (!din_b[27] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_438  ) + ( Xd_0__inst_mult_2_437  ))
// Xd_0__inst_mult_2_453  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[28])))) # (din_a[31] & (!din_b[27] $ (((!din_a[30]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_438  ) + ( Xd_0__inst_mult_2_437  ))
// Xd_0__inst_mult_2_454  = SHARE((din_a[31] & (din_b[27] & (din_a[30] & din_b[28]))))

	.dataa(!din_a[31]),
	.datab(!din_b[27]),
	.datac(!din_a[30]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_437 ),
	.sharein(Xd_0__inst_mult_2_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_452 ),
	.cout(Xd_0__inst_mult_2_453 ),
	.shareout(Xd_0__inst_mult_2_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_139 (
// Equation(s):
// Xd_0__inst_mult_2_456  = SUM(( (din_a[29] & din_b[29]) ) + ( Xd_0__inst_mult_2_442  ) + ( Xd_0__inst_mult_2_441  ))
// Xd_0__inst_mult_2_457  = CARRY(( (din_a[29] & din_b[29]) ) + ( Xd_0__inst_mult_2_442  ) + ( Xd_0__inst_mult_2_441  ))
// Xd_0__inst_mult_2_458  = SHARE((din_a[29] & din_b[30]))

	.dataa(!din_a[29]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_441 ),
	.sharein(Xd_0__inst_mult_2_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_456 ),
	.cout(Xd_0__inst_mult_2_457 ),
	.shareout(Xd_0__inst_mult_2_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_140 (
// Equation(s):
// Xd_0__inst_mult_2_460  = SUM(( (din_a[25] & din_b[33]) ) + ( Xd_0__inst_mult_2_446  ) + ( Xd_0__inst_mult_2_445  ))
// Xd_0__inst_mult_2_461  = CARRY(( (din_a[25] & din_b[33]) ) + ( Xd_0__inst_mult_2_446  ) + ( Xd_0__inst_mult_2_445  ))
// Xd_0__inst_mult_2_462  = SHARE((din_a[25] & din_b[34]))

	.dataa(!din_a[25]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_445 ),
	.sharein(Xd_0__inst_mult_2_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_460 ),
	.cout(Xd_0__inst_mult_2_461 ),
	.shareout(Xd_0__inst_mult_2_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_141 (
// Equation(s):
// Xd_0__inst_mult_2_464  = SUM(( (!din_a[27] & (((din_a[26] & din_b[32])))) # (din_a[27] & (!din_b[31] $ (((!din_a[26]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_586  ) + ( Xd_0__inst_mult_2_585  ))
// Xd_0__inst_mult_2_465  = CARRY(( (!din_a[27] & (((din_a[26] & din_b[32])))) # (din_a[27] & (!din_b[31] $ (((!din_a[26]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_586  ) + ( Xd_0__inst_mult_2_585  ))
// Xd_0__inst_mult_2_466  = SHARE((din_a[27] & (din_b[31] & (din_a[26] & din_b[32]))))

	.dataa(!din_a[27]),
	.datab(!din_b[31]),
	.datac(!din_a[26]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_585 ),
	.sharein(Xd_0__inst_mult_2_586 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_464 ),
	.cout(Xd_0__inst_mult_2_465 ),
	.shareout(Xd_0__inst_mult_2_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_144 (
// Equation(s):
// Xd_0__inst_mult_3_488  = SUM(( (din_a[44] & din_b[38]) ) + ( Xd_0__inst_mult_3_474  ) + ( Xd_0__inst_mult_3_473  ))
// Xd_0__inst_mult_3_489  = CARRY(( (din_a[44] & din_b[38]) ) + ( Xd_0__inst_mult_3_474  ) + ( Xd_0__inst_mult_3_473  ))
// Xd_0__inst_mult_3_490  = SHARE((din_a[46] & din_b[37]))

	.dataa(!din_a[44]),
	.datab(!din_b[38]),
	.datac(!din_a[46]),
	.datad(!din_b[37]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_473 ),
	.sharein(Xd_0__inst_mult_3_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_488 ),
	.cout(Xd_0__inst_mult_3_489 ),
	.shareout(Xd_0__inst_mult_3_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_145 (
// Equation(s):
// Xd_0__inst_mult_3_492  = SUM(( (!din_a[43] & (((din_a[42] & din_b[40])))) # (din_a[43] & (!din_b[39] $ (((!din_a[42]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_478  ) + ( Xd_0__inst_mult_3_477  ))
// Xd_0__inst_mult_3_493  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[40])))) # (din_a[43] & (!din_b[39] $ (((!din_a[42]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_478  ) + ( Xd_0__inst_mult_3_477  ))
// Xd_0__inst_mult_3_494  = SHARE((din_a[43] & (din_b[39] & (din_a[42] & din_b[40]))))

	.dataa(!din_a[43]),
	.datab(!din_b[39]),
	.datac(!din_a[42]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_477 ),
	.sharein(Xd_0__inst_mult_3_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_492 ),
	.cout(Xd_0__inst_mult_3_493 ),
	.shareout(Xd_0__inst_mult_3_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_146 (
// Equation(s):
// Xd_0__inst_mult_3_496  = SUM(( (din_a[41] & din_b[41]) ) + ( Xd_0__inst_mult_3_482  ) + ( Xd_0__inst_mult_3_481  ))
// Xd_0__inst_mult_3_497  = CARRY(( (din_a[41] & din_b[41]) ) + ( Xd_0__inst_mult_3_482  ) + ( Xd_0__inst_mult_3_481  ))
// Xd_0__inst_mult_3_498  = SHARE((din_a[41] & din_b[42]))

	.dataa(!din_a[41]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_481 ),
	.sharein(Xd_0__inst_mult_3_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_496 ),
	.cout(Xd_0__inst_mult_3_497 ),
	.shareout(Xd_0__inst_mult_3_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_147 (
// Equation(s):
// Xd_0__inst_mult_3_500  = SUM(( (din_a[37] & din_b[45]) ) + ( Xd_0__inst_mult_3_486  ) + ( Xd_0__inst_mult_3_485  ))
// Xd_0__inst_mult_3_501  = CARRY(( (din_a[37] & din_b[45]) ) + ( Xd_0__inst_mult_3_486  ) + ( Xd_0__inst_mult_3_485  ))
// Xd_0__inst_mult_3_502  = SHARE((din_a[37] & din_b[46]))

	.dataa(!din_a[37]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_485 ),
	.sharein(Xd_0__inst_mult_3_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_500 ),
	.cout(Xd_0__inst_mult_3_501 ),
	.shareout(Xd_0__inst_mult_3_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_148 (
// Equation(s):
// Xd_0__inst_mult_3_504  = SUM(( (!din_a[39] & (((din_a[38] & din_b[44])))) # (din_a[39] & (!din_b[43] $ (((!din_a[38]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_578  ) + ( Xd_0__inst_mult_3_577  ))
// Xd_0__inst_mult_3_505  = CARRY(( (!din_a[39] & (((din_a[38] & din_b[44])))) # (din_a[39] & (!din_b[43] $ (((!din_a[38]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_578  ) + ( Xd_0__inst_mult_3_577  ))
// Xd_0__inst_mult_3_506  = SHARE((din_a[39] & (din_b[43] & (din_a[38] & din_b[44]))))

	.dataa(!din_a[39]),
	.datab(!din_b[43]),
	.datac(!din_a[38]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_577 ),
	.sharein(Xd_0__inst_mult_3_578 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_504 ),
	.cout(Xd_0__inst_mult_3_505 ),
	.shareout(Xd_0__inst_mult_3_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_137 (
// Equation(s):
// Xd_0__inst_mult_0_460  = SUM(( (din_a[8] & din_b[2]) ) + ( Xd_0__inst_mult_0_446  ) + ( Xd_0__inst_mult_0_445  ))
// Xd_0__inst_mult_0_461  = CARRY(( (din_a[8] & din_b[2]) ) + ( Xd_0__inst_mult_0_446  ) + ( Xd_0__inst_mult_0_445  ))
// Xd_0__inst_mult_0_462  = SHARE((din_a[10] & din_b[1]))

	.dataa(!din_a[8]),
	.datab(!din_b[2]),
	.datac(!din_a[10]),
	.datad(!din_b[1]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_445 ),
	.sharein(Xd_0__inst_mult_0_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_460 ),
	.cout(Xd_0__inst_mult_0_461 ),
	.shareout(Xd_0__inst_mult_0_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_138 (
// Equation(s):
// Xd_0__inst_mult_0_464  = SUM(( (!din_a[7] & (((din_a[6] & din_b[4])))) # (din_a[7] & (!din_b[3] $ (((!din_a[6]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_450  ) + ( Xd_0__inst_mult_0_449  ))
// Xd_0__inst_mult_0_465  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[4])))) # (din_a[7] & (!din_b[3] $ (((!din_a[6]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_450  ) + ( Xd_0__inst_mult_0_449  ))
// Xd_0__inst_mult_0_466  = SHARE((din_a[7] & (din_b[3] & (din_a[6] & din_b[4]))))

	.dataa(!din_a[7]),
	.datab(!din_b[3]),
	.datac(!din_a[6]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_449 ),
	.sharein(Xd_0__inst_mult_0_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_464 ),
	.cout(Xd_0__inst_mult_0_465 ),
	.shareout(Xd_0__inst_mult_0_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_139 (
// Equation(s):
// Xd_0__inst_mult_0_468  = SUM(( (din_a[5] & din_b[5]) ) + ( Xd_0__inst_mult_0_454  ) + ( Xd_0__inst_mult_0_453  ))
// Xd_0__inst_mult_0_469  = CARRY(( (din_a[5] & din_b[5]) ) + ( Xd_0__inst_mult_0_454  ) + ( Xd_0__inst_mult_0_453  ))
// Xd_0__inst_mult_0_470  = SHARE((din_a[5] & din_b[6]))

	.dataa(!din_a[5]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_453 ),
	.sharein(Xd_0__inst_mult_0_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_468 ),
	.cout(Xd_0__inst_mult_0_469 ),
	.shareout(Xd_0__inst_mult_0_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_140 (
// Equation(s):
// Xd_0__inst_mult_0_472  = SUM(( (din_a[1] & din_b[9]) ) + ( Xd_0__inst_mult_0_458  ) + ( Xd_0__inst_mult_0_457  ))
// Xd_0__inst_mult_0_473  = CARRY(( (din_a[1] & din_b[9]) ) + ( Xd_0__inst_mult_0_458  ) + ( Xd_0__inst_mult_0_457  ))
// Xd_0__inst_mult_0_474  = SHARE((din_a[1] & din_b[10]))

	.dataa(!din_a[1]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_457 ),
	.sharein(Xd_0__inst_mult_0_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_472 ),
	.cout(Xd_0__inst_mult_0_473 ),
	.shareout(Xd_0__inst_mult_0_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_141 (
// Equation(s):
// Xd_0__inst_mult_0_476  = SUM(( (!din_a[3] & (((din_a[2] & din_b[8])))) # (din_a[3] & (!din_b[7] $ (((!din_a[2]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_582  ) + ( Xd_0__inst_mult_0_581  ))
// Xd_0__inst_mult_0_477  = CARRY(( (!din_a[3] & (((din_a[2] & din_b[8])))) # (din_a[3] & (!din_b[7] $ (((!din_a[2]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_582  ) + ( Xd_0__inst_mult_0_581  ))
// Xd_0__inst_mult_0_478  = SHARE((din_a[3] & (din_b[7] & (din_a[2] & din_b[8]))))

	.dataa(!din_a[3]),
	.datab(!din_b[7]),
	.datac(!din_a[2]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_581 ),
	.sharein(Xd_0__inst_mult_0_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_476 ),
	.cout(Xd_0__inst_mult_0_477 ),
	.shareout(Xd_0__inst_mult_0_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_133 (
// Equation(s):
// Xd_0__inst_mult_1_444  = SUM(( (din_a[20] & din_b[14]) ) + ( Xd_0__inst_mult_1_430  ) + ( Xd_0__inst_mult_1_429  ))
// Xd_0__inst_mult_1_445  = CARRY(( (din_a[20] & din_b[14]) ) + ( Xd_0__inst_mult_1_430  ) + ( Xd_0__inst_mult_1_429  ))
// Xd_0__inst_mult_1_446  = SHARE((din_a[22] & din_b[13]))

	.dataa(!din_a[20]),
	.datab(!din_b[14]),
	.datac(!din_a[22]),
	.datad(!din_b[13]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_429 ),
	.sharein(Xd_0__inst_mult_1_430 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_444 ),
	.cout(Xd_0__inst_mult_1_445 ),
	.shareout(Xd_0__inst_mult_1_446 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_134 (
// Equation(s):
// Xd_0__inst_mult_1_448  = SUM(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_434  ) + ( Xd_0__inst_mult_1_433  ))
// Xd_0__inst_mult_1_449  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[16])))) # (din_a[19] & (!din_b[15] $ (((!din_a[18]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_434  ) + ( Xd_0__inst_mult_1_433  ))
// Xd_0__inst_mult_1_450  = SHARE((din_a[19] & (din_b[15] & (din_a[18] & din_b[16]))))

	.dataa(!din_a[19]),
	.datab(!din_b[15]),
	.datac(!din_a[18]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_433 ),
	.sharein(Xd_0__inst_mult_1_434 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_448 ),
	.cout(Xd_0__inst_mult_1_449 ),
	.shareout(Xd_0__inst_mult_1_450 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_135 (
// Equation(s):
// Xd_0__inst_mult_1_452  = SUM(( (din_a[17] & din_b[17]) ) + ( Xd_0__inst_mult_1_438  ) + ( Xd_0__inst_mult_1_437  ))
// Xd_0__inst_mult_1_453  = CARRY(( (din_a[17] & din_b[17]) ) + ( Xd_0__inst_mult_1_438  ) + ( Xd_0__inst_mult_1_437  ))
// Xd_0__inst_mult_1_454  = SHARE((din_a[17] & din_b[18]))

	.dataa(!din_a[17]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_437 ),
	.sharein(Xd_0__inst_mult_1_438 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_452 ),
	.cout(Xd_0__inst_mult_1_453 ),
	.shareout(Xd_0__inst_mult_1_454 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_136 (
// Equation(s):
// Xd_0__inst_mult_1_456  = SUM(( (din_a[13] & din_b[21]) ) + ( Xd_0__inst_mult_1_442  ) + ( Xd_0__inst_mult_1_441  ))
// Xd_0__inst_mult_1_457  = CARRY(( (din_a[13] & din_b[21]) ) + ( Xd_0__inst_mult_1_442  ) + ( Xd_0__inst_mult_1_441  ))
// Xd_0__inst_mult_1_458  = SHARE((din_a[13] & din_b[22]))

	.dataa(!din_a[13]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_441 ),
	.sharein(Xd_0__inst_mult_1_442 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_456 ),
	.cout(Xd_0__inst_mult_1_457 ),
	.shareout(Xd_0__inst_mult_1_458 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_137 (
// Equation(s):
// Xd_0__inst_mult_1_460  = SUM(( (!din_a[15] & (((din_a[14] & din_b[20])))) # (din_a[15] & (!din_b[19] $ (((!din_a[14]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_582  ) + ( Xd_0__inst_mult_1_581  ))
// Xd_0__inst_mult_1_461  = CARRY(( (!din_a[15] & (((din_a[14] & din_b[20])))) # (din_a[15] & (!din_b[19] $ (((!din_a[14]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_582  ) + ( Xd_0__inst_mult_1_581  ))
// Xd_0__inst_mult_1_462  = SHARE((din_a[15] & (din_b[19] & (din_a[14] & din_b[20]))))

	.dataa(!din_a[15]),
	.datab(!din_b[19]),
	.datac(!din_a[14]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_581 ),
	.sharein(Xd_0__inst_mult_1_582 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_460 ),
	.cout(Xd_0__inst_mult_1_461 ),
	.shareout(Xd_0__inst_mult_1_462 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_170 (
// Equation(s):
// Xd_0__inst_mult_6_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_582  = SHARE((din_a[76] & din_b[78]))

	.dataa(!din_a[76]),
	.datab(!din_b[78]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_581 ),
	.shareout(Xd_0__inst_mult_6_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_170 (
// Equation(s):
// Xd_0__inst_mult_7_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_582  = SHARE((din_a[88] & din_b[90]))

	.dataa(!din_a[88]),
	.datab(!din_b[90]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_581 ),
	.shareout(Xd_0__inst_mult_7_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_143 (
// Equation(s):
// Xd_0__inst_mult_4_472  = SUM(( (din_a[57] & din_b[50]) ) + ( Xd_0__inst_mult_4_454  ) + ( Xd_0__inst_mult_4_453  ))
// Xd_0__inst_mult_4_473  = CARRY(( (din_a[57] & din_b[50]) ) + ( Xd_0__inst_mult_4_454  ) + ( Xd_0__inst_mult_4_453  ))
// Xd_0__inst_mult_4_474  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[50]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_453 ),
	.sharein(Xd_0__inst_mult_4_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_472 ),
	.cout(Xd_0__inst_mult_4_473 ),
	.shareout(Xd_0__inst_mult_4_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_144 (
// Equation(s):
// Xd_0__inst_mult_4_476  = SUM(( (!din_a[56] & (((din_a[55] & din_b[52])))) # (din_a[56] & (!din_b[51] $ (((!din_a[55]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_458  ) + ( Xd_0__inst_mult_4_457  ))
// Xd_0__inst_mult_4_477  = CARRY(( (!din_a[56] & (((din_a[55] & din_b[52])))) # (din_a[56] & (!din_b[51] $ (((!din_a[55]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_458  ) + ( Xd_0__inst_mult_4_457  ))
// Xd_0__inst_mult_4_478  = SHARE((din_a[56] & (din_b[51] & (din_a[55] & din_b[52]))))

	.dataa(!din_a[56]),
	.datab(!din_b[51]),
	.datac(!din_a[55]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_457 ),
	.sharein(Xd_0__inst_mult_4_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_476 ),
	.cout(Xd_0__inst_mult_4_477 ),
	.shareout(Xd_0__inst_mult_4_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_145 (
// Equation(s):
// Xd_0__inst_mult_4_480  = SUM(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_4_462  ) + ( Xd_0__inst_mult_4_461  ))
// Xd_0__inst_mult_4_481  = CARRY(( (din_a[54] & din_b[53]) ) + ( Xd_0__inst_mult_4_462  ) + ( Xd_0__inst_mult_4_461  ))
// Xd_0__inst_mult_4_482  = SHARE((din_a[54] & din_b[54]))

	.dataa(!din_a[54]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_461 ),
	.sharein(Xd_0__inst_mult_4_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_480 ),
	.cout(Xd_0__inst_mult_4_481 ),
	.shareout(Xd_0__inst_mult_4_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_146 (
// Equation(s):
// Xd_0__inst_mult_4_484  = SUM(( (din_a[50] & din_b[57]) ) + ( Xd_0__inst_mult_4_466  ) + ( Xd_0__inst_mult_4_465  ))
// Xd_0__inst_mult_4_485  = CARRY(( (din_a[50] & din_b[57]) ) + ( Xd_0__inst_mult_4_466  ) + ( Xd_0__inst_mult_4_465  ))
// Xd_0__inst_mult_4_486  = SHARE((din_a[50] & din_b[58]))

	.dataa(!din_a[50]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_465 ),
	.sharein(Xd_0__inst_mult_4_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_484 ),
	.cout(Xd_0__inst_mult_4_485 ),
	.shareout(Xd_0__inst_mult_4_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_147 (
// Equation(s):
// Xd_0__inst_mult_4_488  = SUM(( (!din_a[52] & (((din_a[51] & din_b[56])))) # (din_a[52] & (!din_b[55] $ (((!din_a[51]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_470  ) + ( Xd_0__inst_mult_4_469  ))
// Xd_0__inst_mult_4_489  = CARRY(( (!din_a[52] & (((din_a[51] & din_b[56])))) # (din_a[52] & (!din_b[55] $ (((!din_a[51]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_470  ) + ( Xd_0__inst_mult_4_469  ))
// Xd_0__inst_mult_4_490  = SHARE((din_a[52] & (din_b[55] & (din_a[51] & din_b[56]))))

	.dataa(!din_a[52]),
	.datab(!din_b[55]),
	.datac(!din_a[51]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_469 ),
	.sharein(Xd_0__inst_mult_4_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_488 ),
	.cout(Xd_0__inst_mult_4_489 ),
	.shareout(Xd_0__inst_mult_4_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_142 (
// Equation(s):
// Xd_0__inst_mult_5_468  = SUM(( (din_a[69] & din_b[62]) ) + ( Xd_0__inst_mult_5_450  ) + ( Xd_0__inst_mult_5_449  ))
// Xd_0__inst_mult_5_469  = CARRY(( (din_a[69] & din_b[62]) ) + ( Xd_0__inst_mult_5_450  ) + ( Xd_0__inst_mult_5_449  ))
// Xd_0__inst_mult_5_470  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[62]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_449 ),
	.sharein(Xd_0__inst_mult_5_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_468 ),
	.cout(Xd_0__inst_mult_5_469 ),
	.shareout(Xd_0__inst_mult_5_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_143 (
// Equation(s):
// Xd_0__inst_mult_5_472  = SUM(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_454  ) + ( Xd_0__inst_mult_5_453  ))
// Xd_0__inst_mult_5_473  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[64])))) # (din_a[68] & (!din_b[63] $ (((!din_a[67]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_454  ) + ( Xd_0__inst_mult_5_453  ))
// Xd_0__inst_mult_5_474  = SHARE((din_a[68] & (din_b[63] & (din_a[67] & din_b[64]))))

	.dataa(!din_a[68]),
	.datab(!din_b[63]),
	.datac(!din_a[67]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_453 ),
	.sharein(Xd_0__inst_mult_5_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_472 ),
	.cout(Xd_0__inst_mult_5_473 ),
	.shareout(Xd_0__inst_mult_5_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_144 (
// Equation(s):
// Xd_0__inst_mult_5_476  = SUM(( (din_a[66] & din_b[65]) ) + ( Xd_0__inst_mult_5_458  ) + ( Xd_0__inst_mult_5_457  ))
// Xd_0__inst_mult_5_477  = CARRY(( (din_a[66] & din_b[65]) ) + ( Xd_0__inst_mult_5_458  ) + ( Xd_0__inst_mult_5_457  ))
// Xd_0__inst_mult_5_478  = SHARE((din_a[66] & din_b[66]))

	.dataa(!din_a[66]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_457 ),
	.sharein(Xd_0__inst_mult_5_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_476 ),
	.cout(Xd_0__inst_mult_5_477 ),
	.shareout(Xd_0__inst_mult_5_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_145 (
// Equation(s):
// Xd_0__inst_mult_5_480  = SUM(( (din_a[62] & din_b[69]) ) + ( Xd_0__inst_mult_5_462  ) + ( Xd_0__inst_mult_5_461  ))
// Xd_0__inst_mult_5_481  = CARRY(( (din_a[62] & din_b[69]) ) + ( Xd_0__inst_mult_5_462  ) + ( Xd_0__inst_mult_5_461  ))
// Xd_0__inst_mult_5_482  = SHARE((din_a[62] & din_b[70]))

	.dataa(!din_a[62]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_461 ),
	.sharein(Xd_0__inst_mult_5_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_480 ),
	.cout(Xd_0__inst_mult_5_481 ),
	.shareout(Xd_0__inst_mult_5_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_146 (
// Equation(s):
// Xd_0__inst_mult_5_484  = SUM(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_466  ) + ( Xd_0__inst_mult_5_465  ))
// Xd_0__inst_mult_5_485  = CARRY(( (!din_a[64] & (((din_a[63] & din_b[68])))) # (din_a[64] & (!din_b[67] $ (((!din_a[63]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_466  ) + ( Xd_0__inst_mult_5_465  ))
// Xd_0__inst_mult_5_486  = SHARE((din_a[64] & (din_b[67] & (din_a[63] & din_b[68]))))

	.dataa(!din_a[64]),
	.datab(!din_b[67]),
	.datac(!din_a[63]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_465 ),
	.sharein(Xd_0__inst_mult_5_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_484 ),
	.cout(Xd_0__inst_mult_5_485 ),
	.shareout(Xd_0__inst_mult_5_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_142 (
// Equation(s):
// Xd_0__inst_mult_2_468  = SUM(( (din_a[33] & din_b[26]) ) + ( Xd_0__inst_mult_2_450  ) + ( Xd_0__inst_mult_2_449  ))
// Xd_0__inst_mult_2_469  = CARRY(( (din_a[33] & din_b[26]) ) + ( Xd_0__inst_mult_2_450  ) + ( Xd_0__inst_mult_2_449  ))
// Xd_0__inst_mult_2_470  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[26]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_449 ),
	.sharein(Xd_0__inst_mult_2_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_468 ),
	.cout(Xd_0__inst_mult_2_469 ),
	.shareout(Xd_0__inst_mult_2_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_143 (
// Equation(s):
// Xd_0__inst_mult_2_472  = SUM(( (!din_a[32] & (((din_a[31] & din_b[28])))) # (din_a[32] & (!din_b[27] $ (((!din_a[31]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_454  ) + ( Xd_0__inst_mult_2_453  ))
// Xd_0__inst_mult_2_473  = CARRY(( (!din_a[32] & (((din_a[31] & din_b[28])))) # (din_a[32] & (!din_b[27] $ (((!din_a[31]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_454  ) + ( Xd_0__inst_mult_2_453  ))
// Xd_0__inst_mult_2_474  = SHARE((din_a[32] & (din_b[27] & (din_a[31] & din_b[28]))))

	.dataa(!din_a[32]),
	.datab(!din_b[27]),
	.datac(!din_a[31]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_453 ),
	.sharein(Xd_0__inst_mult_2_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_472 ),
	.cout(Xd_0__inst_mult_2_473 ),
	.shareout(Xd_0__inst_mult_2_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_144 (
// Equation(s):
// Xd_0__inst_mult_2_476  = SUM(( (din_a[30] & din_b[29]) ) + ( Xd_0__inst_mult_2_458  ) + ( Xd_0__inst_mult_2_457  ))
// Xd_0__inst_mult_2_477  = CARRY(( (din_a[30] & din_b[29]) ) + ( Xd_0__inst_mult_2_458  ) + ( Xd_0__inst_mult_2_457  ))
// Xd_0__inst_mult_2_478  = SHARE((din_a[30] & din_b[30]))

	.dataa(!din_a[30]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_457 ),
	.sharein(Xd_0__inst_mult_2_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_476 ),
	.cout(Xd_0__inst_mult_2_477 ),
	.shareout(Xd_0__inst_mult_2_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_145 (
// Equation(s):
// Xd_0__inst_mult_2_480  = SUM(( (din_a[26] & din_b[33]) ) + ( Xd_0__inst_mult_2_462  ) + ( Xd_0__inst_mult_2_461  ))
// Xd_0__inst_mult_2_481  = CARRY(( (din_a[26] & din_b[33]) ) + ( Xd_0__inst_mult_2_462  ) + ( Xd_0__inst_mult_2_461  ))
// Xd_0__inst_mult_2_482  = SHARE((din_a[26] & din_b[34]))

	.dataa(!din_a[26]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_461 ),
	.sharein(Xd_0__inst_mult_2_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_480 ),
	.cout(Xd_0__inst_mult_2_481 ),
	.shareout(Xd_0__inst_mult_2_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_146 (
// Equation(s):
// Xd_0__inst_mult_2_484  = SUM(( (!din_a[28] & (((din_a[27] & din_b[32])))) # (din_a[28] & (!din_b[31] $ (((!din_a[27]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_466  ) + ( Xd_0__inst_mult_2_465  ))
// Xd_0__inst_mult_2_485  = CARRY(( (!din_a[28] & (((din_a[27] & din_b[32])))) # (din_a[28] & (!din_b[31] $ (((!din_a[27]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_466  ) + ( Xd_0__inst_mult_2_465  ))
// Xd_0__inst_mult_2_486  = SHARE((din_a[28] & (din_b[31] & (din_a[27] & din_b[32]))))

	.dataa(!din_a[28]),
	.datab(!din_b[31]),
	.datac(!din_a[27]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_465 ),
	.sharein(Xd_0__inst_mult_2_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_484 ),
	.cout(Xd_0__inst_mult_2_485 ),
	.shareout(Xd_0__inst_mult_2_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_149 (
// Equation(s):
// Xd_0__inst_mult_3_508  = SUM(( (din_a[45] & din_b[38]) ) + ( Xd_0__inst_mult_3_490  ) + ( Xd_0__inst_mult_3_489  ))
// Xd_0__inst_mult_3_509  = CARRY(( (din_a[45] & din_b[38]) ) + ( Xd_0__inst_mult_3_490  ) + ( Xd_0__inst_mult_3_489  ))
// Xd_0__inst_mult_3_510  = SHARE(GND)

	.dataa(!din_a[45]),
	.datab(!din_b[38]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_489 ),
	.sharein(Xd_0__inst_mult_3_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_508 ),
	.cout(Xd_0__inst_mult_3_509 ),
	.shareout(Xd_0__inst_mult_3_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_150 (
// Equation(s):
// Xd_0__inst_mult_3_512  = SUM(( (!din_a[44] & (((din_a[43] & din_b[40])))) # (din_a[44] & (!din_b[39] $ (((!din_a[43]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_494  ) + ( Xd_0__inst_mult_3_493  ))
// Xd_0__inst_mult_3_513  = CARRY(( (!din_a[44] & (((din_a[43] & din_b[40])))) # (din_a[44] & (!din_b[39] $ (((!din_a[43]) # (!din_b[40]))))) ) + ( Xd_0__inst_mult_3_494  ) + ( Xd_0__inst_mult_3_493  ))
// Xd_0__inst_mult_3_514  = SHARE((din_a[44] & (din_b[39] & (din_a[43] & din_b[40]))))

	.dataa(!din_a[44]),
	.datab(!din_b[39]),
	.datac(!din_a[43]),
	.datad(!din_b[40]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_493 ),
	.sharein(Xd_0__inst_mult_3_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_512 ),
	.cout(Xd_0__inst_mult_3_513 ),
	.shareout(Xd_0__inst_mult_3_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_151 (
// Equation(s):
// Xd_0__inst_mult_3_516  = SUM(( (din_a[42] & din_b[41]) ) + ( Xd_0__inst_mult_3_498  ) + ( Xd_0__inst_mult_3_497  ))
// Xd_0__inst_mult_3_517  = CARRY(( (din_a[42] & din_b[41]) ) + ( Xd_0__inst_mult_3_498  ) + ( Xd_0__inst_mult_3_497  ))
// Xd_0__inst_mult_3_518  = SHARE((din_a[42] & din_b[42]))

	.dataa(!din_a[42]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_497 ),
	.sharein(Xd_0__inst_mult_3_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_516 ),
	.cout(Xd_0__inst_mult_3_517 ),
	.shareout(Xd_0__inst_mult_3_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_152 (
// Equation(s):
// Xd_0__inst_mult_3_520  = SUM(( (din_a[38] & din_b[45]) ) + ( Xd_0__inst_mult_3_502  ) + ( Xd_0__inst_mult_3_501  ))
// Xd_0__inst_mult_3_521  = CARRY(( (din_a[38] & din_b[45]) ) + ( Xd_0__inst_mult_3_502  ) + ( Xd_0__inst_mult_3_501  ))
// Xd_0__inst_mult_3_522  = SHARE((din_a[38] & din_b[46]))

	.dataa(!din_a[38]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_501 ),
	.sharein(Xd_0__inst_mult_3_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_520 ),
	.cout(Xd_0__inst_mult_3_521 ),
	.shareout(Xd_0__inst_mult_3_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_153 (
// Equation(s):
// Xd_0__inst_mult_3_524  = SUM(( (!din_a[40] & (((din_a[39] & din_b[44])))) # (din_a[40] & (!din_b[43] $ (((!din_a[39]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_506  ) + ( Xd_0__inst_mult_3_505  ))
// Xd_0__inst_mult_3_525  = CARRY(( (!din_a[40] & (((din_a[39] & din_b[44])))) # (din_a[40] & (!din_b[43] $ (((!din_a[39]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_506  ) + ( Xd_0__inst_mult_3_505  ))
// Xd_0__inst_mult_3_526  = SHARE((din_a[40] & (din_b[43] & (din_a[39] & din_b[44]))))

	.dataa(!din_a[40]),
	.datab(!din_b[43]),
	.datac(!din_a[39]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_505 ),
	.sharein(Xd_0__inst_mult_3_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_524 ),
	.cout(Xd_0__inst_mult_3_525 ),
	.shareout(Xd_0__inst_mult_3_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_142 (
// Equation(s):
// Xd_0__inst_mult_0_480  = SUM(( (din_a[9] & din_b[2]) ) + ( Xd_0__inst_mult_0_462  ) + ( Xd_0__inst_mult_0_461  ))
// Xd_0__inst_mult_0_481  = CARRY(( (din_a[9] & din_b[2]) ) + ( Xd_0__inst_mult_0_462  ) + ( Xd_0__inst_mult_0_461  ))
// Xd_0__inst_mult_0_482  = SHARE(GND)

	.dataa(!din_a[9]),
	.datab(!din_b[2]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_461 ),
	.sharein(Xd_0__inst_mult_0_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_480 ),
	.cout(Xd_0__inst_mult_0_481 ),
	.shareout(Xd_0__inst_mult_0_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_143 (
// Equation(s):
// Xd_0__inst_mult_0_484  = SUM(( (!din_a[8] & (((din_a[7] & din_b[4])))) # (din_a[8] & (!din_b[3] $ (((!din_a[7]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_466  ) + ( Xd_0__inst_mult_0_465  ))
// Xd_0__inst_mult_0_485  = CARRY(( (!din_a[8] & (((din_a[7] & din_b[4])))) # (din_a[8] & (!din_b[3] $ (((!din_a[7]) # (!din_b[4]))))) ) + ( Xd_0__inst_mult_0_466  ) + ( Xd_0__inst_mult_0_465  ))
// Xd_0__inst_mult_0_486  = SHARE((din_a[8] & (din_b[3] & (din_a[7] & din_b[4]))))

	.dataa(!din_a[8]),
	.datab(!din_b[3]),
	.datac(!din_a[7]),
	.datad(!din_b[4]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_465 ),
	.sharein(Xd_0__inst_mult_0_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_484 ),
	.cout(Xd_0__inst_mult_0_485 ),
	.shareout(Xd_0__inst_mult_0_486 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_144 (
// Equation(s):
// Xd_0__inst_mult_0_488  = SUM(( (din_a[6] & din_b[5]) ) + ( Xd_0__inst_mult_0_470  ) + ( Xd_0__inst_mult_0_469  ))
// Xd_0__inst_mult_0_489  = CARRY(( (din_a[6] & din_b[5]) ) + ( Xd_0__inst_mult_0_470  ) + ( Xd_0__inst_mult_0_469  ))
// Xd_0__inst_mult_0_490  = SHARE((din_a[6] & din_b[6]))

	.dataa(!din_a[6]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_469 ),
	.sharein(Xd_0__inst_mult_0_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_488 ),
	.cout(Xd_0__inst_mult_0_489 ),
	.shareout(Xd_0__inst_mult_0_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_145 (
// Equation(s):
// Xd_0__inst_mult_0_492  = SUM(( (din_a[2] & din_b[9]) ) + ( Xd_0__inst_mult_0_474  ) + ( Xd_0__inst_mult_0_473  ))
// Xd_0__inst_mult_0_493  = CARRY(( (din_a[2] & din_b[9]) ) + ( Xd_0__inst_mult_0_474  ) + ( Xd_0__inst_mult_0_473  ))
// Xd_0__inst_mult_0_494  = SHARE((din_a[2] & din_b[10]))

	.dataa(!din_a[2]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_473 ),
	.sharein(Xd_0__inst_mult_0_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_492 ),
	.cout(Xd_0__inst_mult_0_493 ),
	.shareout(Xd_0__inst_mult_0_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_146 (
// Equation(s):
// Xd_0__inst_mult_0_496  = SUM(( (!din_a[4] & (((din_a[3] & din_b[8])))) # (din_a[4] & (!din_b[7] $ (((!din_a[3]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_478  ) + ( Xd_0__inst_mult_0_477  ))
// Xd_0__inst_mult_0_497  = CARRY(( (!din_a[4] & (((din_a[3] & din_b[8])))) # (din_a[4] & (!din_b[7] $ (((!din_a[3]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_478  ) + ( Xd_0__inst_mult_0_477  ))
// Xd_0__inst_mult_0_498  = SHARE((din_a[4] & (din_b[7] & (din_a[3] & din_b[8]))))

	.dataa(!din_a[4]),
	.datab(!din_b[7]),
	.datac(!din_a[3]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_477 ),
	.sharein(Xd_0__inst_mult_0_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_496 ),
	.cout(Xd_0__inst_mult_0_497 ),
	.shareout(Xd_0__inst_mult_0_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_138 (
// Equation(s):
// Xd_0__inst_mult_1_464  = SUM(( (din_a[21] & din_b[14]) ) + ( Xd_0__inst_mult_1_446  ) + ( Xd_0__inst_mult_1_445  ))
// Xd_0__inst_mult_1_465  = CARRY(( (din_a[21] & din_b[14]) ) + ( Xd_0__inst_mult_1_446  ) + ( Xd_0__inst_mult_1_445  ))
// Xd_0__inst_mult_1_466  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[14]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_445 ),
	.sharein(Xd_0__inst_mult_1_446 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_464 ),
	.cout(Xd_0__inst_mult_1_465 ),
	.shareout(Xd_0__inst_mult_1_466 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_139 (
// Equation(s):
// Xd_0__inst_mult_1_468  = SUM(( (!din_a[20] & (((din_a[19] & din_b[16])))) # (din_a[20] & (!din_b[15] $ (((!din_a[19]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_450  ) + ( Xd_0__inst_mult_1_449  ))
// Xd_0__inst_mult_1_469  = CARRY(( (!din_a[20] & (((din_a[19] & din_b[16])))) # (din_a[20] & (!din_b[15] $ (((!din_a[19]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_450  ) + ( Xd_0__inst_mult_1_449  ))
// Xd_0__inst_mult_1_470  = SHARE((din_a[20] & (din_b[15] & (din_a[19] & din_b[16]))))

	.dataa(!din_a[20]),
	.datab(!din_b[15]),
	.datac(!din_a[19]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_449 ),
	.sharein(Xd_0__inst_mult_1_450 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_468 ),
	.cout(Xd_0__inst_mult_1_469 ),
	.shareout(Xd_0__inst_mult_1_470 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_140 (
// Equation(s):
// Xd_0__inst_mult_1_472  = SUM(( (din_a[18] & din_b[17]) ) + ( Xd_0__inst_mult_1_454  ) + ( Xd_0__inst_mult_1_453  ))
// Xd_0__inst_mult_1_473  = CARRY(( (din_a[18] & din_b[17]) ) + ( Xd_0__inst_mult_1_454  ) + ( Xd_0__inst_mult_1_453  ))
// Xd_0__inst_mult_1_474  = SHARE((din_a[18] & din_b[18]))

	.dataa(!din_a[18]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_453 ),
	.sharein(Xd_0__inst_mult_1_454 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_472 ),
	.cout(Xd_0__inst_mult_1_473 ),
	.shareout(Xd_0__inst_mult_1_474 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_141 (
// Equation(s):
// Xd_0__inst_mult_1_476  = SUM(( (din_a[14] & din_b[21]) ) + ( Xd_0__inst_mult_1_458  ) + ( Xd_0__inst_mult_1_457  ))
// Xd_0__inst_mult_1_477  = CARRY(( (din_a[14] & din_b[21]) ) + ( Xd_0__inst_mult_1_458  ) + ( Xd_0__inst_mult_1_457  ))
// Xd_0__inst_mult_1_478  = SHARE((din_a[14] & din_b[22]))

	.dataa(!din_a[14]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_457 ),
	.sharein(Xd_0__inst_mult_1_458 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_476 ),
	.cout(Xd_0__inst_mult_1_477 ),
	.shareout(Xd_0__inst_mult_1_478 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_142 (
// Equation(s):
// Xd_0__inst_mult_1_480  = SUM(( (!din_a[16] & (((din_a[15] & din_b[20])))) # (din_a[16] & (!din_b[19] $ (((!din_a[15]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_462  ) + ( Xd_0__inst_mult_1_461  ))
// Xd_0__inst_mult_1_481  = CARRY(( (!din_a[16] & (((din_a[15] & din_b[20])))) # (din_a[16] & (!din_b[19] $ (((!din_a[15]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_462  ) + ( Xd_0__inst_mult_1_461  ))
// Xd_0__inst_mult_1_482  = SHARE((din_a[16] & (din_b[19] & (din_a[15] & din_b[20]))))

	.dataa(!din_a[16]),
	.datab(!din_b[19]),
	.datac(!din_a[15]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_461 ),
	.sharein(Xd_0__inst_mult_1_462 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_480 ),
	.cout(Xd_0__inst_mult_1_481 ),
	.shareout(Xd_0__inst_mult_1_482 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_148 (
// Equation(s):
// Xd_0__inst_mult_4_492  = SUM(( GND ) + ( Xd_0__inst_mult_4_474  ) + ( Xd_0__inst_mult_4_473  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_473 ),
	.sharein(Xd_0__inst_mult_4_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_492 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_149 (
// Equation(s):
// Xd_0__inst_mult_4_496  = SUM(( (!din_a[57] & (((din_a[56] & din_b[52])))) # (din_a[57] & (!din_b[51] $ (((!din_a[56]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_478  ) + ( Xd_0__inst_mult_4_477  ))
// Xd_0__inst_mult_4_497  = CARRY(( (!din_a[57] & (((din_a[56] & din_b[52])))) # (din_a[57] & (!din_b[51] $ (((!din_a[56]) # (!din_b[52]))))) ) + ( Xd_0__inst_mult_4_478  ) + ( Xd_0__inst_mult_4_477  ))
// Xd_0__inst_mult_4_498  = SHARE((din_a[57] & (din_b[51] & (din_a[56] & din_b[52]))))

	.dataa(!din_a[57]),
	.datab(!din_b[51]),
	.datac(!din_a[56]),
	.datad(!din_b[52]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_477 ),
	.sharein(Xd_0__inst_mult_4_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_496 ),
	.cout(Xd_0__inst_mult_4_497 ),
	.shareout(Xd_0__inst_mult_4_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_150 (
// Equation(s):
// Xd_0__inst_mult_4_500  = SUM(( (din_a[55] & din_b[53]) ) + ( Xd_0__inst_mult_4_482  ) + ( Xd_0__inst_mult_4_481  ))
// Xd_0__inst_mult_4_501  = CARRY(( (din_a[55] & din_b[53]) ) + ( Xd_0__inst_mult_4_482  ) + ( Xd_0__inst_mult_4_481  ))
// Xd_0__inst_mult_4_502  = SHARE((din_a[55] & din_b[54]))

	.dataa(!din_a[55]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_481 ),
	.sharein(Xd_0__inst_mult_4_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_500 ),
	.cout(Xd_0__inst_mult_4_501 ),
	.shareout(Xd_0__inst_mult_4_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_151 (
// Equation(s):
// Xd_0__inst_mult_4_504  = SUM(( (din_a[51] & din_b[57]) ) + ( Xd_0__inst_mult_4_486  ) + ( Xd_0__inst_mult_4_485  ))
// Xd_0__inst_mult_4_505  = CARRY(( (din_a[51] & din_b[57]) ) + ( Xd_0__inst_mult_4_486  ) + ( Xd_0__inst_mult_4_485  ))
// Xd_0__inst_mult_4_506  = SHARE((din_a[51] & din_b[58]))

	.dataa(!din_a[51]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_485 ),
	.sharein(Xd_0__inst_mult_4_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_504 ),
	.cout(Xd_0__inst_mult_4_505 ),
	.shareout(Xd_0__inst_mult_4_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_152 (
// Equation(s):
// Xd_0__inst_mult_4_508  = SUM(( (!din_a[53] & (((din_a[52] & din_b[56])))) # (din_a[53] & (!din_b[55] $ (((!din_a[52]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_490  ) + ( Xd_0__inst_mult_4_489  ))
// Xd_0__inst_mult_4_509  = CARRY(( (!din_a[53] & (((din_a[52] & din_b[56])))) # (din_a[53] & (!din_b[55] $ (((!din_a[52]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_490  ) + ( Xd_0__inst_mult_4_489  ))
// Xd_0__inst_mult_4_510  = SHARE((din_a[53] & (din_b[55] & (din_a[52] & din_b[56]))))

	.dataa(!din_a[53]),
	.datab(!din_b[55]),
	.datac(!din_a[52]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_489 ),
	.sharein(Xd_0__inst_mult_4_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_508 ),
	.cout(Xd_0__inst_mult_4_509 ),
	.shareout(Xd_0__inst_mult_4_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_147 (
// Equation(s):
// Xd_0__inst_mult_5_488  = SUM(( GND ) + ( Xd_0__inst_mult_5_470  ) + ( Xd_0__inst_mult_5_469  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_469 ),
	.sharein(Xd_0__inst_mult_5_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_488 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_148 (
// Equation(s):
// Xd_0__inst_mult_5_492  = SUM(( (!din_a[69] & (((din_a[68] & din_b[64])))) # (din_a[69] & (!din_b[63] $ (((!din_a[68]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_474  ) + ( Xd_0__inst_mult_5_473  ))
// Xd_0__inst_mult_5_493  = CARRY(( (!din_a[69] & (((din_a[68] & din_b[64])))) # (din_a[69] & (!din_b[63] $ (((!din_a[68]) # (!din_b[64]))))) ) + ( Xd_0__inst_mult_5_474  ) + ( Xd_0__inst_mult_5_473  ))
// Xd_0__inst_mult_5_494  = SHARE((din_a[69] & (din_b[63] & (din_a[68] & din_b[64]))))

	.dataa(!din_a[69]),
	.datab(!din_b[63]),
	.datac(!din_a[68]),
	.datad(!din_b[64]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_473 ),
	.sharein(Xd_0__inst_mult_5_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_492 ),
	.cout(Xd_0__inst_mult_5_493 ),
	.shareout(Xd_0__inst_mult_5_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_149 (
// Equation(s):
// Xd_0__inst_mult_5_496  = SUM(( (din_a[67] & din_b[65]) ) + ( Xd_0__inst_mult_5_478  ) + ( Xd_0__inst_mult_5_477  ))
// Xd_0__inst_mult_5_497  = CARRY(( (din_a[67] & din_b[65]) ) + ( Xd_0__inst_mult_5_478  ) + ( Xd_0__inst_mult_5_477  ))
// Xd_0__inst_mult_5_498  = SHARE((din_a[67] & din_b[66]))

	.dataa(!din_a[67]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_477 ),
	.sharein(Xd_0__inst_mult_5_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_496 ),
	.cout(Xd_0__inst_mult_5_497 ),
	.shareout(Xd_0__inst_mult_5_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_150 (
// Equation(s):
// Xd_0__inst_mult_5_500  = SUM(( (din_a[63] & din_b[69]) ) + ( Xd_0__inst_mult_5_482  ) + ( Xd_0__inst_mult_5_481  ))
// Xd_0__inst_mult_5_501  = CARRY(( (din_a[63] & din_b[69]) ) + ( Xd_0__inst_mult_5_482  ) + ( Xd_0__inst_mult_5_481  ))
// Xd_0__inst_mult_5_502  = SHARE((din_a[63] & din_b[70]))

	.dataa(!din_a[63]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_481 ),
	.sharein(Xd_0__inst_mult_5_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_500 ),
	.cout(Xd_0__inst_mult_5_501 ),
	.shareout(Xd_0__inst_mult_5_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_151 (
// Equation(s):
// Xd_0__inst_mult_5_504  = SUM(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_486  ) + ( Xd_0__inst_mult_5_485  ))
// Xd_0__inst_mult_5_505  = CARRY(( (!din_a[65] & (((din_a[64] & din_b[68])))) # (din_a[65] & (!din_b[67] $ (((!din_a[64]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_486  ) + ( Xd_0__inst_mult_5_485  ))
// Xd_0__inst_mult_5_506  = SHARE((din_a[65] & (din_b[67] & (din_a[64] & din_b[68]))))

	.dataa(!din_a[65]),
	.datab(!din_b[67]),
	.datac(!din_a[64]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_485 ),
	.sharein(Xd_0__inst_mult_5_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_504 ),
	.cout(Xd_0__inst_mult_5_505 ),
	.shareout(Xd_0__inst_mult_5_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_147 (
// Equation(s):
// Xd_0__inst_mult_2_488  = SUM(( GND ) + ( Xd_0__inst_mult_2_470  ) + ( Xd_0__inst_mult_2_469  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_469 ),
	.sharein(Xd_0__inst_mult_2_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_488 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_148 (
// Equation(s):
// Xd_0__inst_mult_2_492  = SUM(( (!din_a[33] & (((din_a[32] & din_b[28])))) # (din_a[33] & (!din_b[27] $ (((!din_a[32]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_474  ) + ( Xd_0__inst_mult_2_473  ))
// Xd_0__inst_mult_2_493  = CARRY(( (!din_a[33] & (((din_a[32] & din_b[28])))) # (din_a[33] & (!din_b[27] $ (((!din_a[32]) # (!din_b[28]))))) ) + ( Xd_0__inst_mult_2_474  ) + ( Xd_0__inst_mult_2_473  ))
// Xd_0__inst_mult_2_494  = SHARE((din_a[33] & (din_b[27] & (din_a[32] & din_b[28]))))

	.dataa(!din_a[33]),
	.datab(!din_b[27]),
	.datac(!din_a[32]),
	.datad(!din_b[28]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_473 ),
	.sharein(Xd_0__inst_mult_2_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_492 ),
	.cout(Xd_0__inst_mult_2_493 ),
	.shareout(Xd_0__inst_mult_2_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_149 (
// Equation(s):
// Xd_0__inst_mult_2_496  = SUM(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_2_478  ) + ( Xd_0__inst_mult_2_477  ))
// Xd_0__inst_mult_2_497  = CARRY(( (din_a[31] & din_b[29]) ) + ( Xd_0__inst_mult_2_478  ) + ( Xd_0__inst_mult_2_477  ))
// Xd_0__inst_mult_2_498  = SHARE((din_a[31] & din_b[30]))

	.dataa(!din_a[31]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_477 ),
	.sharein(Xd_0__inst_mult_2_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_496 ),
	.cout(Xd_0__inst_mult_2_497 ),
	.shareout(Xd_0__inst_mult_2_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_150 (
// Equation(s):
// Xd_0__inst_mult_2_500  = SUM(( (din_a[27] & din_b[33]) ) + ( Xd_0__inst_mult_2_482  ) + ( Xd_0__inst_mult_2_481  ))
// Xd_0__inst_mult_2_501  = CARRY(( (din_a[27] & din_b[33]) ) + ( Xd_0__inst_mult_2_482  ) + ( Xd_0__inst_mult_2_481  ))
// Xd_0__inst_mult_2_502  = SHARE((din_a[27] & din_b[34]))

	.dataa(!din_a[27]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_481 ),
	.sharein(Xd_0__inst_mult_2_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_500 ),
	.cout(Xd_0__inst_mult_2_501 ),
	.shareout(Xd_0__inst_mult_2_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_151 (
// Equation(s):
// Xd_0__inst_mult_2_504  = SUM(( (!din_a[29] & (((din_a[28] & din_b[32])))) # (din_a[29] & (!din_b[31] $ (((!din_a[28]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_486  ) + ( Xd_0__inst_mult_2_485  ))
// Xd_0__inst_mult_2_505  = CARRY(( (!din_a[29] & (((din_a[28] & din_b[32])))) # (din_a[29] & (!din_b[31] $ (((!din_a[28]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_486  ) + ( Xd_0__inst_mult_2_485  ))
// Xd_0__inst_mult_2_506  = SHARE((din_a[29] & (din_b[31] & (din_a[28] & din_b[32]))))

	.dataa(!din_a[29]),
	.datab(!din_b[31]),
	.datac(!din_a[28]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_485 ),
	.sharein(Xd_0__inst_mult_2_486 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_504 ),
	.cout(Xd_0__inst_mult_2_505 ),
	.shareout(Xd_0__inst_mult_2_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_154 (
// Equation(s):
// Xd_0__inst_mult_3_528  = SUM(( (din_a[43] & din_b[41]) ) + ( Xd_0__inst_mult_3_518  ) + ( Xd_0__inst_mult_3_517  ))
// Xd_0__inst_mult_3_529  = CARRY(( (din_a[43] & din_b[41]) ) + ( Xd_0__inst_mult_3_518  ) + ( Xd_0__inst_mult_3_517  ))
// Xd_0__inst_mult_3_530  = SHARE((din_a[43] & din_b[42]))

	.dataa(!din_a[43]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_517 ),
	.sharein(Xd_0__inst_mult_3_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_528 ),
	.cout(Xd_0__inst_mult_3_529 ),
	.shareout(Xd_0__inst_mult_3_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_155 (
// Equation(s):
// Xd_0__inst_mult_3_532  = SUM(( (din_a[39] & din_b[45]) ) + ( Xd_0__inst_mult_3_522  ) + ( Xd_0__inst_mult_3_521  ))
// Xd_0__inst_mult_3_533  = CARRY(( (din_a[39] & din_b[45]) ) + ( Xd_0__inst_mult_3_522  ) + ( Xd_0__inst_mult_3_521  ))
// Xd_0__inst_mult_3_534  = SHARE((din_a[39] & din_b[46]))

	.dataa(!din_a[39]),
	.datab(!din_b[45]),
	.datac(!din_b[46]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_521 ),
	.sharein(Xd_0__inst_mult_3_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_532 ),
	.cout(Xd_0__inst_mult_3_533 ),
	.shareout(Xd_0__inst_mult_3_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_156 (
// Equation(s):
// Xd_0__inst_mult_3_536  = SUM(( (!din_a[41] & (((din_a[40] & din_b[44])))) # (din_a[41] & (!din_b[43] $ (((!din_a[40]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_526  ) + ( Xd_0__inst_mult_3_525  ))
// Xd_0__inst_mult_3_537  = CARRY(( (!din_a[41] & (((din_a[40] & din_b[44])))) # (din_a[41] & (!din_b[43] $ (((!din_a[40]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_526  ) + ( Xd_0__inst_mult_3_525  ))
// Xd_0__inst_mult_3_538  = SHARE((din_a[41] & (din_b[43] & (din_a[40] & din_b[44]))))

	.dataa(!din_a[41]),
	.datab(!din_b[43]),
	.datac(!din_a[40]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_525 ),
	.sharein(Xd_0__inst_mult_3_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_536 ),
	.cout(Xd_0__inst_mult_3_537 ),
	.shareout(Xd_0__inst_mult_3_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_147 (
// Equation(s):
// Xd_0__inst_mult_0_500  = SUM(( (din_a[7] & din_b[5]) ) + ( Xd_0__inst_mult_0_490  ) + ( Xd_0__inst_mult_0_489  ))
// Xd_0__inst_mult_0_501  = CARRY(( (din_a[7] & din_b[5]) ) + ( Xd_0__inst_mult_0_490  ) + ( Xd_0__inst_mult_0_489  ))
// Xd_0__inst_mult_0_502  = SHARE((din_a[7] & din_b[6]))

	.dataa(!din_a[7]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_489 ),
	.sharein(Xd_0__inst_mult_0_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_500 ),
	.cout(Xd_0__inst_mult_0_501 ),
	.shareout(Xd_0__inst_mult_0_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_148 (
// Equation(s):
// Xd_0__inst_mult_0_504  = SUM(( (din_a[3] & din_b[9]) ) + ( Xd_0__inst_mult_0_494  ) + ( Xd_0__inst_mult_0_493  ))
// Xd_0__inst_mult_0_505  = CARRY(( (din_a[3] & din_b[9]) ) + ( Xd_0__inst_mult_0_494  ) + ( Xd_0__inst_mult_0_493  ))
// Xd_0__inst_mult_0_506  = SHARE((din_a[3] & din_b[10]))

	.dataa(!din_a[3]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_493 ),
	.sharein(Xd_0__inst_mult_0_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_504 ),
	.cout(Xd_0__inst_mult_0_505 ),
	.shareout(Xd_0__inst_mult_0_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_149 (
// Equation(s):
// Xd_0__inst_mult_0_508  = SUM(( (!din_a[5] & (((din_a[4] & din_b[8])))) # (din_a[5] & (!din_b[7] $ (((!din_a[4]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_498  ) + ( Xd_0__inst_mult_0_497  ))
// Xd_0__inst_mult_0_509  = CARRY(( (!din_a[5] & (((din_a[4] & din_b[8])))) # (din_a[5] & (!din_b[7] $ (((!din_a[4]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_498  ) + ( Xd_0__inst_mult_0_497  ))
// Xd_0__inst_mult_0_510  = SHARE((din_a[5] & (din_b[7] & (din_a[4] & din_b[8]))))

	.dataa(!din_a[5]),
	.datab(!din_b[7]),
	.datac(!din_a[4]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_497 ),
	.sharein(Xd_0__inst_mult_0_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_508 ),
	.cout(Xd_0__inst_mult_0_509 ),
	.shareout(Xd_0__inst_mult_0_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_143 (
// Equation(s):
// Xd_0__inst_mult_1_484  = SUM(( GND ) + ( Xd_0__inst_mult_1_466  ) + ( Xd_0__inst_mult_1_465  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_465 ),
	.sharein(Xd_0__inst_mult_1_466 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_484 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_144 (
// Equation(s):
// Xd_0__inst_mult_1_488  = SUM(( (!din_a[21] & (((din_a[20] & din_b[16])))) # (din_a[21] & (!din_b[15] $ (((!din_a[20]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_470  ) + ( Xd_0__inst_mult_1_469  ))
// Xd_0__inst_mult_1_489  = CARRY(( (!din_a[21] & (((din_a[20] & din_b[16])))) # (din_a[21] & (!din_b[15] $ (((!din_a[20]) # (!din_b[16]))))) ) + ( Xd_0__inst_mult_1_470  ) + ( Xd_0__inst_mult_1_469  ))
// Xd_0__inst_mult_1_490  = SHARE((din_a[21] & (din_b[15] & (din_a[20] & din_b[16]))))

	.dataa(!din_a[21]),
	.datab(!din_b[15]),
	.datac(!din_a[20]),
	.datad(!din_b[16]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_469 ),
	.sharein(Xd_0__inst_mult_1_470 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_488 ),
	.cout(Xd_0__inst_mult_1_489 ),
	.shareout(Xd_0__inst_mult_1_490 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_145 (
// Equation(s):
// Xd_0__inst_mult_1_492  = SUM(( (din_a[19] & din_b[17]) ) + ( Xd_0__inst_mult_1_474  ) + ( Xd_0__inst_mult_1_473  ))
// Xd_0__inst_mult_1_493  = CARRY(( (din_a[19] & din_b[17]) ) + ( Xd_0__inst_mult_1_474  ) + ( Xd_0__inst_mult_1_473  ))
// Xd_0__inst_mult_1_494  = SHARE((din_a[19] & din_b[18]))

	.dataa(!din_a[19]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_473 ),
	.sharein(Xd_0__inst_mult_1_474 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_492 ),
	.cout(Xd_0__inst_mult_1_493 ),
	.shareout(Xd_0__inst_mult_1_494 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_146 (
// Equation(s):
// Xd_0__inst_mult_1_496  = SUM(( (din_a[15] & din_b[21]) ) + ( Xd_0__inst_mult_1_478  ) + ( Xd_0__inst_mult_1_477  ))
// Xd_0__inst_mult_1_497  = CARRY(( (din_a[15] & din_b[21]) ) + ( Xd_0__inst_mult_1_478  ) + ( Xd_0__inst_mult_1_477  ))
// Xd_0__inst_mult_1_498  = SHARE((din_a[15] & din_b[22]))

	.dataa(!din_a[15]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_477 ),
	.sharein(Xd_0__inst_mult_1_478 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_496 ),
	.cout(Xd_0__inst_mult_1_497 ),
	.shareout(Xd_0__inst_mult_1_498 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_147 (
// Equation(s):
// Xd_0__inst_mult_1_500  = SUM(( (!din_a[17] & (((din_a[16] & din_b[20])))) # (din_a[17] & (!din_b[19] $ (((!din_a[16]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_482  ) + ( Xd_0__inst_mult_1_481  ))
// Xd_0__inst_mult_1_501  = CARRY(( (!din_a[17] & (((din_a[16] & din_b[20])))) # (din_a[17] & (!din_b[19] $ (((!din_a[16]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_482  ) + ( Xd_0__inst_mult_1_481  ))
// Xd_0__inst_mult_1_502  = SHARE((din_a[17] & (din_b[19] & (din_a[16] & din_b[20]))))

	.dataa(!din_a[17]),
	.datab(!din_b[19]),
	.datac(!din_a[16]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_481 ),
	.sharein(Xd_0__inst_mult_1_482 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_500 ),
	.cout(Xd_0__inst_mult_1_501 ),
	.shareout(Xd_0__inst_mult_1_502 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_153 (
// Equation(s):
// Xd_0__inst_mult_4_512  = SUM(( (din_a[57] & din_b[52]) ) + ( Xd_0__inst_mult_4_498  ) + ( Xd_0__inst_mult_4_497  ))
// Xd_0__inst_mult_4_513  = CARRY(( (din_a[57] & din_b[52]) ) + ( Xd_0__inst_mult_4_498  ) + ( Xd_0__inst_mult_4_497  ))
// Xd_0__inst_mult_4_514  = SHARE(GND)

	.dataa(!din_a[57]),
	.datab(!din_b[52]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_497 ),
	.sharein(Xd_0__inst_mult_4_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_512 ),
	.cout(Xd_0__inst_mult_4_513 ),
	.shareout(Xd_0__inst_mult_4_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_154 (
// Equation(s):
// Xd_0__inst_mult_4_516  = SUM(( (din_a[56] & din_b[53]) ) + ( Xd_0__inst_mult_4_502  ) + ( Xd_0__inst_mult_4_501  ))
// Xd_0__inst_mult_4_517  = CARRY(( (din_a[56] & din_b[53]) ) + ( Xd_0__inst_mult_4_502  ) + ( Xd_0__inst_mult_4_501  ))
// Xd_0__inst_mult_4_518  = SHARE((din_a[56] & din_b[54]))

	.dataa(!din_a[56]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_501 ),
	.sharein(Xd_0__inst_mult_4_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_516 ),
	.cout(Xd_0__inst_mult_4_517 ),
	.shareout(Xd_0__inst_mult_4_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_155 (
// Equation(s):
// Xd_0__inst_mult_4_520  = SUM(( (din_a[52] & din_b[57]) ) + ( Xd_0__inst_mult_4_506  ) + ( Xd_0__inst_mult_4_505  ))
// Xd_0__inst_mult_4_521  = CARRY(( (din_a[52] & din_b[57]) ) + ( Xd_0__inst_mult_4_506  ) + ( Xd_0__inst_mult_4_505  ))
// Xd_0__inst_mult_4_522  = SHARE((din_a[52] & din_b[58]))

	.dataa(!din_a[52]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_505 ),
	.sharein(Xd_0__inst_mult_4_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_520 ),
	.cout(Xd_0__inst_mult_4_521 ),
	.shareout(Xd_0__inst_mult_4_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_156 (
// Equation(s):
// Xd_0__inst_mult_4_524  = SUM(( (!din_a[54] & (((din_a[53] & din_b[56])))) # (din_a[54] & (!din_b[55] $ (((!din_a[53]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_510  ) + ( Xd_0__inst_mult_4_509  ))
// Xd_0__inst_mult_4_525  = CARRY(( (!din_a[54] & (((din_a[53] & din_b[56])))) # (din_a[54] & (!din_b[55] $ (((!din_a[53]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_510  ) + ( Xd_0__inst_mult_4_509  ))
// Xd_0__inst_mult_4_526  = SHARE((din_a[54] & (din_b[55] & (din_a[53] & din_b[56]))))

	.dataa(!din_a[54]),
	.datab(!din_b[55]),
	.datac(!din_a[53]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_509 ),
	.sharein(Xd_0__inst_mult_4_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_524 ),
	.cout(Xd_0__inst_mult_4_525 ),
	.shareout(Xd_0__inst_mult_4_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_152 (
// Equation(s):
// Xd_0__inst_mult_5_508  = SUM(( (din_a[69] & din_b[64]) ) + ( Xd_0__inst_mult_5_494  ) + ( Xd_0__inst_mult_5_493  ))
// Xd_0__inst_mult_5_509  = CARRY(( (din_a[69] & din_b[64]) ) + ( Xd_0__inst_mult_5_494  ) + ( Xd_0__inst_mult_5_493  ))
// Xd_0__inst_mult_5_510  = SHARE(GND)

	.dataa(!din_a[69]),
	.datab(!din_b[64]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_493 ),
	.sharein(Xd_0__inst_mult_5_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_508 ),
	.cout(Xd_0__inst_mult_5_509 ),
	.shareout(Xd_0__inst_mult_5_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_153 (
// Equation(s):
// Xd_0__inst_mult_5_512  = SUM(( (din_a[68] & din_b[65]) ) + ( Xd_0__inst_mult_5_498  ) + ( Xd_0__inst_mult_5_497  ))
// Xd_0__inst_mult_5_513  = CARRY(( (din_a[68] & din_b[65]) ) + ( Xd_0__inst_mult_5_498  ) + ( Xd_0__inst_mult_5_497  ))
// Xd_0__inst_mult_5_514  = SHARE((din_a[68] & din_b[66]))

	.dataa(!din_a[68]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_497 ),
	.sharein(Xd_0__inst_mult_5_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_512 ),
	.cout(Xd_0__inst_mult_5_513 ),
	.shareout(Xd_0__inst_mult_5_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_154 (
// Equation(s):
// Xd_0__inst_mult_5_516  = SUM(( (din_a[64] & din_b[69]) ) + ( Xd_0__inst_mult_5_502  ) + ( Xd_0__inst_mult_5_501  ))
// Xd_0__inst_mult_5_517  = CARRY(( (din_a[64] & din_b[69]) ) + ( Xd_0__inst_mult_5_502  ) + ( Xd_0__inst_mult_5_501  ))
// Xd_0__inst_mult_5_518  = SHARE((din_a[64] & din_b[70]))

	.dataa(!din_a[64]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_501 ),
	.sharein(Xd_0__inst_mult_5_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_516 ),
	.cout(Xd_0__inst_mult_5_517 ),
	.shareout(Xd_0__inst_mult_5_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_155 (
// Equation(s):
// Xd_0__inst_mult_5_520  = SUM(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_506  ) + ( Xd_0__inst_mult_5_505  ))
// Xd_0__inst_mult_5_521  = CARRY(( (!din_a[66] & (((din_a[65] & din_b[68])))) # (din_a[66] & (!din_b[67] $ (((!din_a[65]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_506  ) + ( Xd_0__inst_mult_5_505  ))
// Xd_0__inst_mult_5_522  = SHARE((din_a[66] & (din_b[67] & (din_a[65] & din_b[68]))))

	.dataa(!din_a[66]),
	.datab(!din_b[67]),
	.datac(!din_a[65]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_505 ),
	.sharein(Xd_0__inst_mult_5_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_520 ),
	.cout(Xd_0__inst_mult_5_521 ),
	.shareout(Xd_0__inst_mult_5_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_152 (
// Equation(s):
// Xd_0__inst_mult_2_508  = SUM(( (din_a[33] & din_b[28]) ) + ( Xd_0__inst_mult_2_494  ) + ( Xd_0__inst_mult_2_493  ))
// Xd_0__inst_mult_2_509  = CARRY(( (din_a[33] & din_b[28]) ) + ( Xd_0__inst_mult_2_494  ) + ( Xd_0__inst_mult_2_493  ))
// Xd_0__inst_mult_2_510  = SHARE(GND)

	.dataa(!din_a[33]),
	.datab(!din_b[28]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_493 ),
	.sharein(Xd_0__inst_mult_2_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_508 ),
	.cout(Xd_0__inst_mult_2_509 ),
	.shareout(Xd_0__inst_mult_2_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_153 (
// Equation(s):
// Xd_0__inst_mult_2_512  = SUM(( (din_a[32] & din_b[29]) ) + ( Xd_0__inst_mult_2_498  ) + ( Xd_0__inst_mult_2_497  ))
// Xd_0__inst_mult_2_513  = CARRY(( (din_a[32] & din_b[29]) ) + ( Xd_0__inst_mult_2_498  ) + ( Xd_0__inst_mult_2_497  ))
// Xd_0__inst_mult_2_514  = SHARE((din_a[32] & din_b[30]))

	.dataa(!din_a[32]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_497 ),
	.sharein(Xd_0__inst_mult_2_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_512 ),
	.cout(Xd_0__inst_mult_2_513 ),
	.shareout(Xd_0__inst_mult_2_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_154 (
// Equation(s):
// Xd_0__inst_mult_2_516  = SUM(( (din_a[28] & din_b[33]) ) + ( Xd_0__inst_mult_2_502  ) + ( Xd_0__inst_mult_2_501  ))
// Xd_0__inst_mult_2_517  = CARRY(( (din_a[28] & din_b[33]) ) + ( Xd_0__inst_mult_2_502  ) + ( Xd_0__inst_mult_2_501  ))
// Xd_0__inst_mult_2_518  = SHARE((din_a[28] & din_b[34]))

	.dataa(!din_a[28]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_501 ),
	.sharein(Xd_0__inst_mult_2_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_516 ),
	.cout(Xd_0__inst_mult_2_517 ),
	.shareout(Xd_0__inst_mult_2_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_155 (
// Equation(s):
// Xd_0__inst_mult_2_520  = SUM(( (!din_a[30] & (((din_a[29] & din_b[32])))) # (din_a[30] & (!din_b[31] $ (((!din_a[29]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_506  ) + ( Xd_0__inst_mult_2_505  ))
// Xd_0__inst_mult_2_521  = CARRY(( (!din_a[30] & (((din_a[29] & din_b[32])))) # (din_a[30] & (!din_b[31] $ (((!din_a[29]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_506  ) + ( Xd_0__inst_mult_2_505  ))
// Xd_0__inst_mult_2_522  = SHARE((din_a[30] & (din_b[31] & (din_a[29] & din_b[32]))))

	.dataa(!din_a[30]),
	.datab(!din_b[31]),
	.datac(!din_a[29]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_505 ),
	.sharein(Xd_0__inst_mult_2_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_520 ),
	.cout(Xd_0__inst_mult_2_521 ),
	.shareout(Xd_0__inst_mult_2_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_157 (
// Equation(s):
// Xd_0__inst_mult_3_540  = SUM(( (din_a[44] & din_b[41]) ) + ( Xd_0__inst_mult_3_530  ) + ( Xd_0__inst_mult_3_529  ))
// Xd_0__inst_mult_3_541  = CARRY(( (din_a[44] & din_b[41]) ) + ( Xd_0__inst_mult_3_530  ) + ( Xd_0__inst_mult_3_529  ))
// Xd_0__inst_mult_3_542  = SHARE((din_a[44] & din_b[42]))

	.dataa(!din_a[44]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_529 ),
	.sharein(Xd_0__inst_mult_3_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_540 ),
	.cout(Xd_0__inst_mult_3_541 ),
	.shareout(Xd_0__inst_mult_3_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_158 (
// Equation(s):
// Xd_0__inst_mult_3_544  = SUM(( (!din_a[42] & (((din_a[41] & din_b[44])))) # (din_a[42] & (!din_b[43] $ (((!din_a[41]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_538  ) + ( Xd_0__inst_mult_3_537  ))
// Xd_0__inst_mult_3_545  = CARRY(( (!din_a[42] & (((din_a[41] & din_b[44])))) # (din_a[42] & (!din_b[43] $ (((!din_a[41]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_538  ) + ( Xd_0__inst_mult_3_537  ))
// Xd_0__inst_mult_3_546  = SHARE((din_a[42] & (din_b[43] & (din_a[41] & din_b[44]))))

	.dataa(!din_a[42]),
	.datab(!din_b[43]),
	.datac(!din_a[41]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_537 ),
	.sharein(Xd_0__inst_mult_3_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_544 ),
	.cout(Xd_0__inst_mult_3_545 ),
	.shareout(Xd_0__inst_mult_3_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_150 (
// Equation(s):
// Xd_0__inst_mult_0_512  = SUM(( (din_a[8] & din_b[5]) ) + ( Xd_0__inst_mult_0_502  ) + ( Xd_0__inst_mult_0_501  ))
// Xd_0__inst_mult_0_513  = CARRY(( (din_a[8] & din_b[5]) ) + ( Xd_0__inst_mult_0_502  ) + ( Xd_0__inst_mult_0_501  ))
// Xd_0__inst_mult_0_514  = SHARE((din_a[8] & din_b[6]))

	.dataa(!din_a[8]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_501 ),
	.sharein(Xd_0__inst_mult_0_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_512 ),
	.cout(Xd_0__inst_mult_0_513 ),
	.shareout(Xd_0__inst_mult_0_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_151 (
// Equation(s):
// Xd_0__inst_mult_0_516  = SUM(( (din_a[4] & din_b[9]) ) + ( Xd_0__inst_mult_0_506  ) + ( Xd_0__inst_mult_0_505  ))
// Xd_0__inst_mult_0_517  = CARRY(( (din_a[4] & din_b[9]) ) + ( Xd_0__inst_mult_0_506  ) + ( Xd_0__inst_mult_0_505  ))
// Xd_0__inst_mult_0_518  = SHARE((din_a[4] & din_b[10]))

	.dataa(!din_a[4]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_505 ),
	.sharein(Xd_0__inst_mult_0_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_516 ),
	.cout(Xd_0__inst_mult_0_517 ),
	.shareout(Xd_0__inst_mult_0_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_152 (
// Equation(s):
// Xd_0__inst_mult_0_520  = SUM(( (!din_a[6] & (((din_a[5] & din_b[8])))) # (din_a[6] & (!din_b[7] $ (((!din_a[5]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_510  ) + ( Xd_0__inst_mult_0_509  ))
// Xd_0__inst_mult_0_521  = CARRY(( (!din_a[6] & (((din_a[5] & din_b[8])))) # (din_a[6] & (!din_b[7] $ (((!din_a[5]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_510  ) + ( Xd_0__inst_mult_0_509  ))
// Xd_0__inst_mult_0_522  = SHARE((din_a[6] & (din_b[7] & (din_a[5] & din_b[8]))))

	.dataa(!din_a[6]),
	.datab(!din_b[7]),
	.datac(!din_a[5]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_509 ),
	.sharein(Xd_0__inst_mult_0_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_520 ),
	.cout(Xd_0__inst_mult_0_521 ),
	.shareout(Xd_0__inst_mult_0_522 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_148 (
// Equation(s):
// Xd_0__inst_mult_1_504  = SUM(( (din_a[21] & din_b[16]) ) + ( Xd_0__inst_mult_1_490  ) + ( Xd_0__inst_mult_1_489  ))
// Xd_0__inst_mult_1_505  = CARRY(( (din_a[21] & din_b[16]) ) + ( Xd_0__inst_mult_1_490  ) + ( Xd_0__inst_mult_1_489  ))
// Xd_0__inst_mult_1_506  = SHARE(GND)

	.dataa(!din_a[21]),
	.datab(!din_b[16]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_489 ),
	.sharein(Xd_0__inst_mult_1_490 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_504 ),
	.cout(Xd_0__inst_mult_1_505 ),
	.shareout(Xd_0__inst_mult_1_506 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_149 (
// Equation(s):
// Xd_0__inst_mult_1_508  = SUM(( (din_a[20] & din_b[17]) ) + ( Xd_0__inst_mult_1_494  ) + ( Xd_0__inst_mult_1_493  ))
// Xd_0__inst_mult_1_509  = CARRY(( (din_a[20] & din_b[17]) ) + ( Xd_0__inst_mult_1_494  ) + ( Xd_0__inst_mult_1_493  ))
// Xd_0__inst_mult_1_510  = SHARE((din_a[20] & din_b[18]))

	.dataa(!din_a[20]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_493 ),
	.sharein(Xd_0__inst_mult_1_494 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_508 ),
	.cout(Xd_0__inst_mult_1_509 ),
	.shareout(Xd_0__inst_mult_1_510 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_150 (
// Equation(s):
// Xd_0__inst_mult_1_512  = SUM(( (din_a[16] & din_b[21]) ) + ( Xd_0__inst_mult_1_498  ) + ( Xd_0__inst_mult_1_497  ))
// Xd_0__inst_mult_1_513  = CARRY(( (din_a[16] & din_b[21]) ) + ( Xd_0__inst_mult_1_498  ) + ( Xd_0__inst_mult_1_497  ))
// Xd_0__inst_mult_1_514  = SHARE((din_a[16] & din_b[22]))

	.dataa(!din_a[16]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_497 ),
	.sharein(Xd_0__inst_mult_1_498 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_512 ),
	.cout(Xd_0__inst_mult_1_513 ),
	.shareout(Xd_0__inst_mult_1_514 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_151 (
// Equation(s):
// Xd_0__inst_mult_1_516  = SUM(( (!din_a[18] & (((din_a[17] & din_b[20])))) # (din_a[18] & (!din_b[19] $ (((!din_a[17]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_502  ) + ( Xd_0__inst_mult_1_501  ))
// Xd_0__inst_mult_1_517  = CARRY(( (!din_a[18] & (((din_a[17] & din_b[20])))) # (din_a[18] & (!din_b[19] $ (((!din_a[17]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_502  ) + ( Xd_0__inst_mult_1_501  ))
// Xd_0__inst_mult_1_518  = SHARE((din_a[18] & (din_b[19] & (din_a[17] & din_b[20]))))

	.dataa(!din_a[18]),
	.datab(!din_b[19]),
	.datac(!din_a[17]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_501 ),
	.sharein(Xd_0__inst_mult_1_502 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_516 ),
	.cout(Xd_0__inst_mult_1_517 ),
	.shareout(Xd_0__inst_mult_1_518 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_157 (
// Equation(s):
// Xd_0__inst_mult_4_528  = SUM(( GND ) + ( Xd_0__inst_mult_4_514  ) + ( Xd_0__inst_mult_4_513  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_513 ),
	.sharein(Xd_0__inst_mult_4_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_528 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_158 (
// Equation(s):
// Xd_0__inst_mult_4_532  = SUM(( (din_a[57] & din_b[53]) ) + ( Xd_0__inst_mult_4_518  ) + ( Xd_0__inst_mult_4_517  ))
// Xd_0__inst_mult_4_533  = CARRY(( (din_a[57] & din_b[53]) ) + ( Xd_0__inst_mult_4_518  ) + ( Xd_0__inst_mult_4_517  ))
// Xd_0__inst_mult_4_534  = SHARE((din_a[57] & din_b[54]))

	.dataa(!din_a[57]),
	.datab(!din_b[53]),
	.datac(!din_b[54]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_517 ),
	.sharein(Xd_0__inst_mult_4_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_532 ),
	.cout(Xd_0__inst_mult_4_533 ),
	.shareout(Xd_0__inst_mult_4_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_159 (
// Equation(s):
// Xd_0__inst_mult_4_536  = SUM(( (din_a[53] & din_b[57]) ) + ( Xd_0__inst_mult_4_522  ) + ( Xd_0__inst_mult_4_521  ))
// Xd_0__inst_mult_4_537  = CARRY(( (din_a[53] & din_b[57]) ) + ( Xd_0__inst_mult_4_522  ) + ( Xd_0__inst_mult_4_521  ))
// Xd_0__inst_mult_4_538  = SHARE((din_a[53] & din_b[58]))

	.dataa(!din_a[53]),
	.datab(!din_b[57]),
	.datac(!din_b[58]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_521 ),
	.sharein(Xd_0__inst_mult_4_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_536 ),
	.cout(Xd_0__inst_mult_4_537 ),
	.shareout(Xd_0__inst_mult_4_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_160 (
// Equation(s):
// Xd_0__inst_mult_4_540  = SUM(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_526  ) + ( Xd_0__inst_mult_4_525  ))
// Xd_0__inst_mult_4_541  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[56])))) # (din_a[55] & (!din_b[55] $ (((!din_a[54]) # (!din_b[56]))))) ) + ( Xd_0__inst_mult_4_526  ) + ( Xd_0__inst_mult_4_525  ))
// Xd_0__inst_mult_4_542  = SHARE((din_a[55] & (din_b[55] & (din_a[54] & din_b[56]))))

	.dataa(!din_a[55]),
	.datab(!din_b[55]),
	.datac(!din_a[54]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_525 ),
	.sharein(Xd_0__inst_mult_4_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_540 ),
	.cout(Xd_0__inst_mult_4_541 ),
	.shareout(Xd_0__inst_mult_4_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_156 (
// Equation(s):
// Xd_0__inst_mult_5_524  = SUM(( GND ) + ( Xd_0__inst_mult_5_510  ) + ( Xd_0__inst_mult_5_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_509 ),
	.sharein(Xd_0__inst_mult_5_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_524 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_157 (
// Equation(s):
// Xd_0__inst_mult_5_528  = SUM(( (din_a[69] & din_b[65]) ) + ( Xd_0__inst_mult_5_514  ) + ( Xd_0__inst_mult_5_513  ))
// Xd_0__inst_mult_5_529  = CARRY(( (din_a[69] & din_b[65]) ) + ( Xd_0__inst_mult_5_514  ) + ( Xd_0__inst_mult_5_513  ))
// Xd_0__inst_mult_5_530  = SHARE((din_a[69] & din_b[66]))

	.dataa(!din_a[69]),
	.datab(!din_b[65]),
	.datac(!din_b[66]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_513 ),
	.sharein(Xd_0__inst_mult_5_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_528 ),
	.cout(Xd_0__inst_mult_5_529 ),
	.shareout(Xd_0__inst_mult_5_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_158 (
// Equation(s):
// Xd_0__inst_mult_5_532  = SUM(( (din_a[65] & din_b[69]) ) + ( Xd_0__inst_mult_5_518  ) + ( Xd_0__inst_mult_5_517  ))
// Xd_0__inst_mult_5_533  = CARRY(( (din_a[65] & din_b[69]) ) + ( Xd_0__inst_mult_5_518  ) + ( Xd_0__inst_mult_5_517  ))
// Xd_0__inst_mult_5_534  = SHARE((din_a[65] & din_b[70]))

	.dataa(!din_a[65]),
	.datab(!din_b[69]),
	.datac(!din_b[70]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_517 ),
	.sharein(Xd_0__inst_mult_5_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_532 ),
	.cout(Xd_0__inst_mult_5_533 ),
	.shareout(Xd_0__inst_mult_5_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_159 (
// Equation(s):
// Xd_0__inst_mult_5_536  = SUM(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_522  ) + ( Xd_0__inst_mult_5_521  ))
// Xd_0__inst_mult_5_537  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[68])))) # (din_a[67] & (!din_b[67] $ (((!din_a[66]) # (!din_b[68]))))) ) + ( Xd_0__inst_mult_5_522  ) + ( Xd_0__inst_mult_5_521  ))
// Xd_0__inst_mult_5_538  = SHARE((din_a[67] & (din_b[67] & (din_a[66] & din_b[68]))))

	.dataa(!din_a[67]),
	.datab(!din_b[67]),
	.datac(!din_a[66]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_521 ),
	.sharein(Xd_0__inst_mult_5_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_536 ),
	.cout(Xd_0__inst_mult_5_537 ),
	.shareout(Xd_0__inst_mult_5_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_156 (
// Equation(s):
// Xd_0__inst_mult_2_524  = SUM(( GND ) + ( Xd_0__inst_mult_2_510  ) + ( Xd_0__inst_mult_2_509  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_509 ),
	.sharein(Xd_0__inst_mult_2_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_524 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_157 (
// Equation(s):
// Xd_0__inst_mult_2_528  = SUM(( (din_a[33] & din_b[29]) ) + ( Xd_0__inst_mult_2_514  ) + ( Xd_0__inst_mult_2_513  ))
// Xd_0__inst_mult_2_529  = CARRY(( (din_a[33] & din_b[29]) ) + ( Xd_0__inst_mult_2_514  ) + ( Xd_0__inst_mult_2_513  ))
// Xd_0__inst_mult_2_530  = SHARE((din_a[33] & din_b[30]))

	.dataa(!din_a[33]),
	.datab(!din_b[29]),
	.datac(!din_b[30]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_513 ),
	.sharein(Xd_0__inst_mult_2_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_528 ),
	.cout(Xd_0__inst_mult_2_529 ),
	.shareout(Xd_0__inst_mult_2_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_158 (
// Equation(s):
// Xd_0__inst_mult_2_532  = SUM(( (din_a[29] & din_b[33]) ) + ( Xd_0__inst_mult_2_518  ) + ( Xd_0__inst_mult_2_517  ))
// Xd_0__inst_mult_2_533  = CARRY(( (din_a[29] & din_b[33]) ) + ( Xd_0__inst_mult_2_518  ) + ( Xd_0__inst_mult_2_517  ))
// Xd_0__inst_mult_2_534  = SHARE((din_a[29] & din_b[34]))

	.dataa(!din_a[29]),
	.datab(!din_b[33]),
	.datac(!din_b[34]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_517 ),
	.sharein(Xd_0__inst_mult_2_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_532 ),
	.cout(Xd_0__inst_mult_2_533 ),
	.shareout(Xd_0__inst_mult_2_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_159 (
// Equation(s):
// Xd_0__inst_mult_2_536  = SUM(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_522  ) + ( Xd_0__inst_mult_2_521  ))
// Xd_0__inst_mult_2_537  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[32])))) # (din_a[31] & (!din_b[31] $ (((!din_a[30]) # (!din_b[32]))))) ) + ( Xd_0__inst_mult_2_522  ) + ( Xd_0__inst_mult_2_521  ))
// Xd_0__inst_mult_2_538  = SHARE((din_a[31] & (din_b[31] & (din_a[30] & din_b[32]))))

	.dataa(!din_a[31]),
	.datab(!din_b[31]),
	.datac(!din_a[30]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_521 ),
	.sharein(Xd_0__inst_mult_2_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_536 ),
	.cout(Xd_0__inst_mult_2_537 ),
	.shareout(Xd_0__inst_mult_2_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_159 (
// Equation(s):
// Xd_0__inst_mult_3_548  = SUM(( (din_a[45] & din_b[41]) ) + ( Xd_0__inst_mult_3_542  ) + ( Xd_0__inst_mult_3_541  ))
// Xd_0__inst_mult_3_549  = CARRY(( (din_a[45] & din_b[41]) ) + ( Xd_0__inst_mult_3_542  ) + ( Xd_0__inst_mult_3_541  ))
// Xd_0__inst_mult_3_550  = SHARE((din_a[45] & din_b[42]))

	.dataa(!din_a[45]),
	.datab(!din_b[41]),
	.datac(!din_b[42]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_541 ),
	.sharein(Xd_0__inst_mult_3_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_548 ),
	.cout(Xd_0__inst_mult_3_549 ),
	.shareout(Xd_0__inst_mult_3_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_3_160 (
// Equation(s):
// Xd_0__inst_mult_3_552  = SUM(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_546  ) + ( Xd_0__inst_mult_3_545  ))
// Xd_0__inst_mult_3_553  = CARRY(( (!din_a[43] & (((din_a[42] & din_b[44])))) # (din_a[43] & (!din_b[43] $ (((!din_a[42]) # (!din_b[44]))))) ) + ( Xd_0__inst_mult_3_546  ) + ( Xd_0__inst_mult_3_545  ))
// Xd_0__inst_mult_3_554  = SHARE((din_a[43] & (din_b[43] & (din_a[42] & din_b[44]))))

	.dataa(!din_a[43]),
	.datab(!din_b[43]),
	.datac(!din_a[42]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_545 ),
	.sharein(Xd_0__inst_mult_3_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_552 ),
	.cout(Xd_0__inst_mult_3_553 ),
	.shareout(Xd_0__inst_mult_3_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_153 (
// Equation(s):
// Xd_0__inst_mult_0_524  = SUM(( (din_a[9] & din_b[5]) ) + ( Xd_0__inst_mult_0_514  ) + ( Xd_0__inst_mult_0_513  ))
// Xd_0__inst_mult_0_525  = CARRY(( (din_a[9] & din_b[5]) ) + ( Xd_0__inst_mult_0_514  ) + ( Xd_0__inst_mult_0_513  ))
// Xd_0__inst_mult_0_526  = SHARE((din_a[9] & din_b[6]))

	.dataa(!din_a[9]),
	.datab(!din_b[5]),
	.datac(!din_b[6]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_513 ),
	.sharein(Xd_0__inst_mult_0_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_524 ),
	.cout(Xd_0__inst_mult_0_525 ),
	.shareout(Xd_0__inst_mult_0_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_154 (
// Equation(s):
// Xd_0__inst_mult_0_528  = SUM(( (din_a[5] & din_b[9]) ) + ( Xd_0__inst_mult_0_518  ) + ( Xd_0__inst_mult_0_517  ))
// Xd_0__inst_mult_0_529  = CARRY(( (din_a[5] & din_b[9]) ) + ( Xd_0__inst_mult_0_518  ) + ( Xd_0__inst_mult_0_517  ))
// Xd_0__inst_mult_0_530  = SHARE((din_a[5] & din_b[10]))

	.dataa(!din_a[5]),
	.datab(!din_b[9]),
	.datac(!din_b[10]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_517 ),
	.sharein(Xd_0__inst_mult_0_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_528 ),
	.cout(Xd_0__inst_mult_0_529 ),
	.shareout(Xd_0__inst_mult_0_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_155 (
// Equation(s):
// Xd_0__inst_mult_0_532  = SUM(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_522  ) + ( Xd_0__inst_mult_0_521  ))
// Xd_0__inst_mult_0_533  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[8])))) # (din_a[7] & (!din_b[7] $ (((!din_a[6]) # (!din_b[8]))))) ) + ( Xd_0__inst_mult_0_522  ) + ( Xd_0__inst_mult_0_521  ))
// Xd_0__inst_mult_0_534  = SHARE((din_a[7] & (din_b[7] & (din_a[6] & din_b[8]))))

	.dataa(!din_a[7]),
	.datab(!din_b[7]),
	.datac(!din_a[6]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_521 ),
	.sharein(Xd_0__inst_mult_0_522 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_532 ),
	.cout(Xd_0__inst_mult_0_533 ),
	.shareout(Xd_0__inst_mult_0_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_152 (
// Equation(s):
// Xd_0__inst_mult_1_520  = SUM(( GND ) + ( Xd_0__inst_mult_1_506  ) + ( Xd_0__inst_mult_1_505  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_505 ),
	.sharein(Xd_0__inst_mult_1_506 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_520 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_153 (
// Equation(s):
// Xd_0__inst_mult_1_524  = SUM(( (din_a[21] & din_b[17]) ) + ( Xd_0__inst_mult_1_510  ) + ( Xd_0__inst_mult_1_509  ))
// Xd_0__inst_mult_1_525  = CARRY(( (din_a[21] & din_b[17]) ) + ( Xd_0__inst_mult_1_510  ) + ( Xd_0__inst_mult_1_509  ))
// Xd_0__inst_mult_1_526  = SHARE((din_a[21] & din_b[18]))

	.dataa(!din_a[21]),
	.datab(!din_b[17]),
	.datac(!din_b[18]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_509 ),
	.sharein(Xd_0__inst_mult_1_510 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_524 ),
	.cout(Xd_0__inst_mult_1_525 ),
	.shareout(Xd_0__inst_mult_1_526 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000050500001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_154 (
// Equation(s):
// Xd_0__inst_mult_1_528  = SUM(( (din_a[17] & din_b[21]) ) + ( Xd_0__inst_mult_1_514  ) + ( Xd_0__inst_mult_1_513  ))
// Xd_0__inst_mult_1_529  = CARRY(( (din_a[17] & din_b[21]) ) + ( Xd_0__inst_mult_1_514  ) + ( Xd_0__inst_mult_1_513  ))
// Xd_0__inst_mult_1_530  = SHARE((din_a[17] & din_b[22]))

	.dataa(!din_a[17]),
	.datab(!din_b[21]),
	.datac(!din_b[22]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_513 ),
	.sharein(Xd_0__inst_mult_1_514 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_528 ),
	.cout(Xd_0__inst_mult_1_529 ),
	.shareout(Xd_0__inst_mult_1_530 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_155 (
// Equation(s):
// Xd_0__inst_mult_1_532  = SUM(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_518  ) + ( Xd_0__inst_mult_1_517  ))
// Xd_0__inst_mult_1_533  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[20])))) # (din_a[19] & (!din_b[19] $ (((!din_a[18]) # (!din_b[20]))))) ) + ( Xd_0__inst_mult_1_518  ) + ( Xd_0__inst_mult_1_517  ))
// Xd_0__inst_mult_1_534  = SHARE((din_a[19] & (din_b[19] & (din_a[18] & din_b[20]))))

	.dataa(!din_a[19]),
	.datab(!din_b[19]),
	.datac(!din_a[18]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_517 ),
	.sharein(Xd_0__inst_mult_1_518 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_532 ),
	.cout(Xd_0__inst_mult_1_533 ),
	.shareout(Xd_0__inst_mult_1_534 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_161 (
// Equation(s):
// Xd_0__inst_mult_4_544  = SUM(( (din_a[56] & din_b[55]) ) + ( Xd_0__inst_mult_4_534  ) + ( Xd_0__inst_mult_4_533  ))
// Xd_0__inst_mult_4_545  = CARRY(( (din_a[56] & din_b[55]) ) + ( Xd_0__inst_mult_4_534  ) + ( Xd_0__inst_mult_4_533  ))
// Xd_0__inst_mult_4_546  = SHARE((din_b[55] & din_a[57]))

	.dataa(!din_a[56]),
	.datab(!din_b[55]),
	.datac(!din_a[57]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_533 ),
	.sharein(Xd_0__inst_mult_4_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_544 ),
	.cout(Xd_0__inst_mult_4_545 ),
	.shareout(Xd_0__inst_mult_4_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_162 (
// Equation(s):
// Xd_0__inst_mult_4_548  = SUM(( (!din_a[55] & (((din_a[54] & din_b[57])))) # (din_a[55] & (!din_b[56] $ (((!din_a[54]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_4_538  ) + ( Xd_0__inst_mult_4_537  ))
// Xd_0__inst_mult_4_549  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[57])))) # (din_a[55] & (!din_b[56] $ (((!din_a[54]) # (!din_b[57]))))) ) + ( Xd_0__inst_mult_4_538  ) + ( Xd_0__inst_mult_4_537  ))
// Xd_0__inst_mult_4_550  = SHARE((din_a[55] & (din_b[56] & (din_a[54] & din_b[57]))))

	.dataa(!din_a[55]),
	.datab(!din_b[56]),
	.datac(!din_a[54]),
	.datad(!din_b[57]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_537 ),
	.sharein(Xd_0__inst_mult_4_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_548 ),
	.cout(Xd_0__inst_mult_4_549 ),
	.shareout(Xd_0__inst_mult_4_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_160 (
// Equation(s):
// Xd_0__inst_mult_5_540  = SUM(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_5_530  ) + ( Xd_0__inst_mult_5_529  ))
// Xd_0__inst_mult_5_541  = CARRY(( (din_a[68] & din_b[67]) ) + ( Xd_0__inst_mult_5_530  ) + ( Xd_0__inst_mult_5_529  ))
// Xd_0__inst_mult_5_542  = SHARE((din_b[67] & din_a[69]))

	.dataa(!din_a[68]),
	.datab(!din_b[67]),
	.datac(!din_a[69]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_529 ),
	.sharein(Xd_0__inst_mult_5_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_540 ),
	.cout(Xd_0__inst_mult_5_541 ),
	.shareout(Xd_0__inst_mult_5_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_161 (
// Equation(s):
// Xd_0__inst_mult_5_544  = SUM(( (!din_a[67] & (((din_a[66] & din_b[69])))) # (din_a[67] & (!din_b[68] $ (((!din_a[66]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_5_534  ) + ( Xd_0__inst_mult_5_533  ))
// Xd_0__inst_mult_5_545  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[69])))) # (din_a[67] & (!din_b[68] $ (((!din_a[66]) # (!din_b[69]))))) ) + ( Xd_0__inst_mult_5_534  ) + ( Xd_0__inst_mult_5_533  ))
// Xd_0__inst_mult_5_546  = SHARE((din_a[67] & (din_b[68] & (din_a[66] & din_b[69]))))

	.dataa(!din_a[67]),
	.datab(!din_b[68]),
	.datac(!din_a[66]),
	.datad(!din_b[69]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_533 ),
	.sharein(Xd_0__inst_mult_5_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_544 ),
	.cout(Xd_0__inst_mult_5_545 ),
	.shareout(Xd_0__inst_mult_5_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_162 (
// Equation(s):
// Xd_0__inst_mult_5_548  = SUM(( GND ) + ( Xd_0__inst_mult_5_538  ) + ( Xd_0__inst_mult_5_537  ))
// Xd_0__inst_mult_5_549  = CARRY(( GND ) + ( Xd_0__inst_mult_5_538  ) + ( Xd_0__inst_mult_5_537  ))
// Xd_0__inst_mult_5_550  = SHARE(VCC)

	.dataa(!din_a[62]),
	.datab(!din_b[67]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_537 ),
	.sharein(Xd_0__inst_mult_5_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_548 ),
	.cout(Xd_0__inst_mult_5_549 ),
	.shareout(Xd_0__inst_mult_5_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_160 (
// Equation(s):
// Xd_0__inst_mult_2_540  = SUM(( (din_a[32] & din_b[31]) ) + ( Xd_0__inst_mult_2_530  ) + ( Xd_0__inst_mult_2_529  ))
// Xd_0__inst_mult_2_541  = CARRY(( (din_a[32] & din_b[31]) ) + ( Xd_0__inst_mult_2_530  ) + ( Xd_0__inst_mult_2_529  ))
// Xd_0__inst_mult_2_542  = SHARE((din_b[31] & din_a[33]))

	.dataa(!din_a[32]),
	.datab(!din_b[31]),
	.datac(!din_a[33]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_529 ),
	.sharein(Xd_0__inst_mult_2_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_540 ),
	.cout(Xd_0__inst_mult_2_541 ),
	.shareout(Xd_0__inst_mult_2_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_161 (
// Equation(s):
// Xd_0__inst_mult_2_544  = SUM(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_2_534  ) + ( Xd_0__inst_mult_2_533  ))
// Xd_0__inst_mult_2_545  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[33])))) # (din_a[31] & (!din_b[32] $ (((!din_a[30]) # (!din_b[33]))))) ) + ( Xd_0__inst_mult_2_534  ) + ( Xd_0__inst_mult_2_533  ))
// Xd_0__inst_mult_2_546  = SHARE((din_a[31] & (din_b[32] & (din_a[30] & din_b[33]))))

	.dataa(!din_a[31]),
	.datab(!din_b[32]),
	.datac(!din_a[30]),
	.datad(!din_b[33]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_533 ),
	.sharein(Xd_0__inst_mult_2_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_544 ),
	.cout(Xd_0__inst_mult_2_545 ),
	.shareout(Xd_0__inst_mult_2_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_156 (
// Equation(s):
// Xd_0__inst_mult_1_536  = SUM(( GND ) + ( Xd_0__inst_mult_2_538  ) + ( Xd_0__inst_mult_2_537  ))
// Xd_0__inst_mult_1_537  = CARRY(( GND ) + ( Xd_0__inst_mult_2_538  ) + ( Xd_0__inst_mult_2_537  ))
// Xd_0__inst_mult_1_538  = SHARE(VCC)

	.dataa(!din_a[14]),
	.datab(!din_b[19]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_537 ),
	.sharein(Xd_0__inst_mult_2_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_536 ),
	.cout(Xd_0__inst_mult_1_537 ),
	.shareout(Xd_0__inst_mult_1_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_161 (
// Equation(s):
// Xd_0__inst_mult_3_556  = SUM(( (din_a[44] & din_b[43]) ) + ( Xd_0__inst_mult_3_550  ) + ( Xd_0__inst_mult_3_549  ))
// Xd_0__inst_mult_3_557  = CARRY(( (din_a[44] & din_b[43]) ) + ( Xd_0__inst_mult_3_550  ) + ( Xd_0__inst_mult_3_549  ))
// Xd_0__inst_mult_3_558  = SHARE((din_b[43] & din_a[45]))

	.dataa(!din_a[44]),
	.datab(!din_b[43]),
	.datac(!din_a[45]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_549 ),
	.sharein(Xd_0__inst_mult_3_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_556 ),
	.cout(Xd_0__inst_mult_3_557 ),
	.shareout(Xd_0__inst_mult_3_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_162 (
// Equation(s):
// Xd_0__inst_mult_2_548  = SUM(( GND ) + ( Xd_0__inst_mult_3_554  ) + ( Xd_0__inst_mult_3_553  ))
// Xd_0__inst_mult_2_549  = CARRY(( GND ) + ( Xd_0__inst_mult_3_554  ) + ( Xd_0__inst_mult_3_553  ))
// Xd_0__inst_mult_2_550  = SHARE(VCC)

	.dataa(!din_a[26]),
	.datab(!din_b[31]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_553 ),
	.sharein(Xd_0__inst_mult_3_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_548 ),
	.cout(Xd_0__inst_mult_2_549 ),
	.shareout(Xd_0__inst_mult_2_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_156 (
// Equation(s):
// Xd_0__inst_mult_0_536  = SUM(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_0_526  ) + ( Xd_0__inst_mult_0_525  ))
// Xd_0__inst_mult_0_537  = CARRY(( (din_a[8] & din_b[7]) ) + ( Xd_0__inst_mult_0_526  ) + ( Xd_0__inst_mult_0_525  ))
// Xd_0__inst_mult_0_538  = SHARE((din_b[7] & din_a[9]))

	.dataa(!din_a[8]),
	.datab(!din_b[7]),
	.datac(!din_a[9]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_525 ),
	.sharein(Xd_0__inst_mult_0_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_536 ),
	.cout(Xd_0__inst_mult_0_537 ),
	.shareout(Xd_0__inst_mult_0_538 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_157 (
// Equation(s):
// Xd_0__inst_mult_0_540  = SUM(( (!din_a[7] & (((din_a[6] & din_b[9])))) # (din_a[7] & (!din_b[8] $ (((!din_a[6]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_0_530  ) + ( Xd_0__inst_mult_0_529  ))
// Xd_0__inst_mult_0_541  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[9])))) # (din_a[7] & (!din_b[8] $ (((!din_a[6]) # (!din_b[9]))))) ) + ( Xd_0__inst_mult_0_530  ) + ( Xd_0__inst_mult_0_529  ))
// Xd_0__inst_mult_0_542  = SHARE((din_a[7] & (din_b[8] & (din_a[6] & din_b[9]))))

	.dataa(!din_a[7]),
	.datab(!din_b[8]),
	.datac(!din_a[6]),
	.datad(!din_b[9]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_529 ),
	.sharein(Xd_0__inst_mult_0_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_540 ),
	.cout(Xd_0__inst_mult_0_541 ),
	.shareout(Xd_0__inst_mult_0_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_158 (
// Equation(s):
// Xd_0__inst_mult_0_544  = SUM(( GND ) + ( Xd_0__inst_mult_0_534  ) + ( Xd_0__inst_mult_0_533  ))
// Xd_0__inst_mult_0_545  = CARRY(( GND ) + ( Xd_0__inst_mult_0_534  ) + ( Xd_0__inst_mult_0_533  ))
// Xd_0__inst_mult_0_546  = SHARE(VCC)

	.dataa(!din_a[2]),
	.datab(!din_b[7]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_533 ),
	.sharein(Xd_0__inst_mult_0_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_544 ),
	.cout(Xd_0__inst_mult_0_545 ),
	.shareout(Xd_0__inst_mult_0_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000030300001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_157 (
// Equation(s):
// Xd_0__inst_mult_1_540  = SUM(( (din_a[20] & din_b[19]) ) + ( Xd_0__inst_mult_1_526  ) + ( Xd_0__inst_mult_1_525  ))
// Xd_0__inst_mult_1_541  = CARRY(( (din_a[20] & din_b[19]) ) + ( Xd_0__inst_mult_1_526  ) + ( Xd_0__inst_mult_1_525  ))
// Xd_0__inst_mult_1_542  = SHARE((din_b[19] & din_a[21]))

	.dataa(!din_a[20]),
	.datab(!din_b[19]),
	.datac(!din_a[21]),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_525 ),
	.sharein(Xd_0__inst_mult_1_526 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_540 ),
	.cout(Xd_0__inst_mult_1_541 ),
	.shareout(Xd_0__inst_mult_1_542 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_158 (
// Equation(s):
// Xd_0__inst_mult_1_544  = SUM(( (!din_a[19] & (((din_a[18] & din_b[21])))) # (din_a[19] & (!din_b[20] $ (((!din_a[18]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_1_530  ) + ( Xd_0__inst_mult_1_529  ))
// Xd_0__inst_mult_1_545  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[21])))) # (din_a[19] & (!din_b[20] $ (((!din_a[18]) # (!din_b[21]))))) ) + ( Xd_0__inst_mult_1_530  ) + ( Xd_0__inst_mult_1_529  ))
// Xd_0__inst_mult_1_546  = SHARE((din_a[19] & (din_b[20] & (din_a[18] & din_b[21]))))

	.dataa(!din_a[19]),
	.datab(!din_b[20]),
	.datac(!din_a[18]),
	.datad(!din_b[21]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_529 ),
	.sharein(Xd_0__inst_mult_1_530 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_544 ),
	.cout(Xd_0__inst_mult_1_545 ),
	.shareout(Xd_0__inst_mult_1_546 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000FFFF00000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_159 (
// Equation(s):
// Xd_0__inst_mult_1_548  = SUM(( GND ) + ( Xd_0__inst_mult_1_534  ) + ( Xd_0__inst_mult_1_533  ))
// Xd_0__inst_mult_1_549  = CARRY(( GND ) + ( Xd_0__inst_mult_1_534  ) + ( Xd_0__inst_mult_1_533  ))
// Xd_0__inst_mult_1_550  = SHARE(VCC)

	.dataa(!din_a[15]),
	.datab(!din_b[13]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_533 ),
	.sharein(Xd_0__inst_mult_1_534 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_548 ),
	.cout(Xd_0__inst_mult_1_549 ),
	.shareout(Xd_0__inst_mult_1_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_163 (
// Equation(s):
// Xd_0__inst_mult_4_552  = SUM(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_4_546  ) + ( Xd_0__inst_mult_4_545  ))
// Xd_0__inst_mult_4_553  = CARRY(( (din_a[56] & din_b[56]) ) + ( Xd_0__inst_mult_4_546  ) + ( Xd_0__inst_mult_4_545  ))
// Xd_0__inst_mult_4_554  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[56]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_545 ),
	.sharein(Xd_0__inst_mult_4_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_552 ),
	.cout(Xd_0__inst_mult_4_553 ),
	.shareout(Xd_0__inst_mult_4_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_164 (
// Equation(s):
// Xd_0__inst_mult_4_556  = SUM(( (!din_a[55] & (((din_a[54] & din_b[58])))) # (din_a[55] & (!din_b[57] $ (((!din_a[54]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_550  ) + ( Xd_0__inst_mult_4_549  ))
// Xd_0__inst_mult_4_557  = CARRY(( (!din_a[55] & (((din_a[54] & din_b[58])))) # (din_a[55] & (!din_b[57] $ (((!din_a[54]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_550  ) + ( Xd_0__inst_mult_4_549  ))
// Xd_0__inst_mult_4_558  = SHARE((din_a[55] & (din_b[57] & (din_a[54] & din_b[58]))))

	.dataa(!din_a[55]),
	.datab(!din_b[57]),
	.datac(!din_a[54]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_549 ),
	.sharein(Xd_0__inst_mult_4_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_556 ),
	.cout(Xd_0__inst_mult_4_557 ),
	.shareout(Xd_0__inst_mult_4_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_163 (
// Equation(s):
// Xd_0__inst_mult_5_552  = SUM(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_5_542  ) + ( Xd_0__inst_mult_5_541  ))
// Xd_0__inst_mult_5_553  = CARRY(( (din_a[68] & din_b[68]) ) + ( Xd_0__inst_mult_5_542  ) + ( Xd_0__inst_mult_5_541  ))
// Xd_0__inst_mult_5_554  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[68]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_541 ),
	.sharein(Xd_0__inst_mult_5_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_552 ),
	.cout(Xd_0__inst_mult_5_553 ),
	.shareout(Xd_0__inst_mult_5_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_164 (
// Equation(s):
// Xd_0__inst_mult_5_556  = SUM(( (!din_a[67] & (((din_a[66] & din_b[70])))) # (din_a[67] & (!din_b[69] $ (((!din_a[66]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_546  ) + ( Xd_0__inst_mult_5_545  ))
// Xd_0__inst_mult_5_557  = CARRY(( (!din_a[67] & (((din_a[66] & din_b[70])))) # (din_a[67] & (!din_b[69] $ (((!din_a[66]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_546  ) + ( Xd_0__inst_mult_5_545  ))
// Xd_0__inst_mult_5_558  = SHARE((din_a[67] & (din_b[69] & (din_a[66] & din_b[70]))))

	.dataa(!din_a[67]),
	.datab(!din_b[69]),
	.datac(!din_a[66]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_545 ),
	.sharein(Xd_0__inst_mult_5_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_556 ),
	.cout(Xd_0__inst_mult_5_557 ),
	.shareout(Xd_0__inst_mult_5_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_163 (
// Equation(s):
// Xd_0__inst_mult_2_552  = SUM(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_2_542  ) + ( Xd_0__inst_mult_2_541  ))
// Xd_0__inst_mult_2_553  = CARRY(( (din_a[32] & din_b[32]) ) + ( Xd_0__inst_mult_2_542  ) + ( Xd_0__inst_mult_2_541  ))
// Xd_0__inst_mult_2_554  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[32]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_541 ),
	.sharein(Xd_0__inst_mult_2_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_552 ),
	.cout(Xd_0__inst_mult_2_553 ),
	.shareout(Xd_0__inst_mult_2_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_164 (
// Equation(s):
// Xd_0__inst_mult_2_556  = SUM(( (!din_a[31] & (((din_a[30] & din_b[34])))) # (din_a[31] & (!din_b[33] $ (((!din_a[30]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_546  ) + ( Xd_0__inst_mult_2_545  ))
// Xd_0__inst_mult_2_557  = CARRY(( (!din_a[31] & (((din_a[30] & din_b[34])))) # (din_a[31] & (!din_b[33] $ (((!din_a[30]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_546  ) + ( Xd_0__inst_mult_2_545  ))
// Xd_0__inst_mult_2_558  = SHARE((din_a[31] & (din_b[33] & (din_a[30] & din_b[34]))))

	.dataa(!din_a[31]),
	.datab(!din_b[33]),
	.datac(!din_a[30]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_545 ),
	.sharein(Xd_0__inst_mult_2_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_556 ),
	.cout(Xd_0__inst_mult_2_557 ),
	.shareout(Xd_0__inst_mult_2_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_162 (
// Equation(s):
// Xd_0__inst_mult_3_560  = SUM(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_3_558  ) + ( Xd_0__inst_mult_3_557  ))
// Xd_0__inst_mult_3_561  = CARRY(( (din_a[44] & din_b[44]) ) + ( Xd_0__inst_mult_3_558  ) + ( Xd_0__inst_mult_3_557  ))
// Xd_0__inst_mult_3_562  = SHARE(GND)

	.dataa(!din_a[44]),
	.datab(!din_b[44]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_557 ),
	.sharein(Xd_0__inst_mult_3_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_560 ),
	.cout(Xd_0__inst_mult_3_561 ),
	.shareout(Xd_0__inst_mult_3_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_159 (
// Equation(s):
// Xd_0__inst_mult_0_548  = SUM(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_0_538  ) + ( Xd_0__inst_mult_0_537  ))
// Xd_0__inst_mult_0_549  = CARRY(( (din_a[8] & din_b[8]) ) + ( Xd_0__inst_mult_0_538  ) + ( Xd_0__inst_mult_0_537  ))
// Xd_0__inst_mult_0_550  = SHARE(GND)

	.dataa(!din_a[8]),
	.datab(!din_b[8]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_537 ),
	.sharein(Xd_0__inst_mult_0_538 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_548 ),
	.cout(Xd_0__inst_mult_0_549 ),
	.shareout(Xd_0__inst_mult_0_550 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_160 (
// Equation(s):
// Xd_0__inst_mult_0_552  = SUM(( (!din_a[7] & (((din_a[6] & din_b[10])))) # (din_a[7] & (!din_b[9] $ (((!din_a[6]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_542  ) + ( Xd_0__inst_mult_0_541  ))
// Xd_0__inst_mult_0_553  = CARRY(( (!din_a[7] & (((din_a[6] & din_b[10])))) # (din_a[7] & (!din_b[9] $ (((!din_a[6]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_542  ) + ( Xd_0__inst_mult_0_541  ))
// Xd_0__inst_mult_0_554  = SHARE((din_a[7] & (din_b[9] & (din_a[6] & din_b[10]))))

	.dataa(!din_a[7]),
	.datab(!din_b[9]),
	.datac(!din_a[6]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_541 ),
	.sharein(Xd_0__inst_mult_0_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_552 ),
	.cout(Xd_0__inst_mult_0_553 ),
	.shareout(Xd_0__inst_mult_0_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_160 (
// Equation(s):
// Xd_0__inst_mult_1_552  = SUM(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_1_542  ) + ( Xd_0__inst_mult_1_541  ))
// Xd_0__inst_mult_1_553  = CARRY(( (din_a[20] & din_b[20]) ) + ( Xd_0__inst_mult_1_542  ) + ( Xd_0__inst_mult_1_541  ))
// Xd_0__inst_mult_1_554  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[20]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_541 ),
	.sharein(Xd_0__inst_mult_1_542 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_552 ),
	.cout(Xd_0__inst_mult_1_553 ),
	.shareout(Xd_0__inst_mult_1_554 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_161 (
// Equation(s):
// Xd_0__inst_mult_1_556  = SUM(( (!din_a[19] & (((din_a[18] & din_b[22])))) # (din_a[19] & (!din_b[21] $ (((!din_a[18]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_546  ) + ( Xd_0__inst_mult_1_545  ))
// Xd_0__inst_mult_1_557  = CARRY(( (!din_a[19] & (((din_a[18] & din_b[22])))) # (din_a[19] & (!din_b[21] $ (((!din_a[18]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_546  ) + ( Xd_0__inst_mult_1_545  ))
// Xd_0__inst_mult_1_558  = SHARE((din_a[19] & (din_b[21] & (din_a[18] & din_b[22]))))

	.dataa(!din_a[19]),
	.datab(!din_b[21]),
	.datac(!din_a[18]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_545 ),
	.sharein(Xd_0__inst_mult_1_546 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_556 ),
	.cout(Xd_0__inst_mult_1_557 ),
	.shareout(Xd_0__inst_mult_1_558 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_165 (
// Equation(s):
// Xd_0__inst_mult_4_560  = SUM(( GND ) + ( Xd_0__inst_mult_4_554  ) + ( Xd_0__inst_mult_4_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_553 ),
	.sharein(Xd_0__inst_mult_4_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_4_166 (
// Equation(s):
// Xd_0__inst_mult_4_564  = SUM(( (!din_a[56] & (((din_a[55] & din_b[58])))) # (din_a[56] & (!din_b[57] $ (((!din_a[55]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_558  ) + ( Xd_0__inst_mult_4_557  ))
// Xd_0__inst_mult_4_565  = CARRY(( (!din_a[56] & (((din_a[55] & din_b[58])))) # (din_a[56] & (!din_b[57] $ (((!din_a[55]) # (!din_b[58]))))) ) + ( Xd_0__inst_mult_4_558  ) + ( Xd_0__inst_mult_4_557  ))
// Xd_0__inst_mult_4_566  = SHARE((din_a[56] & (din_b[57] & (din_a[55] & din_b[58]))))

	.dataa(!din_a[56]),
	.datab(!din_b[57]),
	.datac(!din_a[55]),
	.datad(!din_b[58]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_557 ),
	.sharein(Xd_0__inst_mult_4_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_564 ),
	.cout(Xd_0__inst_mult_4_565 ),
	.shareout(Xd_0__inst_mult_4_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_165 (
// Equation(s):
// Xd_0__inst_mult_5_560  = SUM(( GND ) + ( Xd_0__inst_mult_5_554  ) + ( Xd_0__inst_mult_5_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_553 ),
	.sharein(Xd_0__inst_mult_5_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_5_166 (
// Equation(s):
// Xd_0__inst_mult_5_564  = SUM(( (!din_a[68] & (((din_a[67] & din_b[70])))) # (din_a[68] & (!din_b[69] $ (((!din_a[67]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_558  ) + ( Xd_0__inst_mult_5_557  ))
// Xd_0__inst_mult_5_565  = CARRY(( (!din_a[68] & (((din_a[67] & din_b[70])))) # (din_a[68] & (!din_b[69] $ (((!din_a[67]) # (!din_b[70]))))) ) + ( Xd_0__inst_mult_5_558  ) + ( Xd_0__inst_mult_5_557  ))
// Xd_0__inst_mult_5_566  = SHARE((din_a[68] & (din_b[69] & (din_a[67] & din_b[70]))))

	.dataa(!din_a[68]),
	.datab(!din_b[69]),
	.datac(!din_a[67]),
	.datad(!din_b[70]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_557 ),
	.sharein(Xd_0__inst_mult_5_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_564 ),
	.cout(Xd_0__inst_mult_5_565 ),
	.shareout(Xd_0__inst_mult_5_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_165 (
// Equation(s):
// Xd_0__inst_mult_2_560  = SUM(( GND ) + ( Xd_0__inst_mult_2_554  ) + ( Xd_0__inst_mult_2_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_553 ),
	.sharein(Xd_0__inst_mult_2_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_2_166 (
// Equation(s):
// Xd_0__inst_mult_2_564  = SUM(( (!din_a[32] & (((din_a[31] & din_b[34])))) # (din_a[32] & (!din_b[33] $ (((!din_a[31]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_558  ) + ( Xd_0__inst_mult_2_557  ))
// Xd_0__inst_mult_2_565  = CARRY(( (!din_a[32] & (((din_a[31] & din_b[34])))) # (din_a[32] & (!din_b[33] $ (((!din_a[31]) # (!din_b[34]))))) ) + ( Xd_0__inst_mult_2_558  ) + ( Xd_0__inst_mult_2_557  ))
// Xd_0__inst_mult_2_566  = SHARE((din_a[32] & (din_b[33] & (din_a[31] & din_b[34]))))

	.dataa(!din_a[32]),
	.datab(!din_b[33]),
	.datac(!din_a[31]),
	.datad(!din_b[34]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_557 ),
	.sharein(Xd_0__inst_mult_2_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_564 ),
	.cout(Xd_0__inst_mult_2_565 ),
	.shareout(Xd_0__inst_mult_2_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_163 (
// Equation(s):
// Xd_0__inst_mult_3_564  = SUM(( GND ) + ( Xd_0__inst_mult_3_562  ) + ( Xd_0__inst_mult_3_561  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_561 ),
	.sharein(Xd_0__inst_mult_3_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_3_564 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_161 (
// Equation(s):
// Xd_0__inst_mult_0_556  = SUM(( GND ) + ( Xd_0__inst_mult_0_550  ) + ( Xd_0__inst_mult_0_549  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_549 ),
	.sharein(Xd_0__inst_mult_0_550 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_556 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_0_162 (
// Equation(s):
// Xd_0__inst_mult_0_560  = SUM(( (!din_a[8] & (((din_a[7] & din_b[10])))) # (din_a[8] & (!din_b[9] $ (((!din_a[7]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_554  ) + ( Xd_0__inst_mult_0_553  ))
// Xd_0__inst_mult_0_561  = CARRY(( (!din_a[8] & (((din_a[7] & din_b[10])))) # (din_a[8] & (!din_b[9] $ (((!din_a[7]) # (!din_b[10]))))) ) + ( Xd_0__inst_mult_0_554  ) + ( Xd_0__inst_mult_0_553  ))
// Xd_0__inst_mult_0_562  = SHARE((din_a[8] & (din_b[9] & (din_a[7] & din_b[10]))))

	.dataa(!din_a[8]),
	.datab(!din_b[9]),
	.datac(!din_a[7]),
	.datad(!din_b[10]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_553 ),
	.sharein(Xd_0__inst_mult_0_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_560 ),
	.cout(Xd_0__inst_mult_0_561 ),
	.shareout(Xd_0__inst_mult_0_562 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_162 (
// Equation(s):
// Xd_0__inst_mult_1_560  = SUM(( GND ) + ( Xd_0__inst_mult_1_554  ) + ( Xd_0__inst_mult_1_553  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_553 ),
	.sharein(Xd_0__inst_mult_1_554 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_560 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h000000010000111E),
	.shared_arith("on")
) Xd_0__inst_mult_1_163 (
// Equation(s):
// Xd_0__inst_mult_1_564  = SUM(( (!din_a[20] & (((din_a[19] & din_b[22])))) # (din_a[20] & (!din_b[21] $ (((!din_a[19]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_558  ) + ( Xd_0__inst_mult_1_557  ))
// Xd_0__inst_mult_1_565  = CARRY(( (!din_a[20] & (((din_a[19] & din_b[22])))) # (din_a[20] & (!din_b[21] $ (((!din_a[19]) # (!din_b[22]))))) ) + ( Xd_0__inst_mult_1_558  ) + ( Xd_0__inst_mult_1_557  ))
// Xd_0__inst_mult_1_566  = SHARE((din_a[20] & (din_b[21] & (din_a[19] & din_b[22]))))

	.dataa(!din_a[20]),
	.datab(!din_b[21]),
	.datac(!din_a[19]),
	.datad(!din_b[22]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_557 ),
	.sharein(Xd_0__inst_mult_1_558 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_564 ),
	.cout(Xd_0__inst_mult_1_565 ),
	.shareout(Xd_0__inst_mult_1_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_167 (
// Equation(s):
// Xd_0__inst_mult_4_568  = SUM(( (din_a[56] & din_b[58]) ) + ( Xd_0__inst_mult_4_566  ) + ( Xd_0__inst_mult_4_565  ))
// Xd_0__inst_mult_4_569  = CARRY(( (din_a[56] & din_b[58]) ) + ( Xd_0__inst_mult_4_566  ) + ( Xd_0__inst_mult_4_565  ))
// Xd_0__inst_mult_4_570  = SHARE(GND)

	.dataa(!din_a[56]),
	.datab(!din_b[58]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_565 ),
	.sharein(Xd_0__inst_mult_4_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_568 ),
	.cout(Xd_0__inst_mult_4_569 ),
	.shareout(Xd_0__inst_mult_4_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_167 (
// Equation(s):
// Xd_0__inst_mult_5_568  = SUM(( (din_a[68] & din_b[70]) ) + ( Xd_0__inst_mult_5_566  ) + ( Xd_0__inst_mult_5_565  ))
// Xd_0__inst_mult_5_569  = CARRY(( (din_a[68] & din_b[70]) ) + ( Xd_0__inst_mult_5_566  ) + ( Xd_0__inst_mult_5_565  ))
// Xd_0__inst_mult_5_570  = SHARE(GND)

	.dataa(!din_a[68]),
	.datab(!din_b[70]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_565 ),
	.sharein(Xd_0__inst_mult_5_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_568 ),
	.cout(Xd_0__inst_mult_5_569 ),
	.shareout(Xd_0__inst_mult_5_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_167 (
// Equation(s):
// Xd_0__inst_mult_2_568  = SUM(( (din_a[32] & din_b[34]) ) + ( Xd_0__inst_mult_2_566  ) + ( Xd_0__inst_mult_2_565  ))
// Xd_0__inst_mult_2_569  = CARRY(( (din_a[32] & din_b[34]) ) + ( Xd_0__inst_mult_2_566  ) + ( Xd_0__inst_mult_2_565  ))
// Xd_0__inst_mult_2_570  = SHARE(GND)

	.dataa(!din_a[32]),
	.datab(!din_b[34]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_565 ),
	.sharein(Xd_0__inst_mult_2_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_568 ),
	.cout(Xd_0__inst_mult_2_569 ),
	.shareout(Xd_0__inst_mult_2_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_163 (
// Equation(s):
// Xd_0__inst_mult_0_564  = SUM(( (din_a[8] & din_b[10]) ) + ( Xd_0__inst_mult_0_562  ) + ( Xd_0__inst_mult_0_561  ))
// Xd_0__inst_mult_0_565  = CARRY(( (din_a[8] & din_b[10]) ) + ( Xd_0__inst_mult_0_562  ) + ( Xd_0__inst_mult_0_561  ))
// Xd_0__inst_mult_0_566  = SHARE(GND)

	.dataa(!din_a[8]),
	.datab(!din_b[10]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_561 ),
	.sharein(Xd_0__inst_mult_0_562 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_564 ),
	.cout(Xd_0__inst_mult_0_565 ),
	.shareout(Xd_0__inst_mult_0_566 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_164 (
// Equation(s):
// Xd_0__inst_mult_1_568  = SUM(( (din_a[20] & din_b[22]) ) + ( Xd_0__inst_mult_1_566  ) + ( Xd_0__inst_mult_1_565  ))
// Xd_0__inst_mult_1_569  = CARRY(( (din_a[20] & din_b[22]) ) + ( Xd_0__inst_mult_1_566  ) + ( Xd_0__inst_mult_1_565  ))
// Xd_0__inst_mult_1_570  = SHARE(GND)

	.dataa(!din_a[20]),
	.datab(!din_b[22]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_565 ),
	.sharein(Xd_0__inst_mult_1_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_568 ),
	.cout(Xd_0__inst_mult_1_569 ),
	.shareout(Xd_0__inst_mult_1_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_168 (
// Equation(s):
// Xd_0__inst_mult_4_572  = SUM(( GND ) + ( Xd_0__inst_mult_4_570  ) + ( Xd_0__inst_mult_4_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_569 ),
	.sharein(Xd_0__inst_mult_4_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_4_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_168 (
// Equation(s):
// Xd_0__inst_mult_5_572  = SUM(( GND ) + ( Xd_0__inst_mult_5_570  ) + ( Xd_0__inst_mult_5_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_569 ),
	.sharein(Xd_0__inst_mult_5_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_5_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_168 (
// Equation(s):
// Xd_0__inst_mult_2_572  = SUM(( GND ) + ( Xd_0__inst_mult_2_570  ) + ( Xd_0__inst_mult_2_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_569 ),
	.sharein(Xd_0__inst_mult_2_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_2_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_164 (
// Equation(s):
// Xd_0__inst_mult_0_568  = SUM(( GND ) + ( Xd_0__inst_mult_0_566  ) + ( Xd_0__inst_mult_0_565  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_565 ),
	.sharein(Xd_0__inst_mult_0_566 ),
	.combout(),
	.sumout(Xd_0__inst_mult_0_568 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000000000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_165 (
// Equation(s):
// Xd_0__inst_mult_1_572  = SUM(( GND ) + ( Xd_0__inst_mult_1_570  ) + ( Xd_0__inst_mult_1_569  ))

	.dataa(gnd),
	.datab(gnd),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_569 ),
	.sharein(Xd_0__inst_mult_1_570 ),
	.combout(),
	.sumout(Xd_0__inst_mult_1_572 ),
	.cout(),
	.shareout());

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_169 (
// Equation(s):
// Xd_0__inst_mult_4_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_578  = SHARE((din_a[51] & din_b[49]))

	.dataa(!din_a[51]),
	.datab(!din_b[49]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_577 ),
	.shareout(Xd_0__inst_mult_4_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_169 (
// Equation(s):
// Xd_0__inst_mult_5_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_578  = SHARE((din_a[63] & din_b[61]))

	.dataa(!din_a[63]),
	.datab(!din_b[61]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_577 ),
	.shareout(Xd_0__inst_mult_5_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_169 (
// Equation(s):
// Xd_0__inst_mult_2_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_578  = SHARE((din_a[27] & din_b[25]))

	.dataa(!din_a[27]),
	.datab(!din_b[25]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_577 ),
	.shareout(Xd_0__inst_mult_2_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_164 (
// Equation(s):
// Xd_0__inst_mult_3_569  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_570  = SHARE((din_a[39] & din_b[37]))

	.dataa(!din_a[39]),
	.datab(!din_b[37]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_569 ),
	.shareout(Xd_0__inst_mult_3_570 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_165 (
// Equation(s):
// Xd_0__inst_mult_0_573  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_574  = SHARE((din_a[3] & din_b[1]))

	.dataa(!din_a[3]),
	.datab(!din_b[1]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_573 ),
	.shareout(Xd_0__inst_mult_0_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_4_170 (
// Equation(s):
// Xd_0__inst_mult_4_581  = CARRY(( (din_a[50] & din_b[55]) ) + ( Xd_0__inst_mult_4_362  ) + ( Xd_0__inst_mult_4_361  ))
// Xd_0__inst_mult_4_582  = SHARE((din_a[49] & din_b[56]))

	.dataa(!din_a[50]),
	.datab(!din_b[55]),
	.datac(!din_a[49]),
	.datad(!din_b[56]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_4_361 ),
	.sharein(Xd_0__inst_mult_4_362 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_581 ),
	.shareout(Xd_0__inst_mult_4_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_5_170 (
// Equation(s):
// Xd_0__inst_mult_5_581  = CARRY(( (din_a[62] & din_b[67]) ) + ( Xd_0__inst_mult_5_550  ) + ( Xd_0__inst_mult_5_549  ))
// Xd_0__inst_mult_5_582  = SHARE((din_a[61] & din_b[68]))

	.dataa(!din_a[62]),
	.datab(!din_b[67]),
	.datac(!din_a[61]),
	.datad(!din_b[68]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_5_549 ),
	.sharein(Xd_0__inst_mult_5_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_581 ),
	.shareout(Xd_0__inst_mult_5_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_2_170 (
// Equation(s):
// Xd_0__inst_mult_2_581  = CARRY(( (din_a[26] & din_b[31]) ) + ( Xd_0__inst_mult_2_550  ) + ( Xd_0__inst_mult_2_549  ))
// Xd_0__inst_mult_2_582  = SHARE((din_a[25] & din_b[32]))

	.dataa(!din_a[26]),
	.datab(!din_b[31]),
	.datac(!din_a[25]),
	.datad(!din_b[32]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_2_549 ),
	.sharein(Xd_0__inst_mult_2_550 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_581 ),
	.shareout(Xd_0__inst_mult_2_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_3_165 (
// Equation(s):
// Xd_0__inst_mult_3_573  = CARRY(( (din_a[38] & din_b[43]) ) + ( Xd_0__inst_mult_3_582  ) + ( Xd_0__inst_mult_3_581  ))
// Xd_0__inst_mult_3_574  = SHARE((din_a[37] & din_b[44]))

	.dataa(!din_a[38]),
	.datab(!din_b[43]),
	.datac(!din_a[37]),
	.datad(!din_b[44]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_3_581 ),
	.sharein(Xd_0__inst_mult_3_582 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_573 ),
	.shareout(Xd_0__inst_mult_3_574 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_0_166 (
// Equation(s):
// Xd_0__inst_mult_0_577  = CARRY(( (din_a[2] & din_b[7]) ) + ( Xd_0__inst_mult_0_546  ) + ( Xd_0__inst_mult_0_545  ))
// Xd_0__inst_mult_0_578  = SHARE((din_a[1] & din_b[8]))

	.dataa(!din_a[2]),
	.datab(!din_b[7]),
	.datac(!din_a[1]),
	.datad(!din_b[8]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_0_545 ),
	.sharein(Xd_0__inst_mult_0_546 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_577 ),
	.shareout(Xd_0__inst_mult_0_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000000F00001111),
	.shared_arith("on")
) Xd_0__inst_mult_1_166 (
// Equation(s):
// Xd_0__inst_mult_1_577  = CARRY(( (din_a[14] & din_b[19]) ) + ( Xd_0__inst_mult_1_538  ) + ( Xd_0__inst_mult_1_537  ))
// Xd_0__inst_mult_1_578  = SHARE((din_a[13] & din_b[20]))

	.dataa(!din_a[14]),
	.datab(!din_b[19]),
	.datac(!din_a[13]),
	.datad(!din_b[20]),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(Xd_0__inst_mult_1_537 ),
	.sharein(Xd_0__inst_mult_1_538 ),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_577 ),
	.shareout(Xd_0__inst_mult_1_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_6_171 (
// Equation(s):
// Xd_0__inst_mult_6_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_6_586  = SHARE((din_a[74] & din_b[79]))

	.dataa(!din_a[74]),
	.datab(!din_b[79]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_6_585 ),
	.shareout(Xd_0__inst_mult_6_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_7_171 (
// Equation(s):
// Xd_0__inst_mult_7_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_7_586  = SHARE((din_a[86] & din_b[91]))

	.dataa(!din_a[86]),
	.datab(!din_b[91]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_7_585 ),
	.shareout(Xd_0__inst_mult_7_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_4_171 (
// Equation(s):
// Xd_0__inst_mult_4_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_4_586  = SHARE((din_a[52] & din_b[54]))

	.dataa(!din_a[52]),
	.datab(!din_b[54]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_4_585 ),
	.shareout(Xd_0__inst_mult_4_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_5_171 (
// Equation(s):
// Xd_0__inst_mult_5_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_5_586  = SHARE((din_a[64] & din_b[66]))

	.dataa(!din_a[64]),
	.datab(!din_b[66]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_5_585 ),
	.shareout(Xd_0__inst_mult_5_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_2_171 (
// Equation(s):
// Xd_0__inst_mult_2_585  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_2_586  = SHARE((din_a[28] & din_b[30]))

	.dataa(!din_a[28]),
	.datab(!din_b[30]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_2_585 ),
	.shareout(Xd_0__inst_mult_2_586 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_166 (
// Equation(s):
// Xd_0__inst_mult_3_577  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_578  = SHARE((din_a[40] & din_b[42]))

	.dataa(!din_a[40]),
	.datab(!din_b[42]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_577 ),
	.shareout(Xd_0__inst_mult_3_578 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_0_167 (
// Equation(s):
// Xd_0__inst_mult_0_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_0_582  = SHARE((din_a[4] & din_b[6]))

	.dataa(!din_a[4]),
	.datab(!din_b[6]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_0_581 ),
	.shareout(Xd_0__inst_mult_0_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_1_167 (
// Equation(s):
// Xd_0__inst_mult_1_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_1_582  = SHARE((din_a[16] & din_b[18]))

	.dataa(!din_a[16]),
	.datab(!din_b[18]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_1_581 ),
	.shareout(Xd_0__inst_mult_1_582 ));

twentynm_lcell_comb #(
	.extended_lut("off"),
	.lut_mask(64'h0000111100000000),
	.shared_arith("on")
) Xd_0__inst_mult_3_167 (
// Equation(s):
// Xd_0__inst_mult_3_581  = CARRY(( GND ) + ( !VCC ) + ( !VCC ))
// Xd_0__inst_mult_3_582  = SHARE((din_a[38] & din_b[43]))

	.dataa(!din_a[38]),
	.datab(!din_b[43]),
	.datac(gnd),
	.datad(gnd),
	.datae(gnd),
	.dataf(gnd),
	.datag(gnd),
	.cin(gnd),
	.sharein(gnd),
	.combout(),
	.sumout(),
	.cout(Xd_0__inst_mult_3_581 ),
	.shareout(Xd_0__inst_mult_3_582 ));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [8]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [9]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [10]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [11]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [12]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [13]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [14]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [15]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [16]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [17]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [18]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [19]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [20]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [21]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [22]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [23]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_inst_add_0_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [24]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_inst_dout_25_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_inst_dout [25]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__5__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__6__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__7__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_33_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__8__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_37_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__9__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_41_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__10__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_45_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__11__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_49_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__12__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_53_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__13__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_57_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__14__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_61_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__15__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_65_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__16__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_69_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__17__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_73_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__18__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_77_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__19__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_81_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__20__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_85_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__21__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_89_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__22__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_93_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_1__25_ (
	.clk(clk),
	.d(Xd_0__inst_r_sum1_3__23__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_1__25__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__24_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_97_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__24__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_inst_first_level_0__25_ (
	.clk(clk),
	.d(Xd_0__inst_inst_add_0_101_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_inst_first_level_0__25__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_3__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_3__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_3__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [8]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [9]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [11]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [12]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [13]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [14]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [15]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [16]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [18]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [19]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [20]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [21]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__22_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__22__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_2__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_2__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_2__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_1__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_1__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_1__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_r_sum1_0__23_ (
	.clk(clk),
	.d(Xd_0__inst_a1_0__adder1_inst_dout [23]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_r_sum1_0__23__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_6_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [6]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_7_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [7]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_6__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_7__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_6__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_6__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_7__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_7__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_4_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [4]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_5_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_2_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [2]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_3_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [3]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__0__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_0_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [0]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign_1_ (
	.clk(clk),
	.d(Xd_0__inst_sign1 [1]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_6_ (
	.clk(clk),
	.d(Xd_0__inst_i29_1_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [6]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_7_ (
	.clk(clk),
	.d(Xd_0__inst_i29_5_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [7]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__1__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__2__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__3__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_4__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_5__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_2__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_3__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_0__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_product1_1__4__q ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_6__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_6_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_6__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_7__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_7_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_7__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__5_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__5__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__6_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__6__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__7_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__7__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__8_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__8__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_188 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__9_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__9__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_192 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__10_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__10__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_196 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__11_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__11__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_200 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__12_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__12__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_204 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__13_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__13__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_208 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__14_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__14__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_212 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__15_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__15__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_216 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__16_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__16__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_220 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__17_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__17__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_224 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__18_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__18__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_228 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__19_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__19__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_232 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__20_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__20__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_4__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_4__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_5__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_5__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_2__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_236 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_2__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_3__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_3__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_0__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_0__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product_1__21_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product_1__21__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_4_ (
	.clk(clk),
	.d(Xd_0__inst_i29_9_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [4]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_5_ (
	.clk(clk),
	.d(Xd_0__inst_i29_13_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [5]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_240 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_2_ (
	.clk(clk),
	.d(Xd_0__inst_i29_17_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [2]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_3_ (
	.clk(clk),
	.d(Xd_0__inst_i29_21_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [3]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__0_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__0__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_0_ (
	.clk(clk),
	.d(Xd_0__inst_i29_25_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [0]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_sign1_1_ (
	.clk(clk),
	.d(Xd_0__inst_i29_29_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_sign1 [1]),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__1_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_180 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__1__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_248 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__2_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__2__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__3_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__3__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_4__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_4_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_4__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_5__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_5_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_5__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_2__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_2_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_2__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_3__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_3_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_3__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_0__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_0_268 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_0__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_product1_1__4_ (
	.clk(clk),
	.d(Xd_0__inst_mult_1_260 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_product1_1__4__q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_256 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_244 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_177 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_22 (
	.clk(clk),
	.d(din_a[82]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_23 (
	.clk(clk),
	.d(din_b[77]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_22 (
	.clk(clk),
	.d(din_a[94]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_23 (
	.clk(clk),
	.d(din_b[89]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_6_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_6_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_6_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_7_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_7_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_7_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_272 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_0 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_0_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_1 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_1_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_280 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_2 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_284 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_2_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_3 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_3_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_288 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_4 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_292 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_4_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_5 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_5_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_6 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_300 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_6_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_7 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_7_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_304 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_8 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_308 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_8_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_9 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_9_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_312 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_10 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_316 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_10_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_11 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_11_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_320 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_12 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_324 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_12_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_13 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_13_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_328 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_296 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_276 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_14 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_332 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_14_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_15 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_15_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_336 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_264 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_252 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_16 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_340 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_16_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_17 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_17_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_344 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_184 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_173 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_18 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_348 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_18_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_19 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_19_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_22 (
	.clk(clk),
	.d(din_a[58]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_23 (
	.clk(clk),
	.d(din_b[53]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_22 (
	.clk(clk),
	.d(din_a[70]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_23 (
	.clk(clk),
	.d(din_b[65]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_352 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_22 (
	.clk(clk),
	.d(din_a[34]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_23 (
	.clk(clk),
	.d(din_b[29]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_176 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_384 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_22 (
	.clk(clk),
	.d(din_a[46]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_23 (
	.clk(clk),
	.d(din_b[41]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_169 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_22 (
	.clk(clk),
	.d(din_a[10]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_23 (
	.clk(clk),
	.d(din_b[5]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_20 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_356 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_20_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_21 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_21_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_22 (
	.clk(clk),
	.d(din_a[22]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_22_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_23 (
	.clk(clk),
	.d(din_b[17]),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_23_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_360 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_388 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_24 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_24_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_25 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_25_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_364 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_392 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_26 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_26_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_27 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_27_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_59_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_368 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_396 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_28 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_28_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_29 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_47_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_29_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_372 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_400 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_51_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_30 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_30_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_31 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_35_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_31_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_4_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_4_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_4_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_5_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_5_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_5_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_376 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_2_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_2_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_2_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_404 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_3_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_3_55_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_3_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_0_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_0_43_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_0_33_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_32 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_380 ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_32_q ),
	.prn(vcc));

dffeas #(
	.is_wysiwyg("true"),
	.power_up("low")
) Xd_0__inst_mult_1_33 (
	.clk(clk),
	.d(Xd_0__inst_mult_1_39_sumout ),
	.asdata(vcc),
	.clrn(vcc),
	.aload(gnd),
	.sclr(gnd),
	.sload(gnd),
	.ena(vcc),
	.devclrn(),
	.devpor(),
	.q(Xd_0__inst_mult_1_33_q ),
	.prn(vcc));

assign dout[0] = Xd_0__inst_inst_inst_dout [0];

assign dout[1] = Xd_0__inst_inst_inst_dout [1];

assign dout[2] = Xd_0__inst_inst_inst_dout [2];

assign dout[3] = Xd_0__inst_inst_inst_dout [3];

assign dout[4] = Xd_0__inst_inst_inst_dout [4];

assign dout[5] = Xd_0__inst_inst_inst_dout [5];

assign dout[6] = Xd_0__inst_inst_inst_dout [6];

assign dout[7] = Xd_0__inst_inst_inst_dout [7];

assign dout[8] = Xd_0__inst_inst_inst_dout [8];

assign dout[9] = Xd_0__inst_inst_inst_dout [9];

assign dout[10] = Xd_0__inst_inst_inst_dout [10];

assign dout[11] = Xd_0__inst_inst_inst_dout [11];

assign dout[12] = Xd_0__inst_inst_inst_dout [12];

assign dout[13] = Xd_0__inst_inst_inst_dout [13];

assign dout[14] = Xd_0__inst_inst_inst_dout [14];

assign dout[15] = Xd_0__inst_inst_inst_dout [15];

assign dout[16] = Xd_0__inst_inst_inst_dout [16];

assign dout[17] = Xd_0__inst_inst_inst_dout [17];

assign dout[18] = Xd_0__inst_inst_inst_dout [18];

assign dout[19] = Xd_0__inst_inst_inst_dout [19];

assign dout[20] = Xd_0__inst_inst_inst_dout [20];

assign dout[21] = Xd_0__inst_inst_inst_dout [21];

assign dout[22] = Xd_0__inst_inst_inst_dout [22];

assign dout[23] = Xd_0__inst_inst_inst_dout [23];

assign dout[24] = Xd_0__inst_inst_inst_dout [24];

assign dout[25] = Xd_0__inst_inst_inst_dout [25];

endmodule
